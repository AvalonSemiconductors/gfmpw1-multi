magic
tech gf180mcuD
magscale 1 10
timestamp 1700061065
<< metal1 >>
rect 1344 42362 44576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 44576 42362
rect 1344 42276 44576 42310
rect 32846 42082 32898 42094
rect 32846 42018 32898 42030
rect 34078 42082 34130 42094
rect 34078 42018 34130 42030
rect 43598 42082 43650 42094
rect 43598 42018 43650 42030
rect 43710 42082 43762 42094
rect 43710 42018 43762 42030
rect 33854 41970 33906 41982
rect 33058 41918 33070 41970
rect 33122 41918 33134 41970
rect 33854 41906 33906 41918
rect 34190 41970 34242 41982
rect 43026 41918 43038 41970
rect 43090 41918 43102 41970
rect 34190 41906 34242 41918
rect 32510 41858 32562 41870
rect 41906 41806 41918 41858
rect 41970 41806 41982 41858
rect 32510 41794 32562 41806
rect 43710 41746 43762 41758
rect 43710 41682 43762 41694
rect 1344 41578 44576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 44576 41578
rect 1344 41492 44576 41526
rect 34626 41246 34638 41298
rect 34690 41246 34702 41298
rect 40898 41246 40910 41298
rect 40962 41246 40974 41298
rect 44146 41246 44158 41298
rect 44210 41246 44222 41298
rect 29934 41186 29986 41198
rect 29934 41122 29986 41134
rect 30158 41186 30210 41198
rect 35534 41186 35586 41198
rect 31826 41134 31838 41186
rect 31890 41134 31902 41186
rect 38098 41134 38110 41186
rect 38162 41134 38174 41186
rect 41234 41134 41246 41186
rect 41298 41134 41310 41186
rect 30158 41122 30210 41134
rect 35534 41122 35586 41134
rect 36094 41074 36146 41086
rect 32498 41022 32510 41074
rect 32562 41022 32574 41074
rect 38770 41022 38782 41074
rect 38834 41022 38846 41074
rect 42018 41022 42030 41074
rect 42082 41022 42094 41074
rect 36094 41010 36146 41022
rect 34862 40962 34914 40974
rect 29586 40910 29598 40962
rect 29650 40910 29662 40962
rect 34862 40898 34914 40910
rect 34974 40962 35026 40974
rect 34974 40898 35026 40910
rect 35198 40962 35250 40974
rect 35198 40898 35250 40910
rect 35870 40962 35922 40974
rect 35870 40898 35922 40910
rect 35982 40962 36034 40974
rect 35982 40898 36034 40910
rect 1344 40794 44576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 44576 40794
rect 1344 40708 44576 40742
rect 32510 40626 32562 40638
rect 32510 40562 32562 40574
rect 38222 40626 38274 40638
rect 38222 40562 38274 40574
rect 39118 40626 39170 40638
rect 39118 40562 39170 40574
rect 39342 40626 39394 40638
rect 39342 40562 39394 40574
rect 31838 40514 31890 40526
rect 39566 40514 39618 40526
rect 33954 40462 33966 40514
rect 34018 40462 34030 40514
rect 36530 40462 36542 40514
rect 36594 40462 36606 40514
rect 31838 40450 31890 40462
rect 39566 40450 39618 40462
rect 39678 40514 39730 40526
rect 39678 40450 39730 40462
rect 40238 40514 40290 40526
rect 40238 40450 40290 40462
rect 40350 40514 40402 40526
rect 40350 40450 40402 40462
rect 30046 40402 30098 40414
rect 26898 40350 26910 40402
rect 26962 40350 26974 40402
rect 30046 40338 30098 40350
rect 30270 40402 30322 40414
rect 30270 40338 30322 40350
rect 30718 40402 30770 40414
rect 32174 40402 32226 40414
rect 31602 40350 31614 40402
rect 31666 40350 31678 40402
rect 30718 40338 30770 40350
rect 32174 40338 32226 40350
rect 33070 40402 33122 40414
rect 33742 40402 33794 40414
rect 39006 40402 39058 40414
rect 33506 40350 33518 40402
rect 33570 40350 33582 40402
rect 37314 40350 37326 40402
rect 37378 40350 37390 40402
rect 33070 40338 33122 40350
rect 33742 40338 33794 40350
rect 39006 40338 39058 40350
rect 39902 40402 39954 40414
rect 40898 40350 40910 40402
rect 40962 40350 40974 40402
rect 39902 40338 39954 40350
rect 30158 40290 30210 40302
rect 27570 40238 27582 40290
rect 27634 40238 27646 40290
rect 29698 40238 29710 40290
rect 29762 40238 29774 40290
rect 30158 40226 30210 40238
rect 34078 40290 34130 40302
rect 38110 40290 38162 40302
rect 34402 40238 34414 40290
rect 34466 40238 34478 40290
rect 34078 40226 34130 40238
rect 38110 40226 38162 40238
rect 38670 40290 38722 40302
rect 41682 40238 41694 40290
rect 41746 40238 41758 40290
rect 43810 40238 43822 40290
rect 43874 40238 43886 40290
rect 38670 40226 38722 40238
rect 38558 40178 38610 40190
rect 38558 40114 38610 40126
rect 40238 40178 40290 40190
rect 40238 40114 40290 40126
rect 1344 40010 44576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 44576 40010
rect 1344 39924 44576 39958
rect 27694 39842 27746 39854
rect 27694 39778 27746 39790
rect 37102 39842 37154 39854
rect 37102 39778 37154 39790
rect 27582 39730 27634 39742
rect 26786 39678 26798 39730
rect 26850 39678 26862 39730
rect 27582 39666 27634 39678
rect 28590 39730 28642 39742
rect 36094 39730 36146 39742
rect 29922 39678 29934 39730
rect 29986 39678 29998 39730
rect 32050 39678 32062 39730
rect 32114 39678 32126 39730
rect 35298 39678 35310 39730
rect 35362 39678 35374 39730
rect 38322 39678 38334 39730
rect 38386 39678 38398 39730
rect 40450 39678 40462 39730
rect 40514 39678 40526 39730
rect 41122 39678 41134 39730
rect 41186 39678 41198 39730
rect 28590 39666 28642 39678
rect 36094 39666 36146 39678
rect 28366 39618 28418 39630
rect 35646 39618 35698 39630
rect 26674 39566 26686 39618
rect 26738 39566 26750 39618
rect 29250 39566 29262 39618
rect 29314 39566 29326 39618
rect 32498 39566 32510 39618
rect 32562 39566 32574 39618
rect 28366 39554 28418 39566
rect 35646 39554 35698 39566
rect 36990 39618 37042 39630
rect 37538 39566 37550 39618
rect 37602 39566 37614 39618
rect 43922 39566 43934 39618
rect 43986 39566 43998 39618
rect 36990 39554 37042 39566
rect 27022 39506 27074 39518
rect 35870 39506 35922 39518
rect 33170 39454 33182 39506
rect 33234 39454 33246 39506
rect 27022 39442 27074 39454
rect 35870 39442 35922 39454
rect 36206 39506 36258 39518
rect 43250 39454 43262 39506
rect 43314 39454 43326 39506
rect 36206 39442 36258 39454
rect 27470 39394 27522 39406
rect 37102 39394 37154 39406
rect 28018 39342 28030 39394
rect 28082 39342 28094 39394
rect 27470 39330 27522 39342
rect 37102 39330 37154 39342
rect 1344 39226 44576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 44576 39226
rect 1344 39140 44576 39174
rect 30382 39058 30434 39070
rect 30382 38994 30434 39006
rect 30830 39058 30882 39070
rect 36318 39058 36370 39070
rect 31938 39006 31950 39058
rect 32002 39006 32014 39058
rect 30830 38994 30882 39006
rect 36318 38994 36370 39006
rect 38670 39058 38722 39070
rect 38670 38994 38722 39006
rect 39790 39058 39842 39070
rect 39790 38994 39842 39006
rect 41246 39058 41298 39070
rect 41246 38994 41298 39006
rect 43150 39058 43202 39070
rect 43150 38994 43202 39006
rect 30494 38946 30546 38958
rect 30494 38882 30546 38894
rect 31278 38946 31330 38958
rect 31278 38882 31330 38894
rect 31502 38946 31554 38958
rect 31502 38882 31554 38894
rect 36430 38946 36482 38958
rect 36430 38882 36482 38894
rect 38222 38946 38274 38958
rect 38222 38882 38274 38894
rect 38782 38946 38834 38958
rect 38782 38882 38834 38894
rect 39678 38946 39730 38958
rect 39678 38882 39730 38894
rect 30606 38834 30658 38846
rect 27234 38782 27246 38834
rect 27298 38782 27310 38834
rect 30606 38770 30658 38782
rect 32510 38834 32562 38846
rect 37886 38834 37938 38846
rect 40014 38834 40066 38846
rect 33058 38782 33070 38834
rect 33122 38782 33134 38834
rect 38546 38782 38558 38834
rect 38610 38782 38622 38834
rect 39218 38782 39230 38834
rect 39282 38782 39294 38834
rect 41010 38782 41022 38834
rect 41074 38782 41086 38834
rect 44146 38782 44158 38834
rect 44210 38782 44222 38834
rect 32510 38770 32562 38782
rect 37886 38770 37938 38782
rect 40014 38770 40066 38782
rect 32286 38722 32338 38734
rect 27906 38670 27918 38722
rect 27970 38670 27982 38722
rect 30034 38670 30046 38722
rect 30098 38670 30110 38722
rect 31602 38670 31614 38722
rect 31666 38670 31678 38722
rect 33842 38670 33854 38722
rect 33906 38670 33918 38722
rect 35970 38670 35982 38722
rect 36034 38670 36046 38722
rect 39666 38670 39678 38722
rect 39730 38670 39742 38722
rect 32286 38658 32338 38670
rect 37998 38610 38050 38622
rect 37998 38546 38050 38558
rect 1344 38442 44576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 44576 38442
rect 1344 38356 44576 38390
rect 43150 38274 43202 38286
rect 43150 38210 43202 38222
rect 29262 38162 29314 38174
rect 29262 38098 29314 38110
rect 30158 38162 30210 38174
rect 30158 38098 30210 38110
rect 33182 38162 33234 38174
rect 34402 38110 34414 38162
rect 34466 38110 34478 38162
rect 33182 38098 33234 38110
rect 29038 38050 29090 38062
rect 29038 37986 29090 37998
rect 29486 38050 29538 38062
rect 29486 37986 29538 37998
rect 29710 38050 29762 38062
rect 29710 37986 29762 37998
rect 30046 38050 30098 38062
rect 30046 37986 30098 37998
rect 30718 38050 30770 38062
rect 30718 37986 30770 37998
rect 33294 38050 33346 38062
rect 35086 38050 35138 38062
rect 40126 38050 40178 38062
rect 34066 37998 34078 38050
rect 34130 37998 34142 38050
rect 37202 37998 37214 38050
rect 37266 37998 37278 38050
rect 33294 37986 33346 37998
rect 35086 37986 35138 37998
rect 40126 37986 40178 37998
rect 40574 38050 40626 38062
rect 40574 37986 40626 37998
rect 40910 38050 40962 38062
rect 40910 37986 40962 37998
rect 41246 38050 41298 38062
rect 41246 37986 41298 37998
rect 41582 38050 41634 38062
rect 41582 37986 41634 37998
rect 43598 38050 43650 38062
rect 43598 37986 43650 37998
rect 43934 38050 43986 38062
rect 43934 37986 43986 37998
rect 30270 37938 30322 37950
rect 30270 37874 30322 37886
rect 33630 37938 33682 37950
rect 40462 37938 40514 37950
rect 35410 37886 35422 37938
rect 35474 37886 35486 37938
rect 36978 37886 36990 37938
rect 37042 37886 37054 37938
rect 33630 37874 33682 37886
rect 40462 37874 40514 37886
rect 40798 37938 40850 37950
rect 40798 37874 40850 37886
rect 41358 37938 41410 37950
rect 42478 37938 42530 37950
rect 41794 37886 41806 37938
rect 41858 37886 41870 37938
rect 41358 37874 41410 37886
rect 42478 37874 42530 37886
rect 43038 37938 43090 37950
rect 43038 37874 43090 37886
rect 43150 37938 43202 37950
rect 43150 37874 43202 37886
rect 43710 37938 43762 37950
rect 43710 37874 43762 37886
rect 31838 37826 31890 37838
rect 31838 37762 31890 37774
rect 33070 37826 33122 37838
rect 33070 37762 33122 37774
rect 40238 37826 40290 37838
rect 40238 37762 40290 37774
rect 42142 37826 42194 37838
rect 42142 37762 42194 37774
rect 42590 37826 42642 37838
rect 42590 37762 42642 37774
rect 42814 37826 42866 37838
rect 42814 37762 42866 37774
rect 1344 37658 44576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 44576 37658
rect 1344 37572 44576 37606
rect 29934 37490 29986 37502
rect 29934 37426 29986 37438
rect 33742 37490 33794 37502
rect 33742 37426 33794 37438
rect 39118 37490 39170 37502
rect 39118 37426 39170 37438
rect 26238 37378 26290 37390
rect 29822 37378 29874 37390
rect 27794 37326 27806 37378
rect 27858 37326 27870 37378
rect 26238 37314 26290 37326
rect 29822 37314 29874 37326
rect 33630 37378 33682 37390
rect 38446 37378 38498 37390
rect 36978 37326 36990 37378
rect 37042 37326 37054 37378
rect 33630 37314 33682 37326
rect 38446 37314 38498 37326
rect 38782 37378 38834 37390
rect 38782 37314 38834 37326
rect 41134 37378 41186 37390
rect 41134 37314 41186 37326
rect 30158 37266 30210 37278
rect 39454 37266 39506 37278
rect 26114 37214 26126 37266
rect 26178 37214 26190 37266
rect 26898 37214 26910 37266
rect 26962 37214 26974 37266
rect 27234 37214 27246 37266
rect 27298 37214 27310 37266
rect 28018 37214 28030 37266
rect 28082 37214 28094 37266
rect 33954 37214 33966 37266
rect 34018 37214 34030 37266
rect 36754 37214 36766 37266
rect 36818 37214 36830 37266
rect 37650 37214 37662 37266
rect 37714 37214 37726 37266
rect 38210 37214 38222 37266
rect 38274 37214 38286 37266
rect 30158 37202 30210 37214
rect 39454 37202 39506 37214
rect 41022 37266 41074 37278
rect 41022 37202 41074 37214
rect 41358 37266 41410 37278
rect 41570 37214 41582 37266
rect 41634 37214 41646 37266
rect 41358 37202 41410 37214
rect 25230 37154 25282 37166
rect 25230 37090 25282 37102
rect 38334 37154 38386 37166
rect 38334 37090 38386 37102
rect 39566 37154 39618 37166
rect 39566 37090 39618 37102
rect 25342 37042 25394 37054
rect 37998 37042 38050 37054
rect 27122 36990 27134 37042
rect 27186 36990 27198 37042
rect 37202 36990 37214 37042
rect 37266 37039 37278 37042
rect 37538 37039 37550 37042
rect 37266 36993 37550 37039
rect 37266 36990 37278 36993
rect 37538 36990 37550 36993
rect 37602 36990 37614 37042
rect 43474 36990 43486 37042
rect 43538 36990 43550 37042
rect 25342 36978 25394 36990
rect 37998 36978 38050 36990
rect 1344 36874 44576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 44576 36874
rect 1344 36788 44576 36822
rect 7298 36542 7310 36594
rect 7362 36542 7374 36594
rect 34850 36542 34862 36594
rect 34914 36542 34926 36594
rect 38658 36542 38670 36594
rect 38722 36542 38734 36594
rect 40786 36542 40798 36594
rect 40850 36542 40862 36594
rect 41122 36542 41134 36594
rect 41186 36542 41198 36594
rect 15598 36482 15650 36494
rect 27134 36482 27186 36494
rect 10098 36430 10110 36482
rect 10162 36430 10174 36482
rect 16034 36430 16046 36482
rect 16098 36430 16110 36482
rect 25890 36430 25902 36482
rect 25954 36430 25966 36482
rect 26450 36430 26462 36482
rect 26514 36430 26526 36482
rect 31938 36430 31950 36482
rect 32002 36430 32014 36482
rect 37874 36430 37886 36482
rect 37938 36430 37950 36482
rect 43922 36430 43934 36482
rect 43986 36430 43998 36482
rect 15598 36418 15650 36430
rect 27134 36418 27186 36430
rect 26910 36370 26962 36382
rect 9426 36318 9438 36370
rect 9490 36318 9502 36370
rect 26910 36306 26962 36318
rect 27470 36370 27522 36382
rect 27470 36306 27522 36318
rect 28030 36370 28082 36382
rect 32722 36318 32734 36370
rect 32786 36318 32798 36370
rect 43250 36318 43262 36370
rect 43314 36318 43326 36370
rect 28030 36306 28082 36318
rect 19070 36258 19122 36270
rect 18274 36206 18286 36258
rect 18338 36206 18350 36258
rect 19070 36194 19122 36206
rect 19406 36258 19458 36270
rect 27246 36258 27298 36270
rect 23538 36206 23550 36258
rect 23602 36206 23614 36258
rect 19406 36194 19458 36206
rect 27246 36194 27298 36206
rect 27358 36258 27410 36270
rect 27358 36194 27410 36206
rect 27918 36258 27970 36270
rect 27918 36194 27970 36206
rect 1344 36090 44576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 44576 36090
rect 1344 36004 44576 36038
rect 17726 35922 17778 35934
rect 10434 35870 10446 35922
rect 10498 35870 10510 35922
rect 17726 35858 17778 35870
rect 35982 35922 36034 35934
rect 40014 35922 40066 35934
rect 39330 35870 39342 35922
rect 39394 35870 39406 35922
rect 35982 35858 36034 35870
rect 40014 35858 40066 35870
rect 15822 35810 15874 35822
rect 15822 35746 15874 35758
rect 16158 35810 16210 35822
rect 16158 35746 16210 35758
rect 16494 35810 16546 35822
rect 16494 35746 16546 35758
rect 17502 35810 17554 35822
rect 18622 35810 18674 35822
rect 18274 35758 18286 35810
rect 18338 35758 18350 35810
rect 17502 35746 17554 35758
rect 18622 35746 18674 35758
rect 19294 35810 19346 35822
rect 19294 35746 19346 35758
rect 23550 35810 23602 35822
rect 23550 35746 23602 35758
rect 31838 35810 31890 35822
rect 31838 35746 31890 35758
rect 35534 35810 35586 35822
rect 36754 35758 36766 35810
rect 36818 35758 36830 35810
rect 43026 35758 43038 35810
rect 43090 35758 43102 35810
rect 35534 35746 35586 35758
rect 10782 35698 10834 35710
rect 17390 35698 17442 35710
rect 16706 35646 16718 35698
rect 16770 35646 16782 35698
rect 10782 35634 10834 35646
rect 17390 35634 17442 35646
rect 17950 35698 18002 35710
rect 24110 35698 24162 35710
rect 18834 35646 18846 35698
rect 18898 35646 18910 35698
rect 19506 35646 19518 35698
rect 19570 35646 19582 35698
rect 20290 35646 20302 35698
rect 20354 35646 20366 35698
rect 17950 35634 18002 35646
rect 24110 35634 24162 35646
rect 24222 35698 24274 35710
rect 24222 35634 24274 35646
rect 24446 35698 24498 35710
rect 29598 35698 29650 35710
rect 24658 35646 24670 35698
rect 24722 35646 24734 35698
rect 25442 35646 25454 35698
rect 25506 35646 25518 35698
rect 26002 35646 26014 35698
rect 26066 35646 26078 35698
rect 29026 35646 29038 35698
rect 29090 35646 29102 35698
rect 29362 35646 29374 35698
rect 29426 35646 29438 35698
rect 24446 35634 24498 35646
rect 29598 35634 29650 35646
rect 32174 35698 32226 35710
rect 32174 35634 32226 35646
rect 32958 35698 33010 35710
rect 32958 35634 33010 35646
rect 33406 35698 33458 35710
rect 33406 35634 33458 35646
rect 33630 35698 33682 35710
rect 36318 35698 36370 35710
rect 35746 35646 35758 35698
rect 35810 35646 35822 35698
rect 37426 35646 37438 35698
rect 37490 35646 37502 35698
rect 37650 35646 37662 35698
rect 37714 35646 37726 35698
rect 38770 35646 38782 35698
rect 38834 35646 38846 35698
rect 38994 35646 39006 35698
rect 39058 35646 39070 35698
rect 39554 35646 39566 35698
rect 39618 35646 39630 35698
rect 40226 35646 40238 35698
rect 40290 35646 40302 35698
rect 43810 35646 43822 35698
rect 43874 35646 43886 35698
rect 33630 35634 33682 35646
rect 36318 35634 36370 35646
rect 24334 35586 24386 35598
rect 28702 35586 28754 35598
rect 20962 35534 20974 35586
rect 21026 35534 21038 35586
rect 23090 35534 23102 35586
rect 23154 35534 23166 35586
rect 28354 35534 28366 35586
rect 28418 35534 28430 35586
rect 24334 35522 24386 35534
rect 28702 35522 28754 35534
rect 28814 35586 28866 35598
rect 28814 35522 28866 35534
rect 33182 35586 33234 35598
rect 35410 35534 35422 35586
rect 35474 35534 35486 35586
rect 40898 35534 40910 35586
rect 40962 35534 40974 35586
rect 33182 35522 33234 35534
rect 23438 35474 23490 35486
rect 23438 35410 23490 35422
rect 29710 35474 29762 35486
rect 29710 35410 29762 35422
rect 36430 35474 36482 35486
rect 36430 35410 36482 35422
rect 37102 35474 37154 35486
rect 37102 35410 37154 35422
rect 1344 35306 44576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 44576 35306
rect 1344 35220 44576 35254
rect 38334 35138 38386 35150
rect 29362 35086 29374 35138
rect 29426 35086 29438 35138
rect 38334 35074 38386 35086
rect 39790 35138 39842 35150
rect 39790 35074 39842 35086
rect 26126 35026 26178 35038
rect 31054 35026 31106 35038
rect 9314 34974 9326 35026
rect 9378 34974 9390 35026
rect 11442 34974 11454 35026
rect 11506 34974 11518 35026
rect 24882 34974 24894 35026
rect 24946 34974 24958 35026
rect 27346 34974 27358 35026
rect 27410 34974 27422 35026
rect 32274 34974 32286 35026
rect 32338 34974 32350 35026
rect 34402 34974 34414 35026
rect 34466 34974 34478 35026
rect 41906 34974 41918 35026
rect 41970 34974 41982 35026
rect 44034 34974 44046 35026
rect 44098 34974 44110 35026
rect 26126 34962 26178 34974
rect 31054 34962 31106 34974
rect 25230 34914 25282 34926
rect 29598 34914 29650 34926
rect 35310 34914 35362 34926
rect 8642 34862 8654 34914
rect 8706 34862 8718 34914
rect 16146 34862 16158 34914
rect 16210 34862 16222 34914
rect 16818 34862 16830 34914
rect 16882 34862 16894 34914
rect 18946 34862 18958 34914
rect 19010 34862 19022 34914
rect 21970 34862 21982 34914
rect 22034 34862 22046 34914
rect 22530 34862 22542 34914
rect 22594 34862 22606 34914
rect 27010 34862 27022 34914
rect 27074 34862 27086 34914
rect 27458 34862 27470 34914
rect 27522 34862 27534 34914
rect 29138 34862 29150 34914
rect 29202 34862 29214 34914
rect 31602 34862 31614 34914
rect 31666 34862 31678 34914
rect 25230 34850 25282 34862
rect 29598 34850 29650 34862
rect 35310 34850 35362 34862
rect 35422 34914 35474 34926
rect 36094 34914 36146 34926
rect 35522 34862 35534 34914
rect 35586 34862 35598 34914
rect 35422 34850 35474 34862
rect 36094 34850 36146 34862
rect 36206 34914 36258 34926
rect 40014 34914 40066 34926
rect 38322 34862 38334 34914
rect 38386 34862 38398 34914
rect 36206 34850 36258 34862
rect 40014 34850 40066 34862
rect 40798 34914 40850 34926
rect 41234 34862 41246 34914
rect 41298 34862 41310 34914
rect 40798 34850 40850 34862
rect 15822 34802 15874 34814
rect 15822 34738 15874 34750
rect 15934 34802 15986 34814
rect 15934 34738 15986 34750
rect 20414 34802 20466 34814
rect 20414 34738 20466 34750
rect 20526 34802 20578 34814
rect 20526 34738 20578 34750
rect 25342 34802 25394 34814
rect 25342 34738 25394 34750
rect 26462 34802 26514 34814
rect 29934 34802 29986 34814
rect 28130 34750 28142 34802
rect 28194 34750 28206 34802
rect 26462 34738 26514 34750
rect 29934 34738 29986 34750
rect 31166 34802 31218 34814
rect 31166 34738 31218 34750
rect 35870 34802 35922 34814
rect 38670 34802 38722 34814
rect 36978 34750 36990 34802
rect 37042 34750 37054 34802
rect 37650 34750 37662 34802
rect 37714 34750 37726 34802
rect 35870 34738 35922 34750
rect 38670 34738 38722 34750
rect 40462 34802 40514 34814
rect 40462 34738 40514 34750
rect 15598 34690 15650 34702
rect 15598 34626 15650 34638
rect 19966 34690 20018 34702
rect 19966 34626 20018 34638
rect 20190 34690 20242 34702
rect 20190 34626 20242 34638
rect 25566 34690 25618 34702
rect 25566 34626 25618 34638
rect 25902 34690 25954 34702
rect 25902 34626 25954 34638
rect 26014 34690 26066 34702
rect 26014 34626 26066 34638
rect 26238 34690 26290 34702
rect 30942 34690 30994 34702
rect 29474 34638 29486 34690
rect 29538 34638 29550 34690
rect 26238 34626 26290 34638
rect 30942 34626 30994 34638
rect 37326 34690 37378 34702
rect 37326 34626 37378 34638
rect 37998 34690 38050 34702
rect 39442 34638 39454 34690
rect 39506 34638 39518 34690
rect 37998 34626 38050 34638
rect 1344 34522 44576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 44576 34522
rect 1344 34436 44576 34470
rect 16270 34354 16322 34366
rect 20974 34354 21026 34366
rect 20178 34302 20190 34354
rect 20242 34302 20254 34354
rect 16270 34290 16322 34302
rect 20974 34290 21026 34302
rect 24558 34354 24610 34366
rect 24558 34290 24610 34302
rect 26462 34354 26514 34366
rect 26462 34290 26514 34302
rect 30942 34354 30994 34366
rect 30942 34290 30994 34302
rect 39678 34354 39730 34366
rect 39678 34290 39730 34302
rect 40350 34354 40402 34366
rect 40350 34290 40402 34302
rect 41806 34354 41858 34366
rect 41806 34290 41858 34302
rect 43262 34354 43314 34366
rect 43262 34290 43314 34302
rect 43486 34354 43538 34366
rect 43486 34290 43538 34302
rect 8206 34242 8258 34254
rect 8206 34178 8258 34190
rect 8654 34242 8706 34254
rect 8654 34178 8706 34190
rect 11230 34242 11282 34254
rect 11230 34178 11282 34190
rect 24446 34242 24498 34254
rect 24446 34178 24498 34190
rect 25790 34242 25842 34254
rect 30382 34242 30434 34254
rect 27346 34190 27358 34242
rect 27410 34190 27422 34242
rect 25790 34178 25842 34190
rect 30382 34178 30434 34190
rect 31054 34242 31106 34254
rect 31054 34178 31106 34190
rect 32286 34242 32338 34254
rect 32286 34178 32338 34190
rect 32510 34242 32562 34254
rect 36990 34242 37042 34254
rect 36642 34190 36654 34242
rect 36706 34190 36718 34242
rect 32510 34178 32562 34190
rect 36990 34178 37042 34190
rect 37774 34242 37826 34254
rect 40014 34242 40066 34254
rect 39330 34190 39342 34242
rect 39394 34190 39406 34242
rect 37774 34178 37826 34190
rect 40014 34178 40066 34190
rect 40910 34242 40962 34254
rect 40910 34178 40962 34190
rect 41246 34242 41298 34254
rect 41246 34178 41298 34190
rect 42590 34242 42642 34254
rect 42590 34178 42642 34190
rect 43150 34242 43202 34254
rect 43150 34178 43202 34190
rect 8990 34130 9042 34142
rect 7970 34078 7982 34130
rect 8034 34078 8046 34130
rect 8990 34066 9042 34078
rect 9886 34130 9938 34142
rect 17278 34130 17330 34142
rect 24782 34130 24834 34142
rect 10546 34078 10558 34130
rect 10610 34078 10622 34130
rect 11442 34078 11454 34130
rect 11506 34078 11518 34130
rect 12674 34078 12686 34130
rect 12738 34078 12750 34130
rect 13122 34078 13134 34130
rect 13186 34078 13198 34130
rect 15362 34078 15374 34130
rect 15426 34078 15438 34130
rect 17938 34078 17950 34130
rect 18002 34078 18014 34130
rect 21186 34078 21198 34130
rect 21250 34078 21262 34130
rect 21970 34078 21982 34130
rect 22034 34078 22046 34130
rect 9886 34066 9938 34078
rect 17278 34066 17330 34078
rect 24782 34066 24834 34078
rect 25678 34130 25730 34142
rect 25678 34066 25730 34078
rect 26238 34130 26290 34142
rect 28926 34130 28978 34142
rect 30606 34130 30658 34142
rect 28242 34078 28254 34130
rect 28306 34078 28318 34130
rect 29474 34078 29486 34130
rect 29538 34078 29550 34130
rect 26238 34066 26290 34078
rect 28926 34066 28978 34078
rect 30606 34066 30658 34078
rect 31278 34130 31330 34142
rect 31278 34066 31330 34078
rect 31950 34130 32002 34142
rect 36430 34130 36482 34142
rect 33058 34078 33070 34130
rect 33122 34078 33134 34130
rect 31950 34066 32002 34078
rect 36430 34066 36482 34078
rect 36542 34130 36594 34142
rect 36542 34066 36594 34078
rect 37214 34130 37266 34142
rect 37214 34066 37266 34078
rect 42142 34130 42194 34142
rect 42142 34066 42194 34078
rect 25454 34018 25506 34030
rect 32062 34018 32114 34030
rect 43822 34018 43874 34030
rect 10322 33966 10334 34018
rect 10386 33966 10398 34018
rect 24098 33966 24110 34018
rect 24162 33966 24174 34018
rect 26786 33966 26798 34018
rect 26850 33966 26862 34018
rect 29922 33966 29934 34018
rect 29986 33966 29998 34018
rect 33842 33966 33854 34018
rect 33906 33966 33918 34018
rect 35970 33966 35982 34018
rect 36034 33966 36046 34018
rect 42466 33966 42478 34018
rect 42530 33966 42542 34018
rect 25454 33954 25506 33966
rect 32062 33954 32114 33966
rect 43822 33954 43874 33966
rect 37326 33906 37378 33918
rect 37326 33842 37378 33854
rect 37662 33906 37714 33918
rect 37662 33842 37714 33854
rect 42814 33906 42866 33918
rect 42814 33842 42866 33854
rect 1344 33738 44576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 44576 33738
rect 1344 33652 44576 33686
rect 35422 33570 35474 33582
rect 14578 33518 14590 33570
rect 14642 33518 14654 33570
rect 41010 33518 41022 33570
rect 41074 33518 41086 33570
rect 35422 33506 35474 33518
rect 8418 33406 8430 33458
rect 8482 33406 8494 33458
rect 10546 33406 10558 33458
rect 10610 33406 10622 33458
rect 22082 33406 22094 33458
rect 22146 33406 22158 33458
rect 24210 33406 24222 33458
rect 24274 33406 24286 33458
rect 27346 33406 27358 33458
rect 27410 33406 27422 33458
rect 34514 33406 34526 33458
rect 34578 33406 34590 33458
rect 18622 33346 18674 33358
rect 7746 33294 7758 33346
rect 7810 33294 7822 33346
rect 15586 33294 15598 33346
rect 15650 33294 15662 33346
rect 17714 33294 17726 33346
rect 17778 33294 17790 33346
rect 18162 33294 18174 33346
rect 18226 33294 18238 33346
rect 18622 33282 18674 33294
rect 18958 33346 19010 33358
rect 29262 33346 29314 33358
rect 35534 33346 35586 33358
rect 38446 33346 38498 33358
rect 21298 33294 21310 33346
rect 21362 33294 21374 33346
rect 25778 33294 25790 33346
rect 25842 33294 25854 33346
rect 27010 33294 27022 33346
rect 27074 33294 27086 33346
rect 29698 33294 29710 33346
rect 29762 33294 29774 33346
rect 31602 33294 31614 33346
rect 31666 33294 31678 33346
rect 36082 33294 36094 33346
rect 36146 33294 36158 33346
rect 36418 33294 36430 33346
rect 36482 33294 36494 33346
rect 37090 33294 37102 33346
rect 37154 33294 37166 33346
rect 18958 33282 19010 33294
rect 29262 33282 29314 33294
rect 35534 33282 35586 33294
rect 38446 33282 38498 33294
rect 39902 33346 39954 33358
rect 40226 33294 40238 33346
rect 40290 33294 40302 33346
rect 44034 33294 44046 33346
rect 44098 33294 44110 33346
rect 39902 33282 39954 33294
rect 6974 33234 7026 33246
rect 6974 33170 7026 33182
rect 7310 33234 7362 33246
rect 7310 33170 7362 33182
rect 18734 33234 18786 33246
rect 30158 33234 30210 33246
rect 35870 33234 35922 33246
rect 25890 33182 25902 33234
rect 25954 33182 25966 33234
rect 26898 33182 26910 33234
rect 26962 33182 26974 33234
rect 32386 33182 32398 33234
rect 32450 33182 32462 33234
rect 18734 33170 18786 33182
rect 30158 33170 30210 33182
rect 35870 33170 35922 33182
rect 37662 33234 37714 33246
rect 37662 33170 37714 33182
rect 37998 33234 38050 33246
rect 37998 33170 38050 33182
rect 38670 33234 38722 33246
rect 38670 33170 38722 33182
rect 38782 33234 38834 33246
rect 38782 33170 38834 33182
rect 40462 33234 40514 33246
rect 40462 33170 40514 33182
rect 40574 33234 40626 33246
rect 40574 33170 40626 33182
rect 25006 33122 25058 33134
rect 24658 33070 24670 33122
rect 24722 33070 24734 33122
rect 25006 33058 25058 33070
rect 36206 33122 36258 33134
rect 43150 33122 43202 33134
rect 37314 33070 37326 33122
rect 37378 33070 37390 33122
rect 39554 33070 39566 33122
rect 39618 33070 39630 33122
rect 36206 33058 36258 33070
rect 43150 33058 43202 33070
rect 1344 32954 44576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 44576 32954
rect 1344 32868 44576 32902
rect 14702 32786 14754 32798
rect 14018 32734 14030 32786
rect 14082 32734 14094 32786
rect 14702 32722 14754 32734
rect 15934 32786 15986 32798
rect 24670 32786 24722 32798
rect 17938 32734 17950 32786
rect 18002 32734 18014 32786
rect 15934 32722 15986 32734
rect 24670 32722 24722 32734
rect 25790 32786 25842 32798
rect 25790 32722 25842 32734
rect 26126 32786 26178 32798
rect 26126 32722 26178 32734
rect 27694 32786 27746 32798
rect 27694 32722 27746 32734
rect 28030 32786 28082 32798
rect 28030 32722 28082 32734
rect 28926 32786 28978 32798
rect 28926 32722 28978 32734
rect 29598 32786 29650 32798
rect 29598 32722 29650 32734
rect 32398 32786 32450 32798
rect 32398 32722 32450 32734
rect 36878 32786 36930 32798
rect 37998 32786 38050 32798
rect 37650 32734 37662 32786
rect 37714 32734 37726 32786
rect 36878 32722 36930 32734
rect 37998 32722 38050 32734
rect 39678 32786 39730 32798
rect 39678 32722 39730 32734
rect 40350 32786 40402 32798
rect 40350 32722 40402 32734
rect 42926 32786 42978 32798
rect 42926 32722 42978 32734
rect 9550 32674 9602 32686
rect 8194 32622 8206 32674
rect 8258 32622 8270 32674
rect 9550 32610 9602 32622
rect 14926 32674 14978 32686
rect 14926 32610 14978 32622
rect 15598 32674 15650 32686
rect 15598 32610 15650 32622
rect 16158 32674 16210 32686
rect 26350 32674 26402 32686
rect 24322 32622 24334 32674
rect 24386 32622 24398 32674
rect 16158 32610 16210 32622
rect 26350 32610 26402 32622
rect 26910 32674 26962 32686
rect 26910 32610 26962 32622
rect 28478 32674 28530 32686
rect 28478 32610 28530 32622
rect 29038 32674 29090 32686
rect 29038 32610 29090 32622
rect 29374 32674 29426 32686
rect 29374 32610 29426 32622
rect 32510 32674 32562 32686
rect 32510 32610 32562 32622
rect 33854 32674 33906 32686
rect 33854 32610 33906 32622
rect 35982 32674 36034 32686
rect 36430 32674 36482 32686
rect 36194 32622 36206 32674
rect 36258 32622 36270 32674
rect 35982 32610 36034 32622
rect 36430 32610 36482 32622
rect 36766 32674 36818 32686
rect 36766 32610 36818 32622
rect 38782 32674 38834 32686
rect 38782 32610 38834 32622
rect 38894 32674 38946 32686
rect 38894 32610 38946 32622
rect 40014 32674 40066 32686
rect 40014 32610 40066 32622
rect 43374 32674 43426 32686
rect 43374 32610 43426 32622
rect 10446 32562 10498 32574
rect 8866 32510 8878 32562
rect 8930 32510 8942 32562
rect 9986 32510 9998 32562
rect 10050 32510 10062 32562
rect 10446 32498 10498 32510
rect 10894 32562 10946 32574
rect 14590 32562 14642 32574
rect 11554 32510 11566 32562
rect 11618 32510 11630 32562
rect 10894 32498 10946 32510
rect 14590 32498 14642 32510
rect 15038 32562 15090 32574
rect 15038 32498 15090 32510
rect 15486 32562 15538 32574
rect 15486 32498 15538 32510
rect 15822 32562 15874 32574
rect 15822 32498 15874 32510
rect 16270 32562 16322 32574
rect 16270 32498 16322 32510
rect 18286 32562 18338 32574
rect 25902 32562 25954 32574
rect 20178 32510 20190 32562
rect 20242 32510 20254 32562
rect 18286 32498 18338 32510
rect 25902 32498 25954 32510
rect 26686 32562 26738 32574
rect 26686 32498 26738 32510
rect 27022 32562 27074 32574
rect 28814 32562 28866 32574
rect 33182 32562 33234 32574
rect 27234 32510 27246 32562
rect 27298 32510 27310 32562
rect 32162 32510 32174 32562
rect 32226 32510 32238 32562
rect 27022 32498 27074 32510
rect 28814 32498 28866 32510
rect 33182 32498 33234 32510
rect 33518 32562 33570 32574
rect 33518 32498 33570 32510
rect 35198 32562 35250 32574
rect 35198 32498 35250 32510
rect 35646 32562 35698 32574
rect 35646 32498 35698 32510
rect 36318 32562 36370 32574
rect 37438 32562 37490 32574
rect 37090 32510 37102 32562
rect 37154 32510 37166 32562
rect 36318 32498 36370 32510
rect 37438 32498 37490 32510
rect 39118 32562 39170 32574
rect 39118 32498 39170 32510
rect 39342 32562 39394 32574
rect 39342 32498 39394 32510
rect 41022 32562 41074 32574
rect 41022 32498 41074 32510
rect 41358 32562 41410 32574
rect 41358 32498 41410 32510
rect 41806 32562 41858 32574
rect 41806 32498 41858 32510
rect 42030 32562 42082 32574
rect 42030 32498 42082 32510
rect 42478 32562 42530 32574
rect 43586 32510 43598 32562
rect 43650 32510 43662 32562
rect 42478 32498 42530 32510
rect 26014 32450 26066 32462
rect 6066 32398 6078 32450
rect 6130 32398 6142 32450
rect 20850 32398 20862 32450
rect 20914 32398 20926 32450
rect 22978 32398 22990 32450
rect 23042 32398 23054 32450
rect 26014 32386 26066 32398
rect 27918 32450 27970 32462
rect 27918 32386 27970 32398
rect 33406 32450 33458 32462
rect 33406 32386 33458 32398
rect 34974 32450 35026 32462
rect 34974 32386 35026 32398
rect 42254 32450 42306 32462
rect 42254 32386 42306 32398
rect 29710 32338 29762 32350
rect 35534 32338 35586 32350
rect 34626 32286 34638 32338
rect 34690 32286 34702 32338
rect 29710 32274 29762 32286
rect 35534 32274 35586 32286
rect 41134 32338 41186 32350
rect 41134 32274 41186 32286
rect 41470 32338 41522 32350
rect 41470 32274 41522 32286
rect 42702 32338 42754 32350
rect 42702 32274 42754 32286
rect 43038 32338 43090 32350
rect 43038 32274 43090 32286
rect 1344 32170 44576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 44576 32170
rect 1344 32084 44576 32118
rect 26910 32002 26962 32014
rect 31826 31950 31838 32002
rect 31890 31950 31902 32002
rect 39666 31950 39678 32002
rect 39730 31950 39742 32002
rect 26910 31938 26962 31950
rect 7970 31838 7982 31890
rect 8034 31838 8046 31890
rect 10098 31838 10110 31890
rect 10162 31838 10174 31890
rect 17154 31838 17166 31890
rect 17218 31838 17230 31890
rect 31042 31838 31054 31890
rect 31106 31838 31118 31890
rect 33506 31838 33518 31890
rect 33570 31838 33582 31890
rect 35634 31838 35646 31890
rect 35698 31838 35710 31890
rect 37762 31838 37774 31890
rect 37826 31838 37838 31890
rect 11454 31778 11506 31790
rect 23438 31778 23490 31790
rect 39118 31778 39170 31790
rect 7186 31726 7198 31778
rect 7250 31726 7262 31778
rect 13458 31726 13470 31778
rect 13522 31726 13534 31778
rect 14018 31726 14030 31778
rect 14082 31726 14094 31778
rect 16146 31726 16158 31778
rect 16210 31726 16222 31778
rect 23874 31726 23886 31778
rect 23938 31726 23950 31778
rect 27346 31726 27358 31778
rect 27410 31726 27422 31778
rect 28018 31726 28030 31778
rect 28082 31726 28094 31778
rect 31266 31726 31278 31778
rect 31330 31726 31342 31778
rect 32722 31726 32734 31778
rect 32786 31726 32798 31778
rect 11454 31714 11506 31726
rect 23438 31714 23490 31726
rect 39118 31714 39170 31726
rect 39342 31778 39394 31790
rect 39342 31714 39394 31726
rect 40350 31778 40402 31790
rect 44034 31726 44046 31778
rect 44098 31726 44110 31778
rect 40350 31714 40402 31726
rect 37326 31666 37378 31678
rect 38670 31666 38722 31678
rect 17490 31614 17502 31666
rect 17554 31614 17566 31666
rect 27794 31614 27806 31666
rect 27858 31614 27870 31666
rect 37426 31614 37438 31666
rect 37490 31614 37502 31666
rect 37326 31602 37378 31614
rect 38670 31602 38722 31614
rect 38782 31666 38834 31678
rect 38782 31602 38834 31614
rect 40014 31666 40066 31678
rect 40014 31602 40066 31614
rect 40574 31666 40626 31678
rect 40574 31602 40626 31614
rect 41246 31666 41298 31678
rect 41246 31602 41298 31614
rect 11118 31554 11170 31566
rect 11118 31490 11170 31502
rect 17838 31554 17890 31566
rect 17838 31490 17890 31502
rect 18286 31554 18338 31566
rect 32398 31554 32450 31566
rect 26338 31502 26350 31554
rect 26402 31502 26414 31554
rect 27122 31502 27134 31554
rect 27186 31502 27198 31554
rect 18286 31490 18338 31502
rect 32398 31490 32450 31502
rect 36990 31554 37042 31566
rect 36990 31490 37042 31502
rect 37214 31554 37266 31566
rect 37214 31490 37266 31502
rect 38446 31554 38498 31566
rect 38446 31490 38498 31502
rect 40238 31554 40290 31566
rect 40238 31490 40290 31502
rect 41022 31554 41074 31566
rect 41022 31490 41074 31502
rect 41134 31554 41186 31566
rect 41134 31490 41186 31502
rect 43150 31554 43202 31566
rect 43150 31490 43202 31502
rect 1344 31386 44576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 44576 31386
rect 1344 31300 44576 31334
rect 14478 31218 14530 31230
rect 13906 31166 13918 31218
rect 13970 31166 13982 31218
rect 14478 31154 14530 31166
rect 14814 31218 14866 31230
rect 14814 31154 14866 31166
rect 16382 31218 16434 31230
rect 16382 31154 16434 31166
rect 20078 31218 20130 31230
rect 20078 31154 20130 31166
rect 24222 31218 24274 31230
rect 24222 31154 24274 31166
rect 27022 31218 27074 31230
rect 27022 31154 27074 31166
rect 27918 31218 27970 31230
rect 27918 31154 27970 31166
rect 31726 31218 31778 31230
rect 31726 31154 31778 31166
rect 38894 31218 38946 31230
rect 40338 31166 40350 31218
rect 40402 31166 40414 31218
rect 38894 31154 38946 31166
rect 8318 31106 8370 31118
rect 8318 31042 8370 31054
rect 14926 31106 14978 31118
rect 14926 31042 14978 31054
rect 20526 31106 20578 31118
rect 20526 31042 20578 31054
rect 25678 31106 25730 31118
rect 25678 31042 25730 31054
rect 26014 31106 26066 31118
rect 30270 31106 30322 31118
rect 26674 31054 26686 31106
rect 26738 31054 26750 31106
rect 26014 31042 26066 31054
rect 30270 31042 30322 31054
rect 30942 31106 30994 31118
rect 30942 31042 30994 31054
rect 33070 31106 33122 31118
rect 33070 31042 33122 31054
rect 35086 31106 35138 31118
rect 35086 31042 35138 31054
rect 35422 31106 35474 31118
rect 35422 31042 35474 31054
rect 39118 31106 39170 31118
rect 39118 31042 39170 31054
rect 39678 31106 39730 31118
rect 39678 31042 39730 31054
rect 39902 31106 39954 31118
rect 43026 31054 43038 31106
rect 43090 31054 43102 31106
rect 39902 31042 39954 31054
rect 8654 30994 8706 31006
rect 8654 30930 8706 30942
rect 9550 30994 9602 31006
rect 10782 30994 10834 31006
rect 14590 30994 14642 31006
rect 9986 30942 9998 30994
rect 10050 30942 10062 30994
rect 11442 30942 11454 30994
rect 11506 30942 11518 30994
rect 9550 30930 9602 30942
rect 10782 30930 10834 30942
rect 14590 30930 14642 30942
rect 16718 30994 16770 31006
rect 24558 30994 24610 31006
rect 19842 30942 19854 30994
rect 19906 30942 19918 30994
rect 16718 30930 16770 30942
rect 24558 30930 24610 30942
rect 30606 30994 30658 31006
rect 30606 30930 30658 30942
rect 31278 30994 31330 31006
rect 32510 30994 32562 31006
rect 39230 30994 39282 31006
rect 31714 30942 31726 30994
rect 31778 30942 31790 30994
rect 33282 30942 33294 30994
rect 33346 30942 33358 30994
rect 35746 30942 35758 30994
rect 35810 30942 35822 30994
rect 31278 30930 31330 30942
rect 32510 30930 32562 30942
rect 39230 30930 39282 30942
rect 39790 30994 39842 31006
rect 43698 30942 43710 30994
rect 43762 30942 43774 30994
rect 39790 30930 39842 30942
rect 20974 30882 21026 30894
rect 10322 30830 10334 30882
rect 10386 30830 10398 30882
rect 20974 30818 21026 30830
rect 21422 30882 21474 30894
rect 21422 30818 21474 30830
rect 27582 30882 27634 30894
rect 36530 30830 36542 30882
rect 36594 30830 36606 30882
rect 38658 30830 38670 30882
rect 38722 30830 38734 30882
rect 40898 30830 40910 30882
rect 40962 30830 40974 30882
rect 27582 30818 27634 30830
rect 20414 30770 20466 30782
rect 20414 30706 20466 30718
rect 21310 30770 21362 30782
rect 27234 30718 27246 30770
rect 27298 30767 27310 30770
rect 28018 30767 28030 30770
rect 27298 30721 28030 30767
rect 27298 30718 27310 30721
rect 28018 30718 28030 30721
rect 28082 30718 28094 30770
rect 31490 30718 31502 30770
rect 31554 30718 31566 30770
rect 21310 30706 21362 30718
rect 1344 30602 44576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 44576 30602
rect 1344 30516 44576 30550
rect 27022 30434 27074 30446
rect 27022 30370 27074 30382
rect 33742 30434 33794 30446
rect 33742 30370 33794 30382
rect 33406 30322 33458 30334
rect 17042 30270 17054 30322
rect 17106 30270 17118 30322
rect 20738 30270 20750 30322
rect 20802 30270 20814 30322
rect 30482 30270 30494 30322
rect 30546 30270 30558 30322
rect 31938 30270 31950 30322
rect 32002 30270 32014 30322
rect 39330 30270 39342 30322
rect 39394 30270 39406 30322
rect 33406 30258 33458 30270
rect 13806 30210 13858 30222
rect 23550 30210 23602 30222
rect 36990 30210 37042 30222
rect 14242 30158 14254 30210
rect 14306 30158 14318 30210
rect 17826 30158 17838 30210
rect 17890 30158 17902 30210
rect 18610 30158 18622 30210
rect 18674 30158 18686 30210
rect 23986 30158 23998 30210
rect 24050 30158 24062 30210
rect 27458 30158 27470 30210
rect 27522 30158 27534 30210
rect 30594 30158 30606 30210
rect 30658 30158 30670 30210
rect 32274 30158 32286 30210
rect 32338 30158 32350 30210
rect 32946 30158 32958 30210
rect 33010 30158 33022 30210
rect 34290 30158 34302 30210
rect 34354 30158 34366 30210
rect 13806 30146 13858 30158
rect 23550 30146 23602 30158
rect 36990 30146 37042 30158
rect 37214 30210 37266 30222
rect 37214 30146 37266 30158
rect 37550 30210 37602 30222
rect 42590 30210 42642 30222
rect 37986 30158 37998 30210
rect 38050 30158 38062 30210
rect 41458 30158 41470 30210
rect 41522 30158 41534 30210
rect 42130 30158 42142 30210
rect 42194 30158 42206 30210
rect 37550 30146 37602 30158
rect 42590 30146 42642 30158
rect 42814 30210 42866 30222
rect 43474 30158 43486 30210
rect 43538 30158 43550 30210
rect 42814 30146 42866 30158
rect 21646 30098 21698 30110
rect 21646 30034 21698 30046
rect 28142 30098 28194 30110
rect 28142 30034 28194 30046
rect 29598 30098 29650 30110
rect 29598 30034 29650 30046
rect 29934 30098 29986 30110
rect 29934 30034 29986 30046
rect 31278 30098 31330 30110
rect 37102 30098 37154 30110
rect 34066 30046 34078 30098
rect 34130 30046 34142 30098
rect 35074 30046 35086 30098
rect 35138 30046 35150 30098
rect 31278 30034 31330 30046
rect 37102 30034 37154 30046
rect 38222 30098 38274 30110
rect 38222 30034 38274 30046
rect 21310 29986 21362 29998
rect 27806 29986 27858 29998
rect 16482 29934 16494 29986
rect 16546 29934 16558 29986
rect 26450 29934 26462 29986
rect 26514 29934 26526 29986
rect 27234 29934 27246 29986
rect 27298 29934 27310 29986
rect 21310 29922 21362 29934
rect 27806 29922 27858 29934
rect 28030 29986 28082 29998
rect 28030 29922 28082 29934
rect 32734 29986 32786 29998
rect 32734 29922 32786 29934
rect 33630 29986 33682 29998
rect 33630 29922 33682 29934
rect 34750 29986 34802 29998
rect 34750 29922 34802 29934
rect 38782 29986 38834 29998
rect 38782 29922 38834 29934
rect 1344 29818 44576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 44576 29818
rect 1344 29732 44576 29766
rect 13246 29650 13298 29662
rect 13246 29586 13298 29598
rect 15038 29650 15090 29662
rect 15038 29586 15090 29598
rect 16382 29650 16434 29662
rect 16382 29586 16434 29598
rect 24334 29650 24386 29662
rect 24334 29586 24386 29598
rect 25342 29650 25394 29662
rect 30606 29650 30658 29662
rect 29922 29598 29934 29650
rect 29986 29598 29998 29650
rect 25342 29586 25394 29598
rect 30606 29586 30658 29598
rect 34190 29650 34242 29662
rect 34190 29586 34242 29598
rect 15150 29538 15202 29550
rect 8194 29486 8206 29538
rect 8258 29486 8270 29538
rect 15150 29474 15202 29486
rect 16270 29538 16322 29550
rect 16270 29474 16322 29486
rect 17502 29538 17554 29550
rect 17502 29474 17554 29486
rect 18286 29538 18338 29550
rect 23662 29538 23714 29550
rect 28702 29538 28754 29550
rect 33070 29538 33122 29550
rect 40014 29538 40066 29550
rect 20626 29486 20638 29538
rect 20690 29486 20702 29538
rect 26226 29486 26238 29538
rect 26290 29486 26302 29538
rect 27570 29486 27582 29538
rect 27634 29486 27646 29538
rect 27906 29486 27918 29538
rect 27970 29486 27982 29538
rect 32498 29486 32510 29538
rect 32562 29486 32574 29538
rect 35410 29486 35422 29538
rect 35474 29486 35486 29538
rect 41682 29486 41694 29538
rect 41746 29486 41758 29538
rect 18286 29474 18338 29486
rect 23662 29474 23714 29486
rect 28702 29474 28754 29486
rect 33070 29474 33122 29486
rect 40014 29474 40066 29486
rect 17838 29426 17890 29438
rect 23998 29426 24050 29438
rect 8866 29374 8878 29426
rect 8930 29374 8942 29426
rect 9538 29374 9550 29426
rect 9602 29374 9614 29426
rect 10098 29374 10110 29426
rect 10162 29374 10174 29426
rect 12226 29374 12238 29426
rect 12290 29374 12302 29426
rect 19842 29374 19854 29426
rect 19906 29374 19918 29426
rect 17838 29362 17890 29374
rect 23998 29362 24050 29374
rect 24670 29426 24722 29438
rect 24670 29362 24722 29374
rect 25678 29426 25730 29438
rect 27022 29426 27074 29438
rect 26450 29374 26462 29426
rect 26514 29374 26526 29426
rect 25678 29362 25730 29374
rect 27022 29362 27074 29374
rect 27358 29426 27410 29438
rect 27358 29362 27410 29374
rect 28814 29426 28866 29438
rect 28814 29362 28866 29374
rect 29262 29426 29314 29438
rect 30494 29426 30546 29438
rect 29698 29374 29710 29426
rect 29762 29374 29774 29426
rect 30258 29374 30270 29426
rect 30322 29374 30334 29426
rect 29262 29362 29314 29374
rect 30494 29362 30546 29374
rect 30718 29426 30770 29438
rect 30718 29362 30770 29374
rect 30830 29426 30882 29438
rect 31938 29374 31950 29426
rect 32002 29374 32014 29426
rect 33394 29374 33406 29426
rect 33458 29374 33470 29426
rect 34738 29374 34750 29426
rect 34802 29374 34814 29426
rect 40226 29374 40238 29426
rect 40290 29374 40302 29426
rect 40898 29374 40910 29426
rect 40962 29374 40974 29426
rect 30830 29362 30882 29374
rect 13918 29314 13970 29326
rect 6066 29262 6078 29314
rect 6130 29262 6142 29314
rect 13918 29250 13970 29262
rect 16830 29314 16882 29326
rect 33182 29314 33234 29326
rect 22754 29262 22766 29314
rect 22818 29262 22830 29314
rect 16830 29250 16882 29262
rect 33182 29250 33234 29262
rect 33966 29314 34018 29326
rect 33966 29250 34018 29262
rect 34302 29314 34354 29326
rect 37538 29262 37550 29314
rect 37602 29262 37614 29314
rect 43810 29262 43822 29314
rect 43874 29262 43886 29314
rect 34302 29250 34354 29262
rect 14030 29202 14082 29214
rect 14030 29138 14082 29150
rect 16718 29202 16770 29214
rect 16718 29138 16770 29150
rect 18398 29202 18450 29214
rect 18398 29138 18450 29150
rect 28702 29202 28754 29214
rect 28702 29138 28754 29150
rect 32398 29202 32450 29214
rect 32398 29138 32450 29150
rect 1344 29034 44576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 44576 29034
rect 1344 28948 44576 28982
rect 30718 28866 30770 28878
rect 30718 28802 30770 28814
rect 8306 28702 8318 28754
rect 8370 28702 8382 28754
rect 10434 28702 10446 28754
rect 10498 28702 10510 28754
rect 19170 28702 19182 28754
rect 19234 28702 19246 28754
rect 30930 28702 30942 28754
rect 30994 28702 31006 28754
rect 33058 28702 33070 28754
rect 33122 28702 33134 28754
rect 41906 28702 41918 28754
rect 41970 28702 41982 28754
rect 44034 28702 44046 28754
rect 44098 28702 44110 28754
rect 15934 28642 15986 28654
rect 20638 28642 20690 28654
rect 7634 28590 7646 28642
rect 7698 28590 7710 28642
rect 16370 28590 16382 28642
rect 16434 28590 16446 28642
rect 15934 28578 15986 28590
rect 20638 28578 20690 28590
rect 24782 28642 24834 28654
rect 24782 28578 24834 28590
rect 25006 28642 25058 28654
rect 28702 28642 28754 28654
rect 25554 28590 25566 28642
rect 25618 28590 25630 28642
rect 25006 28578 25058 28590
rect 28702 28578 28754 28590
rect 29710 28642 29762 28654
rect 34302 28642 34354 28654
rect 30258 28590 30270 28642
rect 30322 28590 30334 28642
rect 33730 28590 33742 28642
rect 33794 28590 33806 28642
rect 41234 28590 41246 28642
rect 41298 28590 41310 28642
rect 29710 28578 29762 28590
rect 34302 28578 34354 28590
rect 18610 28478 18622 28530
rect 18674 28478 18686 28530
rect 29810 28478 29822 28530
rect 29874 28478 29886 28530
rect 30146 28478 30158 28530
rect 30210 28478 30222 28530
rect 24446 28418 24498 28430
rect 20290 28366 20302 28418
rect 20354 28366 20366 28418
rect 28018 28366 28030 28418
rect 28082 28366 28094 28418
rect 24446 28354 24498 28366
rect 1344 28250 44576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 44576 28250
rect 1344 28164 44576 28198
rect 13022 28082 13074 28094
rect 13022 28018 13074 28030
rect 24670 28082 24722 28094
rect 24670 28018 24722 28030
rect 26014 28082 26066 28094
rect 26014 28018 26066 28030
rect 28030 28082 28082 28094
rect 28030 28018 28082 28030
rect 28254 28082 28306 28094
rect 28254 28018 28306 28030
rect 17390 27970 17442 27982
rect 13794 27918 13806 27970
rect 13858 27918 13870 27970
rect 17390 27906 17442 27918
rect 17502 27970 17554 27982
rect 17502 27906 17554 27918
rect 18174 27970 18226 27982
rect 25230 27970 25282 27982
rect 21410 27918 21422 27970
rect 21474 27918 21486 27970
rect 18174 27906 18226 27918
rect 25230 27906 25282 27918
rect 25902 27970 25954 27982
rect 28366 27970 28418 27982
rect 27458 27918 27470 27970
rect 27522 27918 27534 27970
rect 25902 27906 25954 27918
rect 28366 27906 28418 27918
rect 29150 27970 29202 27982
rect 43810 27918 43822 27970
rect 43874 27918 43886 27970
rect 29150 27906 29202 27918
rect 18734 27858 18786 27870
rect 25566 27858 25618 27870
rect 10994 27806 11006 27858
rect 11058 27806 11070 27858
rect 16034 27806 16046 27858
rect 16098 27806 16110 27858
rect 16594 27806 16606 27858
rect 16658 27806 16670 27858
rect 19170 27806 19182 27858
rect 19234 27806 19246 27858
rect 24434 27806 24446 27858
rect 24498 27806 24510 27858
rect 18734 27794 18786 27806
rect 25566 27794 25618 27806
rect 26574 27858 26626 27870
rect 26574 27794 26626 27806
rect 26910 27858 26962 27870
rect 44158 27858 44210 27870
rect 27346 27806 27358 27858
rect 27410 27806 27422 27858
rect 29586 27806 29598 27858
rect 29650 27806 29662 27858
rect 26910 27794 26962 27806
rect 44158 27794 44210 27806
rect 11566 27746 11618 27758
rect 11106 27694 11118 27746
rect 11170 27694 11182 27746
rect 11566 27682 11618 27694
rect 12014 27746 12066 27758
rect 23998 27746 24050 27758
rect 21970 27694 21982 27746
rect 22034 27694 22046 27746
rect 12014 27682 12066 27694
rect 23998 27682 24050 27694
rect 29262 27746 29314 27758
rect 43150 27746 43202 27758
rect 30370 27694 30382 27746
rect 30434 27694 30446 27746
rect 32498 27694 32510 27746
rect 32562 27694 32574 27746
rect 29262 27682 29314 27694
rect 43150 27682 43202 27694
rect 43598 27746 43650 27758
rect 43598 27682 43650 27694
rect 11902 27634 11954 27646
rect 11902 27570 11954 27582
rect 18286 27634 18338 27646
rect 18286 27570 18338 27582
rect 26014 27634 26066 27646
rect 26014 27570 26066 27582
rect 1344 27466 44576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 44576 27466
rect 1344 27380 44576 27414
rect 15822 27298 15874 27310
rect 15822 27234 15874 27246
rect 20190 27298 20242 27310
rect 20190 27234 20242 27246
rect 21422 27298 21474 27310
rect 21422 27234 21474 27246
rect 27806 27298 27858 27310
rect 27806 27234 27858 27246
rect 9214 27186 9266 27198
rect 20302 27186 20354 27198
rect 35086 27186 35138 27198
rect 19618 27134 19630 27186
rect 19682 27134 19694 27186
rect 29586 27134 29598 27186
rect 29650 27134 29662 27186
rect 9214 27122 9266 27134
rect 20302 27122 20354 27134
rect 35086 27122 35138 27134
rect 37102 27186 37154 27198
rect 44146 27134 44158 27186
rect 44210 27134 44222 27186
rect 37102 27122 37154 27134
rect 9662 27074 9714 27086
rect 11006 27074 11058 27086
rect 16270 27074 16322 27086
rect 24334 27074 24386 27086
rect 10098 27022 10110 27074
rect 10162 27022 10174 27074
rect 11218 27022 11230 27074
rect 11282 27022 11294 27074
rect 12450 27022 12462 27074
rect 12514 27022 12526 27074
rect 16594 27022 16606 27074
rect 16658 27022 16670 27074
rect 24770 27022 24782 27074
rect 24834 27022 24846 27074
rect 32386 27022 32398 27074
rect 32450 27022 32462 27074
rect 41010 27022 41022 27074
rect 41074 27022 41086 27074
rect 41794 27022 41806 27074
rect 41858 27022 41870 27074
rect 9662 27010 9714 27022
rect 11006 27010 11058 27022
rect 16270 27010 16322 27022
rect 24334 27010 24386 27022
rect 10558 26962 10610 26974
rect 10558 26898 10610 26910
rect 11902 26962 11954 26974
rect 11902 26898 11954 26910
rect 12238 26962 12290 26974
rect 12238 26898 12290 26910
rect 15374 26962 15426 26974
rect 15374 26898 15426 26910
rect 15710 26962 15762 26974
rect 21310 26962 21362 26974
rect 18946 26910 18958 26962
rect 19010 26910 19022 26962
rect 15710 26898 15762 26910
rect 21310 26898 21362 26910
rect 27022 26962 27074 26974
rect 34750 26962 34802 26974
rect 31714 26910 31726 26962
rect 31778 26910 31790 26962
rect 27022 26898 27074 26910
rect 34750 26898 34802 26910
rect 35646 26962 35698 26974
rect 35646 26898 35698 26910
rect 36094 26962 36146 26974
rect 36094 26898 36146 26910
rect 38558 26962 38610 26974
rect 38558 26898 38610 26910
rect 39230 26962 39282 26974
rect 39230 26898 39282 26910
rect 40798 26962 40850 26974
rect 40798 26898 40850 26910
rect 35982 26850 36034 26862
rect 35982 26786 36034 26798
rect 38222 26850 38274 26862
rect 38222 26786 38274 26798
rect 38894 26850 38946 26862
rect 38894 26786 38946 26798
rect 1344 26682 44576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 44576 26682
rect 1344 26596 44576 26630
rect 13918 26514 13970 26526
rect 13122 26462 13134 26514
rect 13186 26462 13198 26514
rect 13918 26450 13970 26462
rect 19070 26514 19122 26526
rect 19070 26450 19122 26462
rect 25902 26514 25954 26526
rect 25902 26450 25954 26462
rect 30942 26514 30994 26526
rect 30942 26450 30994 26462
rect 34190 26514 34242 26526
rect 37538 26462 37550 26514
rect 37602 26462 37614 26514
rect 44146 26462 44158 26514
rect 44210 26462 44222 26514
rect 34190 26450 34242 26462
rect 30830 26402 30882 26414
rect 23538 26350 23550 26402
rect 23602 26350 23614 26402
rect 26562 26350 26574 26402
rect 26626 26350 26638 26402
rect 27010 26350 27022 26402
rect 27074 26350 27086 26402
rect 30830 26338 30882 26350
rect 8990 26290 9042 26302
rect 16830 26290 16882 26302
rect 20862 26290 20914 26302
rect 26238 26290 26290 26302
rect 8530 26238 8542 26290
rect 8594 26238 8606 26290
rect 10098 26238 10110 26290
rect 10162 26238 10174 26290
rect 10658 26238 10670 26290
rect 10722 26238 10734 26290
rect 14130 26238 14142 26290
rect 14194 26238 14206 26290
rect 19282 26238 19294 26290
rect 19346 26238 19358 26290
rect 21298 26238 21310 26290
rect 21362 26238 21374 26290
rect 8990 26226 9042 26238
rect 16830 26226 16882 26238
rect 20862 26226 20914 26238
rect 26238 26226 26290 26238
rect 34638 26290 34690 26302
rect 34962 26238 34974 26290
rect 35026 26238 35038 26290
rect 39442 26238 39454 26290
rect 39506 26238 39518 26290
rect 41010 26238 41022 26290
rect 41074 26238 41086 26290
rect 41794 26238 41806 26290
rect 41858 26238 41870 26290
rect 34638 26226 34690 26238
rect 9662 26178 9714 26190
rect 17502 26178 17554 26190
rect 13458 26126 13470 26178
rect 13522 26126 13534 26178
rect 9662 26114 9714 26126
rect 17502 26114 17554 26126
rect 19854 26178 19906 26190
rect 19854 26114 19906 26126
rect 20302 26178 20354 26190
rect 27582 26178 27634 26190
rect 24098 26126 24110 26178
rect 24162 26126 24174 26178
rect 20302 26114 20354 26126
rect 27582 26114 27634 26126
rect 34078 26178 34130 26190
rect 37874 26126 37886 26178
rect 37938 26126 37950 26178
rect 38882 26126 38894 26178
rect 38946 26126 38958 26178
rect 34078 26114 34130 26126
rect 9774 26066 9826 26078
rect 9774 26002 9826 26014
rect 17390 26066 17442 26078
rect 17390 26002 17442 26014
rect 19742 26066 19794 26078
rect 39218 26014 39230 26066
rect 39282 26014 39294 26066
rect 19742 26002 19794 26014
rect 1344 25898 44576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 44576 25898
rect 1344 25812 44576 25846
rect 19742 25730 19794 25742
rect 19742 25666 19794 25678
rect 22542 25730 22594 25742
rect 22542 25666 22594 25678
rect 23998 25730 24050 25742
rect 37538 25678 37550 25730
rect 37602 25678 37614 25730
rect 38658 25678 38670 25730
rect 38722 25678 38734 25730
rect 23998 25666 24050 25678
rect 8318 25618 8370 25630
rect 21422 25618 21474 25630
rect 9538 25566 9550 25618
rect 9602 25566 9614 25618
rect 8318 25554 8370 25566
rect 21422 25554 21474 25566
rect 22430 25618 22482 25630
rect 22430 25554 22482 25566
rect 24110 25618 24162 25630
rect 24110 25554 24162 25566
rect 28030 25618 28082 25630
rect 41470 25618 41522 25630
rect 37874 25566 37886 25618
rect 37938 25566 37950 25618
rect 28030 25554 28082 25566
rect 41470 25554 41522 25566
rect 7310 25506 7362 25518
rect 7310 25442 7362 25454
rect 7870 25506 7922 25518
rect 12798 25506 12850 25518
rect 26350 25506 26402 25518
rect 12338 25454 12350 25506
rect 12402 25454 12414 25506
rect 16146 25454 16158 25506
rect 16210 25454 16222 25506
rect 16706 25454 16718 25506
rect 16770 25454 16782 25506
rect 25666 25454 25678 25506
rect 25730 25454 25742 25506
rect 7870 25442 7922 25454
rect 12798 25442 12850 25454
rect 26350 25442 26402 25454
rect 33070 25506 33122 25518
rect 38782 25506 38834 25518
rect 33506 25454 33518 25506
rect 33570 25454 33582 25506
rect 37426 25454 37438 25506
rect 37490 25454 37502 25506
rect 39442 25454 39454 25506
rect 39506 25454 39518 25506
rect 33070 25442 33122 25454
rect 38782 25442 38834 25454
rect 15710 25394 15762 25406
rect 42254 25394 42306 25406
rect 10098 25342 10110 25394
rect 10162 25342 10174 25394
rect 19954 25342 19966 25394
rect 20018 25342 20030 25394
rect 25106 25342 25118 25394
rect 25170 25342 25182 25394
rect 15710 25330 15762 25342
rect 42254 25330 42306 25342
rect 15822 25282 15874 25294
rect 20302 25282 20354 25294
rect 19170 25230 19182 25282
rect 19234 25230 19246 25282
rect 15822 25218 15874 25230
rect 20302 25218 20354 25230
rect 21310 25282 21362 25294
rect 28590 25282 28642 25294
rect 25442 25230 25454 25282
rect 25506 25230 25518 25282
rect 21310 25218 21362 25230
rect 28590 25218 28642 25230
rect 29262 25282 29314 25294
rect 36542 25282 36594 25294
rect 35858 25230 35870 25282
rect 35922 25230 35934 25282
rect 29262 25218 29314 25230
rect 36542 25218 36594 25230
rect 41358 25282 41410 25294
rect 41358 25218 41410 25230
rect 41918 25282 41970 25294
rect 41918 25218 41970 25230
rect 44158 25282 44210 25294
rect 44158 25218 44210 25230
rect 1344 25114 44576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 44576 25114
rect 1344 25028 44576 25062
rect 6974 24946 7026 24958
rect 6974 24882 7026 24894
rect 7758 24946 7810 24958
rect 7758 24882 7810 24894
rect 10334 24946 10386 24958
rect 21982 24946 22034 24958
rect 10882 24894 10894 24946
rect 10946 24894 10958 24946
rect 21298 24894 21310 24946
rect 21362 24894 21374 24946
rect 37986 24894 37998 24946
rect 38050 24894 38062 24946
rect 10334 24882 10386 24894
rect 21982 24882 22034 24894
rect 17950 24834 18002 24846
rect 17950 24770 18002 24782
rect 22542 24834 22594 24846
rect 22542 24770 22594 24782
rect 25230 24834 25282 24846
rect 27806 24834 27858 24846
rect 27234 24782 27246 24834
rect 27298 24782 27310 24834
rect 25230 24770 25282 24782
rect 27806 24770 27858 24782
rect 43038 24834 43090 24846
rect 43038 24770 43090 24782
rect 8094 24722 8146 24734
rect 13806 24722 13858 24734
rect 13346 24670 13358 24722
rect 13410 24670 13422 24722
rect 8094 24658 8146 24670
rect 13806 24658 13858 24670
rect 18062 24722 18114 24734
rect 18062 24658 18114 24670
rect 18510 24722 18562 24734
rect 25566 24722 25618 24734
rect 18834 24670 18846 24722
rect 18898 24670 18910 24722
rect 18510 24658 18562 24670
rect 25566 24658 25618 24670
rect 26126 24722 26178 24734
rect 35086 24722 35138 24734
rect 42702 24722 42754 24734
rect 27122 24670 27134 24722
rect 27186 24670 27198 24722
rect 29026 24670 29038 24722
rect 29090 24670 29102 24722
rect 34066 24670 34078 24722
rect 34130 24670 34142 24722
rect 35522 24670 35534 24722
rect 35586 24670 35598 24722
rect 41458 24670 41470 24722
rect 41522 24670 41534 24722
rect 26126 24658 26178 24670
rect 35086 24658 35138 24670
rect 42702 24658 42754 24670
rect 7198 24610 7250 24622
rect 7198 24546 7250 24558
rect 8654 24610 8706 24622
rect 8654 24546 8706 24558
rect 26462 24610 26514 24622
rect 32174 24610 32226 24622
rect 34638 24610 34690 24622
rect 42254 24610 42306 24622
rect 29698 24558 29710 24610
rect 29762 24558 29774 24610
rect 31826 24558 31838 24610
rect 31890 24558 31902 24610
rect 33730 24558 33742 24610
rect 33794 24558 33806 24610
rect 38322 24558 38334 24610
rect 38386 24558 38398 24610
rect 41682 24558 41694 24610
rect 41746 24558 41758 24610
rect 26462 24546 26514 24558
rect 32174 24546 32226 24558
rect 34638 24546 34690 24558
rect 42254 24546 42306 24558
rect 22430 24498 22482 24510
rect 22430 24434 22482 24446
rect 32286 24498 32338 24510
rect 32286 24434 32338 24446
rect 1344 24330 44576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 44576 24330
rect 1344 24244 44576 24278
rect 19406 24162 19458 24174
rect 19406 24098 19458 24110
rect 19742 24162 19794 24174
rect 19742 24098 19794 24110
rect 29262 24050 29314 24062
rect 33294 24050 33346 24062
rect 8754 23998 8766 24050
rect 8818 23998 8830 24050
rect 15474 23998 15486 24050
rect 15538 23998 15550 24050
rect 24770 23998 24782 24050
rect 24834 23998 24846 24050
rect 26898 23998 26910 24050
rect 26962 23998 26974 24050
rect 32946 23998 32958 24050
rect 33010 23998 33022 24050
rect 44034 23998 44046 24050
rect 44098 23998 44110 24050
rect 29262 23986 29314 23998
rect 33294 23986 33346 23998
rect 7758 23938 7810 23950
rect 12462 23938 12514 23950
rect 29486 23938 29538 23950
rect 7186 23886 7198 23938
rect 7250 23886 7262 23938
rect 8530 23886 8542 23938
rect 8594 23886 8606 23938
rect 18274 23886 18286 23938
rect 18338 23886 18350 23938
rect 18834 23886 18846 23938
rect 18898 23886 18910 23938
rect 24098 23886 24110 23938
rect 24162 23886 24174 23938
rect 7758 23874 7810 23886
rect 12462 23874 12514 23886
rect 29486 23874 29538 23886
rect 29598 23938 29650 23950
rect 35198 23938 35250 23950
rect 30034 23886 30046 23938
rect 30098 23886 30110 23938
rect 34962 23886 34974 23938
rect 35026 23886 35038 23938
rect 29598 23874 29650 23886
rect 35198 23874 35250 23886
rect 35422 23938 35474 23950
rect 35422 23874 35474 23886
rect 37550 23938 37602 23950
rect 40674 23886 40686 23938
rect 40738 23886 40750 23938
rect 41234 23886 41246 23938
rect 41298 23886 41310 23938
rect 37550 23874 37602 23886
rect 7870 23826 7922 23838
rect 7870 23762 7922 23774
rect 9214 23826 9266 23838
rect 9214 23762 9266 23774
rect 9550 23826 9602 23838
rect 9550 23762 9602 23774
rect 9886 23826 9938 23838
rect 19294 23826 19346 23838
rect 16034 23774 16046 23826
rect 16098 23774 16110 23826
rect 9886 23762 9938 23774
rect 19294 23762 19346 23774
rect 19854 23826 19906 23838
rect 19854 23762 19906 23774
rect 29150 23826 29202 23838
rect 36318 23826 36370 23838
rect 30818 23774 30830 23826
rect 30882 23774 30894 23826
rect 29150 23762 29202 23774
rect 36318 23762 36370 23774
rect 37214 23826 37266 23838
rect 43474 23774 43486 23826
rect 43538 23774 43550 23826
rect 37214 23762 37266 23774
rect 6526 23714 6578 23726
rect 6178 23662 6190 23714
rect 6242 23662 6254 23714
rect 6526 23650 6578 23662
rect 12798 23714 12850 23726
rect 12798 23650 12850 23662
rect 20302 23714 20354 23726
rect 20302 23650 20354 23662
rect 28142 23714 28194 23726
rect 28142 23650 28194 23662
rect 33406 23714 33458 23726
rect 33406 23650 33458 23662
rect 35310 23714 35362 23726
rect 35310 23650 35362 23662
rect 35534 23714 35586 23726
rect 35534 23650 35586 23662
rect 36206 23714 36258 23726
rect 36206 23650 36258 23662
rect 1344 23546 44576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 44576 23546
rect 1344 23460 44576 23494
rect 21534 23378 21586 23390
rect 13570 23326 13582 23378
rect 13634 23326 13646 23378
rect 21534 23314 21586 23326
rect 30830 23378 30882 23390
rect 30830 23314 30882 23326
rect 31614 23378 31666 23390
rect 31614 23314 31666 23326
rect 35534 23378 35586 23390
rect 35534 23314 35586 23326
rect 39790 23378 39842 23390
rect 39790 23314 39842 23326
rect 8654 23266 8706 23278
rect 8654 23202 8706 23214
rect 20190 23266 20242 23278
rect 20190 23202 20242 23214
rect 20862 23266 20914 23278
rect 20862 23202 20914 23214
rect 21198 23266 21250 23278
rect 21198 23202 21250 23214
rect 31054 23266 31106 23278
rect 31054 23202 31106 23214
rect 35086 23266 35138 23278
rect 35086 23202 35138 23214
rect 36542 23266 36594 23278
rect 36542 23202 36594 23214
rect 36990 23266 37042 23278
rect 36990 23202 37042 23214
rect 37886 23266 37938 23278
rect 37886 23202 37938 23214
rect 42478 23266 42530 23278
rect 42478 23202 42530 23214
rect 43822 23266 43874 23278
rect 43822 23202 43874 23214
rect 6414 23154 6466 23166
rect 7758 23154 7810 23166
rect 6066 23102 6078 23154
rect 6130 23102 6142 23154
rect 7186 23102 7198 23154
rect 7250 23102 7262 23154
rect 6414 23090 6466 23102
rect 7758 23090 7810 23102
rect 7870 23154 7922 23166
rect 7870 23090 7922 23102
rect 8318 23154 8370 23166
rect 17838 23154 17890 23166
rect 19518 23154 19570 23166
rect 10770 23102 10782 23154
rect 10834 23102 10846 23154
rect 11218 23102 11230 23154
rect 11282 23102 11294 23154
rect 18386 23102 18398 23154
rect 18450 23102 18462 23154
rect 19170 23102 19182 23154
rect 19234 23102 19246 23154
rect 8318 23090 8370 23102
rect 17838 23090 17890 23102
rect 19518 23090 19570 23102
rect 20526 23154 20578 23166
rect 28702 23154 28754 23166
rect 21746 23102 21758 23154
rect 21810 23102 21822 23154
rect 25330 23102 25342 23154
rect 25394 23102 25406 23154
rect 28466 23102 28478 23154
rect 28530 23102 28542 23154
rect 20526 23090 20578 23102
rect 28702 23090 28754 23102
rect 28926 23154 28978 23166
rect 28926 23090 28978 23102
rect 29038 23154 29090 23166
rect 30606 23154 30658 23166
rect 30370 23102 30382 23154
rect 30434 23102 30446 23154
rect 29038 23090 29090 23102
rect 30606 23090 30658 23102
rect 31166 23154 31218 23166
rect 32398 23154 32450 23166
rect 35982 23154 36034 23166
rect 36766 23154 36818 23166
rect 31826 23102 31838 23154
rect 31890 23102 31902 23154
rect 35298 23102 35310 23154
rect 35362 23102 35374 23154
rect 36306 23102 36318 23154
rect 36370 23102 36382 23154
rect 31166 23090 31218 23102
rect 32398 23090 32450 23102
rect 35982 23090 36034 23102
rect 36766 23090 36818 23102
rect 37774 23154 37826 23166
rect 42814 23154 42866 23166
rect 44158 23154 44210 23166
rect 38882 23102 38894 23154
rect 38946 23102 38958 23154
rect 41570 23102 41582 23154
rect 41634 23102 41646 23154
rect 43250 23102 43262 23154
rect 43314 23102 43326 23154
rect 37774 23090 37826 23102
rect 42814 23090 42866 23102
rect 44158 23090 44210 23102
rect 5518 23042 5570 23054
rect 28814 23042 28866 23054
rect 14130 22990 14142 23042
rect 14194 22990 14206 23042
rect 26002 22990 26014 23042
rect 26066 22990 26078 23042
rect 28130 22990 28142 23042
rect 28194 22990 28206 23042
rect 5518 22978 5570 22990
rect 28814 22978 28866 22990
rect 29710 23042 29762 23054
rect 38446 23042 38498 23054
rect 34962 22990 34974 23042
rect 35026 22990 35038 23042
rect 36418 22990 36430 23042
rect 36482 22990 36494 23042
rect 29710 22978 29762 22990
rect 38446 22978 38498 22990
rect 40350 23042 40402 23054
rect 41682 22990 41694 23042
rect 41746 22990 41758 23042
rect 40350 22978 40402 22990
rect 30046 22930 30098 22942
rect 18498 22878 18510 22930
rect 18562 22878 18574 22930
rect 30046 22866 30098 22878
rect 30382 22930 30434 22942
rect 30382 22866 30434 22878
rect 35870 22930 35922 22942
rect 35870 22866 35922 22878
rect 1344 22762 44576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 44576 22762
rect 1344 22676 44576 22710
rect 10446 22594 10498 22606
rect 10446 22530 10498 22542
rect 11790 22594 11842 22606
rect 34974 22594 35026 22606
rect 18834 22542 18846 22594
rect 18898 22591 18910 22594
rect 19282 22591 19294 22594
rect 18898 22545 19294 22591
rect 18898 22542 18910 22545
rect 19282 22542 19294 22545
rect 19346 22542 19358 22594
rect 11790 22530 11842 22542
rect 34974 22530 35026 22542
rect 38558 22594 38610 22606
rect 38558 22530 38610 22542
rect 19294 22482 19346 22494
rect 12786 22430 12798 22482
rect 12850 22430 12862 22482
rect 15250 22430 15262 22482
rect 15314 22430 15326 22482
rect 19294 22418 19346 22430
rect 23998 22482 24050 22494
rect 23998 22418 24050 22430
rect 29598 22482 29650 22494
rect 33966 22482 34018 22494
rect 44270 22482 44322 22494
rect 33058 22430 33070 22482
rect 33122 22430 33134 22482
rect 42354 22430 42366 22482
rect 42418 22430 42430 22482
rect 29598 22418 29650 22430
rect 33966 22418 34018 22430
rect 44270 22418 44322 22430
rect 5966 22370 6018 22382
rect 4834 22318 4846 22370
rect 4898 22318 4910 22370
rect 5966 22306 6018 22318
rect 6526 22370 6578 22382
rect 6526 22306 6578 22318
rect 6974 22370 7026 22382
rect 12350 22370 12402 22382
rect 7410 22318 7422 22370
rect 7474 22318 7486 22370
rect 10882 22318 10894 22370
rect 10946 22318 10958 22370
rect 6974 22306 7026 22318
rect 12350 22306 12402 22318
rect 12686 22370 12738 22382
rect 12686 22306 12738 22318
rect 13582 22370 13634 22382
rect 21758 22370 21810 22382
rect 26686 22370 26738 22382
rect 28254 22370 28306 22382
rect 33742 22370 33794 22382
rect 18162 22318 18174 22370
rect 18226 22318 18238 22370
rect 20402 22318 20414 22370
rect 20466 22318 20478 22370
rect 23762 22318 23774 22370
rect 23826 22318 23838 22370
rect 25554 22318 25566 22370
rect 25618 22318 25630 22370
rect 27122 22318 27134 22370
rect 27186 22318 27198 22370
rect 30258 22318 30270 22370
rect 30322 22318 30334 22370
rect 13582 22306 13634 22318
rect 21758 22306 21810 22318
rect 26686 22306 26738 22318
rect 28254 22306 28306 22318
rect 33742 22306 33794 22318
rect 34190 22370 34242 22382
rect 34190 22306 34242 22318
rect 35198 22370 35250 22382
rect 35198 22306 35250 22318
rect 35422 22370 35474 22382
rect 37438 22370 37490 22382
rect 35634 22318 35646 22370
rect 35698 22318 35710 22370
rect 36978 22318 36990 22370
rect 37042 22318 37054 22370
rect 35422 22306 35474 22318
rect 37438 22306 37490 22318
rect 39118 22370 39170 22382
rect 39442 22318 39454 22370
rect 39506 22318 39518 22370
rect 39118 22306 39170 22318
rect 11678 22258 11730 22270
rect 9650 22206 9662 22258
rect 9714 22206 9726 22258
rect 11678 22194 11730 22206
rect 12462 22258 12514 22270
rect 12462 22194 12514 22206
rect 12798 22258 12850 22270
rect 24110 22258 24162 22270
rect 17378 22206 17390 22258
rect 17442 22206 17454 22258
rect 22082 22206 22094 22258
rect 22146 22206 22158 22258
rect 22530 22206 22542 22258
rect 22594 22206 22606 22258
rect 12798 22194 12850 22206
rect 24110 22194 24162 22206
rect 25790 22258 25842 22270
rect 28590 22258 28642 22270
rect 27458 22206 27470 22258
rect 27522 22206 27534 22258
rect 25790 22194 25842 22206
rect 28590 22194 28642 22206
rect 29486 22258 29538 22270
rect 34414 22258 34466 22270
rect 30930 22206 30942 22258
rect 30994 22206 31006 22258
rect 29486 22194 29538 22206
rect 34414 22194 34466 22206
rect 37214 22258 37266 22270
rect 37214 22194 37266 22206
rect 38670 22258 38722 22270
rect 38670 22194 38722 22206
rect 5070 22146 5122 22158
rect 5070 22082 5122 22094
rect 10670 22146 10722 22158
rect 10670 22082 10722 22094
rect 13694 22146 13746 22158
rect 13694 22082 13746 22094
rect 13806 22146 13858 22158
rect 13806 22082 13858 22094
rect 13918 22146 13970 22158
rect 13918 22082 13970 22094
rect 14030 22146 14082 22158
rect 14030 22082 14082 22094
rect 19742 22146 19794 22158
rect 19742 22082 19794 22094
rect 20190 22146 20242 22158
rect 20190 22082 20242 22094
rect 21422 22146 21474 22158
rect 21422 22082 21474 22094
rect 23102 22146 23154 22158
rect 23102 22082 23154 22094
rect 26350 22146 26402 22158
rect 26350 22082 26402 22094
rect 29710 22146 29762 22158
rect 29710 22082 29762 22094
rect 34302 22146 34354 22158
rect 34302 22082 34354 22094
rect 35086 22146 35138 22158
rect 35086 22082 35138 22094
rect 37326 22146 37378 22158
rect 37326 22082 37378 22094
rect 37550 22146 37602 22158
rect 41906 22094 41918 22146
rect 41970 22094 41982 22146
rect 37550 22082 37602 22094
rect 1344 21978 44576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 44576 21978
rect 1344 21892 44576 21926
rect 11006 21810 11058 21822
rect 11006 21746 11058 21758
rect 12910 21810 12962 21822
rect 12910 21746 12962 21758
rect 15486 21810 15538 21822
rect 15486 21746 15538 21758
rect 17502 21810 17554 21822
rect 17502 21746 17554 21758
rect 18846 21810 18898 21822
rect 18846 21746 18898 21758
rect 30942 21810 30994 21822
rect 30942 21746 30994 21758
rect 36094 21810 36146 21822
rect 36094 21746 36146 21758
rect 39790 21810 39842 21822
rect 39790 21746 39842 21758
rect 7646 21698 7698 21710
rect 6626 21646 6638 21698
rect 6690 21646 6702 21698
rect 7646 21634 7698 21646
rect 10558 21698 10610 21710
rect 10558 21634 10610 21646
rect 14478 21698 14530 21710
rect 14478 21634 14530 21646
rect 15822 21698 15874 21710
rect 15822 21634 15874 21646
rect 15934 21698 15986 21710
rect 15934 21634 15986 21646
rect 16494 21698 16546 21710
rect 16494 21634 16546 21646
rect 17726 21698 17778 21710
rect 17726 21634 17778 21646
rect 19630 21698 19682 21710
rect 19630 21634 19682 21646
rect 28590 21698 28642 21710
rect 28590 21634 28642 21646
rect 34414 21698 34466 21710
rect 34414 21634 34466 21646
rect 34974 21698 35026 21710
rect 34974 21634 35026 21646
rect 36542 21698 36594 21710
rect 36542 21634 36594 21646
rect 3950 21586 4002 21598
rect 7758 21586 7810 21598
rect 4386 21534 4398 21586
rect 4450 21534 4462 21586
rect 3950 21522 4002 21534
rect 7758 21522 7810 21534
rect 11342 21586 11394 21598
rect 11342 21522 11394 21534
rect 11566 21586 11618 21598
rect 11566 21522 11618 21534
rect 11790 21586 11842 21598
rect 11790 21522 11842 21534
rect 12014 21586 12066 21598
rect 13358 21586 13410 21598
rect 13122 21534 13134 21586
rect 13186 21534 13198 21586
rect 12014 21522 12066 21534
rect 13358 21522 13410 21534
rect 14142 21586 14194 21598
rect 14142 21522 14194 21534
rect 14254 21586 14306 21598
rect 16382 21586 16434 21598
rect 14690 21534 14702 21586
rect 14754 21534 14766 21586
rect 14254 21522 14306 21534
rect 16382 21522 16434 21534
rect 16942 21586 16994 21598
rect 16942 21522 16994 21534
rect 17278 21586 17330 21598
rect 17278 21522 17330 21534
rect 17950 21586 18002 21598
rect 17950 21522 18002 21534
rect 18734 21586 18786 21598
rect 28478 21586 28530 21598
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 19954 21534 19966 21586
rect 20018 21534 20030 21586
rect 25330 21534 25342 21586
rect 25394 21534 25406 21586
rect 18734 21522 18786 21534
rect 28478 21522 28530 21534
rect 29150 21586 29202 21598
rect 29150 21522 29202 21534
rect 31278 21586 31330 21598
rect 31278 21522 31330 21534
rect 31726 21586 31778 21598
rect 31726 21522 31778 21534
rect 33966 21586 34018 21598
rect 33966 21522 34018 21534
rect 34190 21586 34242 21598
rect 34190 21522 34242 21534
rect 34638 21586 34690 21598
rect 34638 21522 34690 21534
rect 35422 21586 35474 21598
rect 35422 21522 35474 21534
rect 36430 21586 36482 21598
rect 36430 21522 36482 21534
rect 36654 21586 36706 21598
rect 36654 21522 36706 21534
rect 36878 21586 36930 21598
rect 36878 21522 36930 21534
rect 37102 21586 37154 21598
rect 41906 21534 41918 21586
rect 41970 21534 41982 21586
rect 37102 21522 37154 21534
rect 10894 21474 10946 21486
rect 7186 21422 7198 21474
rect 7250 21422 7262 21474
rect 10894 21410 10946 21422
rect 11902 21474 11954 21486
rect 14366 21474 14418 21486
rect 13458 21422 13470 21474
rect 13522 21422 13534 21474
rect 11902 21410 11954 21422
rect 14366 21410 14418 21422
rect 15374 21474 15426 21486
rect 15374 21410 15426 21422
rect 16718 21474 16770 21486
rect 29598 21474 29650 21486
rect 20738 21422 20750 21474
rect 20802 21422 20814 21474
rect 22866 21422 22878 21474
rect 22930 21422 22942 21474
rect 26002 21422 26014 21474
rect 26066 21422 26078 21474
rect 28130 21422 28142 21474
rect 28194 21422 28206 21474
rect 40226 21422 40238 21474
rect 40290 21422 40302 21474
rect 41682 21422 41694 21474
rect 41746 21422 41758 21474
rect 16718 21410 16770 21422
rect 29598 21410 29650 21422
rect 10446 21362 10498 21374
rect 10446 21298 10498 21310
rect 12462 21362 12514 21374
rect 12462 21298 12514 21310
rect 12574 21362 12626 21374
rect 12574 21298 12626 21310
rect 18622 21362 18674 21374
rect 18622 21298 18674 21310
rect 28590 21362 28642 21374
rect 34078 21362 34130 21374
rect 29138 21310 29150 21362
rect 29202 21359 29214 21362
rect 29586 21359 29598 21362
rect 29202 21313 29598 21359
rect 29202 21310 29214 21313
rect 29586 21310 29598 21313
rect 29650 21310 29662 21362
rect 28590 21298 28642 21310
rect 34078 21298 34130 21310
rect 35198 21362 35250 21374
rect 35198 21298 35250 21310
rect 35646 21362 35698 21374
rect 42242 21310 42254 21362
rect 42306 21310 42318 21362
rect 35646 21298 35698 21310
rect 1344 21194 44576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 44576 21194
rect 1344 21108 44576 21142
rect 13694 21026 13746 21038
rect 13694 20962 13746 20974
rect 19294 21026 19346 21038
rect 19294 20962 19346 20974
rect 21534 21026 21586 21038
rect 21534 20962 21586 20974
rect 26350 21026 26402 21038
rect 26350 20962 26402 20974
rect 31502 21026 31554 21038
rect 31502 20962 31554 20974
rect 31838 21026 31890 21038
rect 31838 20962 31890 20974
rect 35870 21026 35922 21038
rect 35870 20962 35922 20974
rect 4398 20914 4450 20926
rect 19182 20914 19234 20926
rect 35310 20914 35362 20926
rect 5954 20862 5966 20914
rect 6018 20862 6030 20914
rect 15362 20862 15374 20914
rect 15426 20862 15438 20914
rect 17490 20862 17502 20914
rect 17554 20862 17566 20914
rect 27906 20862 27918 20914
rect 27970 20862 27982 20914
rect 33954 20862 33966 20914
rect 34018 20862 34030 20914
rect 4398 20850 4450 20862
rect 19182 20850 19234 20862
rect 35310 20850 35362 20862
rect 35982 20914 36034 20926
rect 42366 20914 42418 20926
rect 37090 20862 37102 20914
rect 37154 20862 37166 20914
rect 41458 20862 41470 20914
rect 41522 20862 41534 20914
rect 35982 20850 36034 20862
rect 42366 20850 42418 20862
rect 13918 20802 13970 20814
rect 6066 20750 6078 20802
rect 6130 20750 6142 20802
rect 11554 20750 11566 20802
rect 11618 20750 11630 20802
rect 12002 20750 12014 20802
rect 12066 20750 12078 20802
rect 13918 20738 13970 20750
rect 14142 20802 14194 20814
rect 21870 20802 21922 20814
rect 26014 20802 26066 20814
rect 29822 20802 29874 20814
rect 18162 20750 18174 20802
rect 18226 20750 18238 20802
rect 18946 20750 18958 20802
rect 19010 20750 19022 20802
rect 20514 20750 20526 20802
rect 20578 20750 20590 20802
rect 25330 20750 25342 20802
rect 25394 20750 25406 20802
rect 27122 20750 27134 20802
rect 27186 20750 27198 20802
rect 27794 20750 27806 20802
rect 27858 20750 27870 20802
rect 14142 20738 14194 20750
rect 21870 20738 21922 20750
rect 26014 20738 26066 20750
rect 29822 20738 29874 20750
rect 30046 20802 30098 20814
rect 30046 20738 30098 20750
rect 30606 20802 30658 20814
rect 33070 20802 33122 20814
rect 32274 20750 32286 20802
rect 32338 20750 32350 20802
rect 30606 20738 30658 20750
rect 33070 20738 33122 20750
rect 33854 20802 33906 20814
rect 33854 20738 33906 20750
rect 34750 20802 34802 20814
rect 34750 20738 34802 20750
rect 34974 20802 35026 20814
rect 42926 20802 42978 20814
rect 38098 20750 38110 20802
rect 38162 20750 38174 20802
rect 38658 20750 38670 20802
rect 38722 20750 38734 20802
rect 43474 20750 43486 20802
rect 43538 20750 43550 20802
rect 34974 20738 35026 20750
rect 42926 20738 42978 20750
rect 5070 20690 5122 20702
rect 5070 20626 5122 20638
rect 5630 20690 5682 20702
rect 13470 20690 13522 20702
rect 9202 20638 9214 20690
rect 9266 20638 9278 20690
rect 5630 20626 5682 20638
rect 13470 20626 13522 20638
rect 14590 20690 14642 20702
rect 14590 20626 14642 20638
rect 19742 20690 19794 20702
rect 19742 20626 19794 20638
rect 20078 20690 20130 20702
rect 20078 20626 20130 20638
rect 20750 20690 20802 20702
rect 23214 20690 23266 20702
rect 29262 20690 29314 20702
rect 22082 20638 22094 20690
rect 22146 20638 22158 20690
rect 22642 20638 22654 20690
rect 22706 20638 22718 20690
rect 26898 20638 26910 20690
rect 26962 20638 26974 20690
rect 28130 20638 28142 20690
rect 28194 20638 28206 20690
rect 20750 20626 20802 20638
rect 23214 20626 23266 20638
rect 29262 20626 29314 20638
rect 29486 20690 29538 20702
rect 29486 20626 29538 20638
rect 30494 20690 30546 20702
rect 34190 20690 34242 20702
rect 32386 20638 32398 20690
rect 32450 20638 32462 20690
rect 30494 20626 30546 20638
rect 34190 20626 34242 20638
rect 34414 20690 34466 20702
rect 34414 20626 34466 20638
rect 35198 20690 35250 20702
rect 35198 20626 35250 20638
rect 37214 20690 37266 20702
rect 37214 20626 37266 20638
rect 37662 20690 37714 20702
rect 37662 20626 37714 20638
rect 4286 20578 4338 20590
rect 4286 20514 4338 20526
rect 4734 20578 4786 20590
rect 4734 20514 4786 20526
rect 8430 20578 8482 20590
rect 8430 20514 8482 20526
rect 25566 20578 25618 20590
rect 25566 20514 25618 20526
rect 29598 20578 29650 20590
rect 29598 20514 29650 20526
rect 30270 20578 30322 20590
rect 30270 20514 30322 20526
rect 33406 20578 33458 20590
rect 33406 20514 33458 20526
rect 33966 20578 34018 20590
rect 33966 20514 34018 20526
rect 35422 20578 35474 20590
rect 35422 20514 35474 20526
rect 36430 20578 36482 20590
rect 36430 20514 36482 20526
rect 37102 20578 37154 20590
rect 37102 20514 37154 20526
rect 37438 20578 37490 20590
rect 43262 20578 43314 20590
rect 41122 20526 41134 20578
rect 41186 20526 41198 20578
rect 37438 20514 37490 20526
rect 43262 20514 43314 20526
rect 44270 20578 44322 20590
rect 44270 20514 44322 20526
rect 1344 20410 44576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 44576 20410
rect 1344 20324 44576 20358
rect 11454 20242 11506 20254
rect 4834 20190 4846 20242
rect 4898 20190 4910 20242
rect 11454 20178 11506 20190
rect 14478 20242 14530 20254
rect 35534 20242 35586 20254
rect 26562 20190 26574 20242
rect 26626 20190 26638 20242
rect 39106 20190 39118 20242
rect 39170 20190 39182 20242
rect 14478 20178 14530 20190
rect 35534 20178 35586 20190
rect 5630 20130 5682 20142
rect 5630 20066 5682 20078
rect 11342 20130 11394 20142
rect 11342 20066 11394 20078
rect 12350 20130 12402 20142
rect 12350 20066 12402 20078
rect 12574 20130 12626 20142
rect 12574 20066 12626 20078
rect 12686 20130 12738 20142
rect 12686 20066 12738 20078
rect 12910 20130 12962 20142
rect 12910 20066 12962 20078
rect 14254 20130 14306 20142
rect 14254 20066 14306 20078
rect 17838 20130 17890 20142
rect 25902 20130 25954 20142
rect 32062 20130 32114 20142
rect 19170 20078 19182 20130
rect 19234 20078 19246 20130
rect 20626 20078 20638 20130
rect 20690 20078 20702 20130
rect 26786 20078 26798 20130
rect 26850 20078 26862 20130
rect 27906 20078 27918 20130
rect 27970 20078 27982 20130
rect 29250 20078 29262 20130
rect 29314 20078 29326 20130
rect 31714 20078 31726 20130
rect 31778 20078 31790 20130
rect 17838 20066 17890 20078
rect 25902 20066 25954 20078
rect 32062 20066 32114 20078
rect 32510 20130 32562 20142
rect 32510 20066 32562 20078
rect 33070 20130 33122 20142
rect 33070 20066 33122 20078
rect 34190 20130 34242 20142
rect 34190 20066 34242 20078
rect 40014 20130 40066 20142
rect 40014 20066 40066 20078
rect 40350 20130 40402 20142
rect 40350 20066 40402 20078
rect 40910 20130 40962 20142
rect 40910 20066 40962 20078
rect 43822 20130 43874 20142
rect 43822 20066 43874 20078
rect 12014 20018 12066 20030
rect 2034 19966 2046 20018
rect 2098 19966 2110 20018
rect 2594 19966 2606 20018
rect 2658 19966 2670 20018
rect 12014 19954 12066 19966
rect 12126 20018 12178 20030
rect 14590 20018 14642 20030
rect 13346 19966 13358 20018
rect 13410 19966 13422 20018
rect 12126 19954 12178 19966
rect 14590 19954 14642 19966
rect 14702 20018 14754 20030
rect 14702 19954 14754 19966
rect 14814 20018 14866 20030
rect 18286 20018 18338 20030
rect 25790 20018 25842 20030
rect 17602 19966 17614 20018
rect 17666 19966 17678 20018
rect 19394 19966 19406 20018
rect 19458 19966 19470 20018
rect 19954 19966 19966 20018
rect 20018 19966 20030 20018
rect 14814 19954 14866 19966
rect 18286 19954 18338 19966
rect 25790 19954 25842 19966
rect 26126 20018 26178 20030
rect 27582 20018 27634 20030
rect 33406 20018 33458 20030
rect 27010 19966 27022 20018
rect 27074 19966 27086 20018
rect 28578 19966 28590 20018
rect 28642 19966 28654 20018
rect 26126 19954 26178 19966
rect 27582 19954 27634 19966
rect 33406 19954 33458 19966
rect 33966 20018 34018 20030
rect 33966 19954 34018 19966
rect 34638 20018 34690 20030
rect 34638 19954 34690 19966
rect 35198 20018 35250 20030
rect 35198 19954 35250 19966
rect 35422 20018 35474 20030
rect 35422 19954 35474 19966
rect 35646 20018 35698 20030
rect 35646 19954 35698 19966
rect 35982 20018 36034 20030
rect 39678 20018 39730 20030
rect 44158 20018 44210 20030
rect 36530 19966 36542 20018
rect 36594 19966 36606 20018
rect 41794 19966 41806 20018
rect 41858 19966 41870 20018
rect 42802 19966 42814 20018
rect 42866 19966 42878 20018
rect 35982 19954 36034 19966
rect 39678 19954 39730 19966
rect 44158 19954 44210 19966
rect 15262 19906 15314 19918
rect 32398 19906 32450 19918
rect 13794 19854 13806 19906
rect 13858 19854 13870 19906
rect 22754 19854 22766 19906
rect 22818 19854 22830 19906
rect 31378 19854 31390 19906
rect 31442 19854 31454 19906
rect 15262 19842 15314 19854
rect 32398 19842 32450 19854
rect 34414 19906 34466 19918
rect 34414 19842 34466 19854
rect 34974 19906 35026 19918
rect 41682 19854 41694 19906
rect 41746 19854 41758 19906
rect 42578 19854 42590 19906
rect 42642 19854 42654 19906
rect 34974 19842 35026 19854
rect 15374 19794 15426 19806
rect 15374 19730 15426 19742
rect 18622 19794 18674 19806
rect 42690 19742 42702 19794
rect 42754 19742 42766 19794
rect 18622 19730 18674 19742
rect 1344 19626 44576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 44576 19626
rect 1344 19540 44576 19574
rect 27134 19458 27186 19470
rect 27134 19394 27186 19406
rect 28254 19458 28306 19470
rect 28254 19394 28306 19406
rect 32846 19458 32898 19470
rect 32846 19394 32898 19406
rect 36990 19458 37042 19470
rect 36990 19394 37042 19406
rect 12238 19346 12290 19358
rect 28366 19346 28418 19358
rect 37102 19346 37154 19358
rect 6514 19294 6526 19346
rect 6578 19294 6590 19346
rect 14130 19294 14142 19346
rect 14194 19294 14206 19346
rect 18162 19294 18174 19346
rect 18226 19294 18238 19346
rect 20290 19294 20302 19346
rect 20354 19294 20366 19346
rect 22082 19294 22094 19346
rect 22146 19294 22158 19346
rect 29922 19294 29934 19346
rect 29986 19294 29998 19346
rect 32050 19294 32062 19346
rect 32114 19294 32126 19346
rect 33954 19294 33966 19346
rect 34018 19294 34030 19346
rect 36082 19294 36094 19346
rect 36146 19294 36158 19346
rect 44034 19294 44046 19346
rect 44098 19294 44110 19346
rect 12238 19282 12290 19294
rect 28366 19282 28418 19294
rect 37102 19282 37154 19294
rect 3278 19234 3330 19246
rect 4958 19234 5010 19246
rect 4610 19182 4622 19234
rect 4674 19182 4686 19234
rect 3278 19170 3330 19182
rect 4958 19170 5010 19182
rect 5070 19234 5122 19246
rect 5070 19170 5122 19182
rect 5966 19234 6018 19246
rect 27246 19234 27298 19246
rect 6850 19182 6862 19234
rect 6914 19182 6926 19234
rect 11890 19182 11902 19234
rect 11954 19182 11966 19234
rect 17042 19182 17054 19234
rect 17106 19182 17118 19234
rect 17378 19182 17390 19234
rect 17442 19182 17454 19234
rect 22306 19182 22318 19234
rect 22370 19182 22382 19234
rect 29138 19182 29150 19234
rect 29202 19182 29214 19234
rect 32834 19182 32846 19234
rect 32898 19182 32910 19234
rect 33282 19182 33294 19234
rect 33346 19182 33358 19234
rect 40674 19182 40686 19234
rect 40738 19182 40750 19234
rect 41122 19182 41134 19234
rect 41186 19182 41198 19234
rect 5966 19170 6018 19182
rect 27246 19170 27298 19182
rect 3166 19122 3218 19134
rect 3166 19058 3218 19070
rect 7422 19122 7474 19134
rect 7422 19058 7474 19070
rect 12126 19122 12178 19134
rect 27918 19122 27970 19134
rect 16258 19070 16270 19122
rect 16322 19070 16334 19122
rect 21970 19070 21982 19122
rect 22034 19070 22046 19122
rect 12126 19058 12178 19070
rect 27918 19058 27970 19070
rect 32510 19122 32562 19134
rect 32510 19058 32562 19070
rect 40238 19122 40290 19134
rect 40238 19058 40290 19070
rect 5630 19010 5682 19022
rect 5630 18946 5682 18958
rect 12350 19010 12402 19022
rect 12350 18946 12402 18958
rect 12462 19010 12514 19022
rect 12462 18946 12514 18958
rect 20750 19010 20802 19022
rect 20750 18946 20802 18958
rect 27134 19010 27186 19022
rect 28478 19010 28530 19022
rect 27570 18958 27582 19010
rect 27634 18958 27646 19010
rect 27134 18946 27186 18958
rect 28478 18946 28530 18958
rect 40350 19010 40402 19022
rect 43474 18958 43486 19010
rect 43538 18958 43550 19010
rect 40350 18946 40402 18958
rect 1344 18842 44576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 44576 18842
rect 1344 18756 44576 18790
rect 1598 18674 1650 18686
rect 15710 18674 15762 18686
rect 2370 18622 2382 18674
rect 2434 18622 2446 18674
rect 1598 18610 1650 18622
rect 15710 18610 15762 18622
rect 15822 18674 15874 18686
rect 15822 18610 15874 18622
rect 43374 18674 43426 18686
rect 43374 18610 43426 18622
rect 7646 18562 7698 18574
rect 7646 18498 7698 18510
rect 8318 18562 8370 18574
rect 8318 18498 8370 18510
rect 10446 18562 10498 18574
rect 10446 18498 10498 18510
rect 10670 18562 10722 18574
rect 10670 18498 10722 18510
rect 15038 18562 15090 18574
rect 15038 18498 15090 18510
rect 15598 18562 15650 18574
rect 15598 18498 15650 18510
rect 17502 18562 17554 18574
rect 17502 18498 17554 18510
rect 17614 18562 17666 18574
rect 24110 18562 24162 18574
rect 18274 18510 18286 18562
rect 18338 18510 18350 18562
rect 17614 18498 17666 18510
rect 24110 18498 24162 18510
rect 25230 18562 25282 18574
rect 29486 18562 29538 18574
rect 32398 18562 32450 18574
rect 35870 18562 35922 18574
rect 28354 18510 28366 18562
rect 28418 18510 28430 18562
rect 29922 18510 29934 18562
rect 29986 18510 29998 18562
rect 33394 18510 33406 18562
rect 33458 18510 33470 18562
rect 25230 18498 25282 18510
rect 29486 18498 29538 18510
rect 32398 18498 32450 18510
rect 35870 18498 35922 18510
rect 36654 18562 36706 18574
rect 36654 18498 36706 18510
rect 41246 18562 41298 18574
rect 41246 18498 41298 18510
rect 7198 18450 7250 18462
rect 10894 18450 10946 18462
rect 4722 18398 4734 18450
rect 4786 18398 4798 18450
rect 5170 18398 5182 18450
rect 5234 18398 5246 18450
rect 6626 18398 6638 18450
rect 6690 18398 6702 18450
rect 7858 18398 7870 18450
rect 7922 18398 7934 18450
rect 8530 18398 8542 18450
rect 8594 18398 8606 18450
rect 7198 18386 7250 18398
rect 10894 18386 10946 18398
rect 11118 18450 11170 18462
rect 11118 18386 11170 18398
rect 11678 18450 11730 18462
rect 11678 18386 11730 18398
rect 12574 18450 12626 18462
rect 12574 18386 12626 18398
rect 13694 18450 13746 18462
rect 14814 18450 14866 18462
rect 14466 18398 14478 18450
rect 14530 18398 14542 18450
rect 13694 18386 13746 18398
rect 14814 18386 14866 18398
rect 16270 18450 16322 18462
rect 16270 18386 16322 18398
rect 17278 18450 17330 18462
rect 17278 18386 17330 18398
rect 18622 18450 18674 18462
rect 21198 18450 21250 18462
rect 20626 18398 20638 18450
rect 20690 18398 20702 18450
rect 18622 18386 18674 18398
rect 21198 18386 21250 18398
rect 24446 18450 24498 18462
rect 26910 18450 26962 18462
rect 29262 18450 29314 18462
rect 31054 18450 31106 18462
rect 25442 18398 25454 18450
rect 25506 18398 25518 18450
rect 26450 18398 26462 18450
rect 26514 18398 26526 18450
rect 28242 18398 28254 18450
rect 28306 18398 28318 18450
rect 30146 18398 30158 18450
rect 30210 18398 30222 18450
rect 24446 18386 24498 18398
rect 26910 18386 26962 18398
rect 29262 18386 29314 18398
rect 31054 18386 31106 18398
rect 31166 18450 31218 18462
rect 31166 18386 31218 18398
rect 31838 18450 31890 18462
rect 31838 18386 31890 18398
rect 32174 18450 32226 18462
rect 32174 18386 32226 18398
rect 33070 18450 33122 18462
rect 33070 18386 33122 18398
rect 34078 18450 34130 18462
rect 34078 18386 34130 18398
rect 34302 18450 34354 18462
rect 34302 18386 34354 18398
rect 34638 18450 34690 18462
rect 34638 18386 34690 18398
rect 34862 18450 34914 18462
rect 34862 18386 34914 18398
rect 35310 18450 35362 18462
rect 35310 18386 35362 18398
rect 35534 18450 35586 18462
rect 35534 18386 35586 18398
rect 36206 18450 36258 18462
rect 36206 18386 36258 18398
rect 36542 18450 36594 18462
rect 36542 18386 36594 18398
rect 40014 18450 40066 18462
rect 42702 18450 42754 18462
rect 42018 18398 42030 18450
rect 42082 18398 42094 18450
rect 40014 18386 40066 18398
rect 42702 18386 42754 18398
rect 43038 18450 43090 18462
rect 43038 18386 43090 18398
rect 10558 18338 10610 18350
rect 6402 18286 6414 18338
rect 6466 18286 6478 18338
rect 10558 18274 10610 18286
rect 11454 18338 11506 18350
rect 11454 18274 11506 18286
rect 11902 18338 11954 18350
rect 11902 18274 11954 18286
rect 14926 18338 14978 18350
rect 14926 18274 14978 18286
rect 21758 18338 21810 18350
rect 27918 18338 27970 18350
rect 30718 18338 30770 18350
rect 34526 18338 34578 18350
rect 26338 18286 26350 18338
rect 26402 18286 26414 18338
rect 28914 18286 28926 18338
rect 28978 18286 28990 18338
rect 29586 18286 29598 18338
rect 29650 18286 29662 18338
rect 32498 18286 32510 18338
rect 32562 18286 32574 18338
rect 21758 18274 21810 18286
rect 27918 18274 27970 18286
rect 30718 18274 30770 18286
rect 34526 18274 34578 18286
rect 35086 18338 35138 18350
rect 35086 18274 35138 18286
rect 37102 18338 37154 18350
rect 37102 18274 37154 18286
rect 40126 18338 40178 18350
rect 42242 18286 42254 18338
rect 42306 18286 42318 18338
rect 40126 18274 40178 18286
rect 12126 18226 12178 18238
rect 12126 18162 12178 18174
rect 13806 18226 13858 18238
rect 13806 18162 13858 18174
rect 20974 18226 21026 18238
rect 20974 18162 21026 18174
rect 26126 18226 26178 18238
rect 26126 18162 26178 18174
rect 41134 18226 41186 18238
rect 41134 18162 41186 18174
rect 1344 18058 44576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 44576 18058
rect 1344 17972 44576 18006
rect 9774 17890 9826 17902
rect 9774 17826 9826 17838
rect 11454 17890 11506 17902
rect 37102 17890 37154 17902
rect 27682 17838 27694 17890
rect 27746 17838 27758 17890
rect 11454 17826 11506 17838
rect 37102 17826 37154 17838
rect 9662 17778 9714 17790
rect 5954 17726 5966 17778
rect 6018 17726 6030 17778
rect 9662 17714 9714 17726
rect 11678 17778 11730 17790
rect 11678 17714 11730 17726
rect 12014 17778 12066 17790
rect 22318 17778 22370 17790
rect 13458 17726 13470 17778
rect 13522 17726 13534 17778
rect 15586 17726 15598 17778
rect 15650 17726 15662 17778
rect 12014 17714 12066 17726
rect 22318 17714 22370 17726
rect 23438 17778 23490 17790
rect 28142 17778 28194 17790
rect 37550 17778 37602 17790
rect 24658 17726 24670 17778
rect 24722 17726 24734 17778
rect 26786 17726 26798 17778
rect 26850 17726 26862 17778
rect 36418 17726 36430 17778
rect 36482 17726 36494 17778
rect 42130 17726 42142 17778
rect 42194 17726 42206 17778
rect 23438 17714 23490 17726
rect 28142 17714 28194 17726
rect 37550 17714 37602 17726
rect 16606 17666 16658 17678
rect 8866 17614 8878 17666
rect 8930 17614 8942 17666
rect 9314 17614 9326 17666
rect 9378 17614 9390 17666
rect 10322 17614 10334 17666
rect 10386 17614 10398 17666
rect 16258 17614 16270 17666
rect 16322 17614 16334 17666
rect 16606 17602 16658 17614
rect 16942 17666 16994 17678
rect 16942 17602 16994 17614
rect 19182 17666 19234 17678
rect 19182 17602 19234 17614
rect 19854 17666 19906 17678
rect 19854 17602 19906 17614
rect 20302 17666 20354 17678
rect 20302 17602 20354 17614
rect 20526 17666 20578 17678
rect 20526 17602 20578 17614
rect 20862 17666 20914 17678
rect 20862 17602 20914 17614
rect 21534 17666 21586 17678
rect 21534 17602 21586 17614
rect 21870 17666 21922 17678
rect 27134 17666 27186 17678
rect 23986 17614 23998 17666
rect 24050 17614 24062 17666
rect 21870 17602 21922 17614
rect 27134 17602 27186 17614
rect 27358 17666 27410 17678
rect 38894 17666 38946 17678
rect 42590 17666 42642 17678
rect 32274 17614 32286 17666
rect 32338 17614 32350 17666
rect 33058 17614 33070 17666
rect 33122 17614 33134 17666
rect 33506 17614 33518 17666
rect 33570 17614 33582 17666
rect 39330 17614 39342 17666
rect 39394 17614 39406 17666
rect 27358 17602 27410 17614
rect 38894 17602 38946 17614
rect 42590 17602 42642 17614
rect 18846 17554 18898 17566
rect 6514 17502 6526 17554
rect 6578 17502 6590 17554
rect 18846 17490 18898 17502
rect 19518 17554 19570 17566
rect 19518 17490 19570 17502
rect 21310 17554 21362 17566
rect 21310 17490 21362 17502
rect 22206 17554 22258 17566
rect 22206 17490 22258 17502
rect 22430 17554 22482 17566
rect 22430 17490 22482 17502
rect 22990 17554 23042 17566
rect 22990 17490 23042 17502
rect 28030 17554 28082 17566
rect 36990 17554 37042 17566
rect 34290 17502 34302 17554
rect 34354 17502 34366 17554
rect 28030 17490 28082 17502
rect 36990 17490 37042 17502
rect 10110 17442 10162 17454
rect 10110 17378 10162 17390
rect 11902 17442 11954 17454
rect 11902 17378 11954 17390
rect 12126 17442 12178 17454
rect 12126 17378 12178 17390
rect 16830 17442 16882 17454
rect 16830 17378 16882 17390
rect 17502 17442 17554 17454
rect 17502 17378 17554 17390
rect 17838 17442 17890 17454
rect 17838 17378 17890 17390
rect 20526 17442 20578 17454
rect 20526 17378 20578 17390
rect 21422 17442 21474 17454
rect 21422 17378 21474 17390
rect 22878 17442 22930 17454
rect 22878 17378 22930 17390
rect 28254 17442 28306 17454
rect 28254 17378 28306 17390
rect 29374 17442 29426 17454
rect 32846 17442 32898 17454
rect 32498 17390 32510 17442
rect 32562 17390 32574 17442
rect 29374 17378 29426 17390
rect 32846 17378 32898 17390
rect 37438 17442 37490 17454
rect 42926 17442 42978 17454
rect 41794 17390 41806 17442
rect 41858 17390 41870 17442
rect 37438 17378 37490 17390
rect 42926 17378 42978 17390
rect 1344 17274 44576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 44576 17274
rect 1344 17188 44576 17222
rect 18286 17106 18338 17118
rect 6066 17054 6078 17106
rect 6130 17054 6142 17106
rect 18286 17042 18338 17054
rect 18510 17106 18562 17118
rect 18510 17042 18562 17054
rect 23886 17106 23938 17118
rect 23886 17042 23938 17054
rect 25342 17106 25394 17118
rect 25342 17042 25394 17054
rect 27806 17106 27858 17118
rect 27806 17042 27858 17054
rect 30830 17106 30882 17118
rect 40350 17106 40402 17118
rect 39778 17054 39790 17106
rect 39842 17054 39854 17106
rect 30830 17042 30882 17054
rect 40350 17042 40402 17054
rect 41918 17106 41970 17118
rect 43810 17054 43822 17106
rect 43874 17054 43886 17106
rect 41918 17042 41970 17054
rect 13134 16994 13186 17006
rect 13134 16930 13186 16942
rect 23438 16994 23490 17006
rect 28254 16994 28306 17006
rect 26450 16942 26462 16994
rect 26514 16942 26526 16994
rect 34178 16942 34190 16994
rect 34242 16942 34254 16994
rect 23438 16930 23490 16942
rect 28254 16930 28306 16942
rect 5294 16882 5346 16894
rect 8990 16882 9042 16894
rect 19070 16882 19122 16894
rect 23998 16882 24050 16894
rect 8306 16830 8318 16882
rect 8370 16830 8382 16882
rect 9986 16830 9998 16882
rect 10050 16830 10062 16882
rect 10658 16830 10670 16882
rect 10722 16830 10734 16882
rect 13346 16830 13358 16882
rect 13410 16830 13422 16882
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 19394 16830 19406 16882
rect 19458 16830 19470 16882
rect 22866 16830 22878 16882
rect 22930 16830 22942 16882
rect 5294 16818 5346 16830
rect 8990 16818 9042 16830
rect 19070 16818 19122 16830
rect 23998 16818 24050 16830
rect 24782 16882 24834 16894
rect 24782 16818 24834 16830
rect 25678 16882 25730 16894
rect 27470 16882 27522 16894
rect 26338 16830 26350 16882
rect 26402 16830 26414 16882
rect 25678 16818 25730 16830
rect 27470 16818 27522 16830
rect 28478 16882 28530 16894
rect 28478 16818 28530 16830
rect 29934 16882 29986 16894
rect 43598 16882 43650 16894
rect 33394 16830 33406 16882
rect 33458 16830 33470 16882
rect 36754 16830 36766 16882
rect 36818 16830 36830 16882
rect 37314 16830 37326 16882
rect 37378 16830 37390 16882
rect 42130 16830 42142 16882
rect 42194 16830 42206 16882
rect 29934 16818 29986 16830
rect 43598 16818 43650 16830
rect 44158 16882 44210 16894
rect 44158 16818 44210 16830
rect 12786 16718 12798 16770
rect 12850 16718 12862 16770
rect 14690 16718 14702 16770
rect 14754 16718 14766 16770
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 20178 16718 20190 16770
rect 20242 16718 20254 16770
rect 22306 16718 22318 16770
rect 22370 16718 22382 16770
rect 23090 16718 23102 16770
rect 23154 16718 23166 16770
rect 27794 16718 27806 16770
rect 27858 16718 27870 16770
rect 29474 16718 29486 16770
rect 29538 16718 29550 16770
rect 36306 16718 36318 16770
rect 36370 16718 36382 16770
rect 23886 16658 23938 16670
rect 23886 16594 23938 16606
rect 28814 16658 28866 16670
rect 28814 16594 28866 16606
rect 1344 16490 44576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 44576 16490
rect 1344 16404 44576 16438
rect 7198 16322 7250 16334
rect 7198 16258 7250 16270
rect 9886 16322 9938 16334
rect 9886 16258 9938 16270
rect 12798 16322 12850 16334
rect 12798 16258 12850 16270
rect 15934 16322 15986 16334
rect 33966 16322 34018 16334
rect 26898 16270 26910 16322
rect 26962 16270 26974 16322
rect 29138 16270 29150 16322
rect 29202 16270 29214 16322
rect 15934 16258 15986 16270
rect 33966 16258 34018 16270
rect 34302 16322 34354 16334
rect 34302 16258 34354 16270
rect 7086 16210 7138 16222
rect 7086 16146 7138 16158
rect 9102 16210 9154 16222
rect 9102 16146 9154 16158
rect 10446 16210 10498 16222
rect 10446 16146 10498 16158
rect 11230 16210 11282 16222
rect 11230 16146 11282 16158
rect 12462 16210 12514 16222
rect 12462 16146 12514 16158
rect 17278 16210 17330 16222
rect 17278 16146 17330 16158
rect 18846 16210 18898 16222
rect 18846 16146 18898 16158
rect 19966 16210 20018 16222
rect 19966 16146 20018 16158
rect 21758 16210 21810 16222
rect 29710 16210 29762 16222
rect 23426 16158 23438 16210
rect 23490 16158 23502 16210
rect 21758 16146 21810 16158
rect 29710 16146 29762 16158
rect 33070 16210 33122 16222
rect 43922 16158 43934 16210
rect 43986 16158 43998 16210
rect 33070 16146 33122 16158
rect 10110 16098 10162 16110
rect 10110 16034 10162 16046
rect 10334 16098 10386 16110
rect 10334 16034 10386 16046
rect 15150 16098 15202 16110
rect 19070 16098 19122 16110
rect 20078 16098 20130 16110
rect 16594 16046 16606 16098
rect 16658 16046 16670 16098
rect 19730 16046 19742 16098
rect 19794 16046 19806 16098
rect 15150 16034 15202 16046
rect 19070 16034 19122 16046
rect 20078 16034 20130 16046
rect 20750 16098 20802 16110
rect 20750 16034 20802 16046
rect 21310 16098 21362 16110
rect 21310 16034 21362 16046
rect 21646 16098 21698 16110
rect 21646 16034 21698 16046
rect 21870 16098 21922 16110
rect 23886 16098 23938 16110
rect 23090 16046 23102 16098
rect 23154 16046 23166 16098
rect 21870 16034 21922 16046
rect 23886 16034 23938 16046
rect 25342 16098 25394 16110
rect 28478 16098 28530 16110
rect 25778 16046 25790 16098
rect 25842 16046 25854 16098
rect 27906 16046 27918 16098
rect 27970 16046 27982 16098
rect 25342 16034 25394 16046
rect 28478 16034 28530 16046
rect 29486 16098 29538 16110
rect 29486 16034 29538 16046
rect 31950 16098 32002 16110
rect 40014 16098 40066 16110
rect 32498 16046 32510 16098
rect 32562 16046 32574 16098
rect 34290 16046 34302 16098
rect 34354 16046 34366 16098
rect 39330 16046 39342 16098
rect 39394 16046 39406 16098
rect 31950 16034 32002 16046
rect 40014 16034 40066 16046
rect 40686 16098 40738 16110
rect 41122 16046 41134 16098
rect 41186 16046 41198 16098
rect 40686 16034 40738 16046
rect 9550 15986 9602 15998
rect 14142 15986 14194 15998
rect 11778 15934 11790 15986
rect 11842 15934 11854 15986
rect 12226 15934 12238 15986
rect 12290 15934 12302 15986
rect 9550 15922 9602 15934
rect 14142 15922 14194 15934
rect 14478 15986 14530 15998
rect 14478 15922 14530 15934
rect 14814 15986 14866 15998
rect 24894 15986 24946 15998
rect 40238 15986 40290 15998
rect 16706 15934 16718 15986
rect 16770 15934 16782 15986
rect 22194 15934 22206 15986
rect 22258 15934 22270 15986
rect 30034 15934 30046 15986
rect 30098 15934 30110 15986
rect 43362 15934 43374 15986
rect 43426 15934 43438 15986
rect 14814 15922 14866 15934
rect 24894 15922 24946 15934
rect 40238 15922 40290 15934
rect 9438 15874 9490 15886
rect 9438 15810 9490 15822
rect 10558 15874 10610 15886
rect 10558 15810 10610 15822
rect 11118 15874 11170 15886
rect 13806 15874 13858 15886
rect 13458 15822 13470 15874
rect 13522 15822 13534 15874
rect 11118 15810 11170 15822
rect 13806 15810 13858 15822
rect 15598 15874 15650 15886
rect 15598 15810 15650 15822
rect 17726 15874 17778 15886
rect 17726 15810 17778 15822
rect 19406 15874 19458 15886
rect 19406 15810 19458 15822
rect 20526 15874 20578 15886
rect 20526 15810 20578 15822
rect 20638 15874 20690 15886
rect 20638 15810 20690 15822
rect 22542 15874 22594 15886
rect 22542 15810 22594 15822
rect 24446 15874 24498 15886
rect 24446 15810 24498 15822
rect 28366 15874 28418 15886
rect 28366 15810 28418 15822
rect 30382 15874 30434 15886
rect 30382 15810 30434 15822
rect 30718 15874 30770 15886
rect 31614 15874 31666 15886
rect 31042 15822 31054 15874
rect 31106 15822 31118 15874
rect 30718 15810 30770 15822
rect 31614 15810 31666 15822
rect 32286 15874 32338 15886
rect 32286 15810 32338 15822
rect 38782 15874 38834 15886
rect 38782 15810 38834 15822
rect 1344 15706 44576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 44576 15706
rect 1344 15620 44576 15654
rect 8766 15538 8818 15550
rect 8766 15474 8818 15486
rect 13134 15538 13186 15550
rect 13134 15474 13186 15486
rect 14142 15538 14194 15550
rect 14142 15474 14194 15486
rect 14590 15538 14642 15550
rect 14590 15474 14642 15486
rect 15150 15538 15202 15550
rect 15150 15474 15202 15486
rect 19070 15538 19122 15550
rect 30046 15538 30098 15550
rect 27010 15486 27022 15538
rect 27074 15486 27086 15538
rect 19070 15474 19122 15486
rect 30046 15474 30098 15486
rect 30606 15538 30658 15550
rect 30606 15474 30658 15486
rect 32398 15538 32450 15550
rect 32398 15474 32450 15486
rect 40910 15538 40962 15550
rect 40910 15474 40962 15486
rect 8990 15426 9042 15438
rect 8990 15362 9042 15374
rect 13358 15426 13410 15438
rect 13358 15362 13410 15374
rect 15486 15426 15538 15438
rect 15486 15362 15538 15374
rect 19518 15426 19570 15438
rect 25230 15426 25282 15438
rect 24322 15374 24334 15426
rect 24386 15374 24398 15426
rect 19518 15362 19570 15374
rect 25230 15362 25282 15374
rect 25454 15426 25506 15438
rect 25454 15362 25506 15374
rect 25678 15426 25730 15438
rect 30382 15426 30434 15438
rect 39902 15426 39954 15438
rect 26338 15374 26350 15426
rect 26402 15374 26414 15426
rect 26786 15374 26798 15426
rect 26850 15374 26862 15426
rect 27570 15374 27582 15426
rect 27634 15374 27646 15426
rect 28130 15374 28142 15426
rect 28194 15374 28206 15426
rect 28578 15374 28590 15426
rect 28642 15374 28654 15426
rect 31378 15374 31390 15426
rect 31442 15374 31454 15426
rect 25678 15362 25730 15374
rect 30382 15362 30434 15374
rect 39902 15362 39954 15374
rect 8878 15314 8930 15326
rect 12686 15314 12738 15326
rect 8418 15262 8430 15314
rect 8482 15262 8494 15314
rect 9650 15262 9662 15314
rect 9714 15262 9726 15314
rect 8878 15250 8930 15262
rect 12686 15250 12738 15262
rect 19294 15314 19346 15326
rect 19294 15250 19346 15262
rect 19630 15314 19682 15326
rect 19954 15262 19966 15314
rect 20018 15262 20030 15314
rect 20738 15262 20750 15314
rect 20802 15262 20814 15314
rect 24210 15262 24222 15314
rect 24274 15262 24286 15314
rect 26114 15262 26126 15314
rect 26178 15262 26190 15314
rect 27682 15262 27694 15314
rect 27746 15262 27758 15314
rect 28466 15262 28478 15314
rect 28530 15262 28542 15314
rect 31266 15262 31278 15314
rect 31330 15262 31342 15314
rect 39666 15262 39678 15314
rect 39730 15262 39742 15314
rect 41122 15262 41134 15314
rect 41186 15262 41198 15314
rect 42466 15262 42478 15314
rect 42530 15262 42542 15314
rect 43474 15262 43486 15314
rect 43538 15262 43550 15314
rect 19630 15250 19682 15262
rect 13246 15202 13298 15214
rect 23662 15202 23714 15214
rect 10322 15150 10334 15202
rect 10386 15150 10398 15202
rect 12450 15150 12462 15202
rect 12514 15150 12526 15202
rect 22866 15150 22878 15202
rect 22930 15150 22942 15202
rect 13246 15138 13298 15150
rect 23662 15138 23714 15150
rect 29486 15202 29538 15214
rect 29486 15138 29538 15150
rect 30494 15202 30546 15214
rect 30494 15138 30546 15150
rect 39230 15202 39282 15214
rect 43038 15202 43090 15214
rect 42018 15150 42030 15202
rect 42082 15150 42094 15202
rect 39230 15138 39282 15150
rect 43038 15138 43090 15150
rect 23326 15090 23378 15102
rect 23326 15026 23378 15038
rect 25790 15090 25842 15102
rect 25790 15026 25842 15038
rect 28590 15090 28642 15102
rect 28590 15026 28642 15038
rect 32062 15090 32114 15102
rect 41906 15038 41918 15090
rect 41970 15038 41982 15090
rect 32062 15026 32114 15038
rect 1344 14922 44576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 44576 14922
rect 1344 14836 44576 14870
rect 13582 14754 13634 14766
rect 13582 14690 13634 14702
rect 21310 14754 21362 14766
rect 26562 14702 26574 14754
rect 26626 14702 26638 14754
rect 21310 14690 21362 14702
rect 14254 14642 14306 14654
rect 9762 14590 9774 14642
rect 9826 14590 9838 14642
rect 11890 14590 11902 14642
rect 11954 14590 11966 14642
rect 14254 14578 14306 14590
rect 21422 14642 21474 14654
rect 21422 14578 21474 14590
rect 21870 14642 21922 14654
rect 25442 14590 25454 14642
rect 25506 14590 25518 14642
rect 28242 14590 28254 14642
rect 28306 14590 28318 14642
rect 31938 14590 31950 14642
rect 32002 14590 32014 14642
rect 34066 14590 34078 14642
rect 34130 14590 34142 14642
rect 34738 14590 34750 14642
rect 34802 14590 34814 14642
rect 21870 14578 21922 14590
rect 12238 14530 12290 14542
rect 9090 14478 9102 14530
rect 9154 14478 9166 14530
rect 12238 14466 12290 14478
rect 12574 14530 12626 14542
rect 12574 14466 12626 14478
rect 13694 14530 13746 14542
rect 13694 14466 13746 14478
rect 15150 14530 15202 14542
rect 15150 14466 15202 14478
rect 18734 14530 18786 14542
rect 19518 14530 19570 14542
rect 19170 14478 19182 14530
rect 19234 14478 19246 14530
rect 18734 14466 18786 14478
rect 19518 14466 19570 14478
rect 20078 14530 20130 14542
rect 21646 14530 21698 14542
rect 26014 14530 26066 14542
rect 41246 14530 41298 14542
rect 20514 14478 20526 14530
rect 20578 14478 20590 14530
rect 22642 14478 22654 14530
rect 22706 14478 22718 14530
rect 25778 14478 25790 14530
rect 25842 14478 25854 14530
rect 27794 14478 27806 14530
rect 27858 14478 27870 14530
rect 28130 14478 28142 14530
rect 28194 14478 28206 14530
rect 29138 14478 29150 14530
rect 29202 14478 29214 14530
rect 30594 14478 30606 14530
rect 30658 14478 30670 14530
rect 30930 14478 30942 14530
rect 30994 14478 31006 14530
rect 31154 14478 31166 14530
rect 31218 14478 31230 14530
rect 40786 14478 40798 14530
rect 40850 14478 40862 14530
rect 20078 14466 20130 14478
rect 21646 14466 21698 14478
rect 26014 14466 26066 14478
rect 16718 14418 16770 14430
rect 26126 14418 26178 14430
rect 15474 14366 15486 14418
rect 15538 14366 15550 14418
rect 15698 14366 15710 14418
rect 15762 14366 15774 14418
rect 20738 14366 20750 14418
rect 20802 14366 20814 14418
rect 23314 14366 23326 14418
rect 23378 14366 23390 14418
rect 29250 14366 29262 14418
rect 29314 14366 29326 14418
rect 30594 14366 30606 14418
rect 30658 14415 30670 14418
rect 30945 14415 30991 14478
rect 41246 14466 41298 14478
rect 41806 14530 41858 14542
rect 42018 14478 42030 14530
rect 42082 14478 42094 14530
rect 41806 14466 41858 14478
rect 30658 14369 30991 14415
rect 34414 14418 34466 14430
rect 30658 14366 30670 14369
rect 16718 14354 16770 14366
rect 26126 14354 26178 14366
rect 34414 14354 34466 14366
rect 34638 14418 34690 14430
rect 34638 14354 34690 14366
rect 41582 14418 41634 14430
rect 41582 14354 41634 14366
rect 12350 14306 12402 14318
rect 12350 14242 12402 14254
rect 13022 14306 13074 14318
rect 13022 14242 13074 14254
rect 13582 14306 13634 14318
rect 13582 14242 13634 14254
rect 14814 14306 14866 14318
rect 14814 14242 14866 14254
rect 16382 14306 16434 14318
rect 16382 14242 16434 14254
rect 17166 14306 17218 14318
rect 17166 14242 17218 14254
rect 18174 14306 18226 14318
rect 18174 14242 18226 14254
rect 18622 14306 18674 14318
rect 18622 14242 18674 14254
rect 18846 14306 18898 14318
rect 18846 14242 18898 14254
rect 18958 14306 19010 14318
rect 18958 14242 19010 14254
rect 21982 14306 22034 14318
rect 21982 14242 22034 14254
rect 22206 14306 22258 14318
rect 35758 14306 35810 14318
rect 28018 14254 28030 14306
rect 28082 14254 28094 14306
rect 30258 14254 30270 14306
rect 30322 14254 30334 14306
rect 30482 14254 30494 14306
rect 30546 14254 30558 14306
rect 22206 14242 22258 14254
rect 35758 14242 35810 14254
rect 1344 14138 44576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 44576 14138
rect 1344 14052 44576 14086
rect 17502 13970 17554 13982
rect 17502 13906 17554 13918
rect 18734 13970 18786 13982
rect 18734 13906 18786 13918
rect 19406 13970 19458 13982
rect 19406 13906 19458 13918
rect 23102 13970 23154 13982
rect 27134 13970 27186 13982
rect 25330 13918 25342 13970
rect 25394 13918 25406 13970
rect 26226 13918 26238 13970
rect 26290 13918 26302 13970
rect 23102 13906 23154 13918
rect 27134 13906 27186 13918
rect 27358 13970 27410 13982
rect 27358 13906 27410 13918
rect 28702 13970 28754 13982
rect 28702 13906 28754 13918
rect 30830 13970 30882 13982
rect 40014 13970 40066 13982
rect 39106 13918 39118 13970
rect 39170 13918 39182 13970
rect 30830 13906 30882 13918
rect 40014 13906 40066 13918
rect 42702 13970 42754 13982
rect 42702 13906 42754 13918
rect 18958 13858 19010 13870
rect 16594 13806 16606 13858
rect 16658 13806 16670 13858
rect 18958 13794 19010 13806
rect 19070 13858 19122 13870
rect 19070 13794 19122 13806
rect 20302 13858 20354 13870
rect 27022 13858 27074 13870
rect 26562 13806 26574 13858
rect 26626 13806 26638 13858
rect 20302 13794 20354 13806
rect 27022 13794 27074 13806
rect 29150 13858 29202 13870
rect 31838 13858 31890 13870
rect 30482 13806 30494 13858
rect 30546 13806 30558 13858
rect 31490 13806 31502 13858
rect 31554 13806 31566 13858
rect 29150 13794 29202 13806
rect 31838 13794 31890 13806
rect 32062 13858 32114 13870
rect 32062 13794 32114 13806
rect 33070 13858 33122 13870
rect 33070 13794 33122 13806
rect 33406 13858 33458 13870
rect 33406 13794 33458 13806
rect 34190 13858 34242 13870
rect 34190 13794 34242 13806
rect 34750 13858 34802 13870
rect 34750 13794 34802 13806
rect 35086 13858 35138 13870
rect 35086 13794 35138 13806
rect 15934 13746 15986 13758
rect 28366 13746 28418 13758
rect 34526 13746 34578 13758
rect 35982 13746 36034 13758
rect 40350 13746 40402 13758
rect 10882 13694 10894 13746
rect 10946 13694 10958 13746
rect 16482 13694 16494 13746
rect 16546 13694 16558 13746
rect 20402 13694 20414 13746
rect 20466 13694 20478 13746
rect 20850 13694 20862 13746
rect 20914 13694 20926 13746
rect 22866 13694 22878 13746
rect 22930 13694 22942 13746
rect 25554 13694 25566 13746
rect 25618 13694 25630 13746
rect 26450 13694 26462 13746
rect 26514 13694 26526 13746
rect 28578 13694 28590 13746
rect 28642 13694 28654 13746
rect 31266 13694 31278 13746
rect 31330 13694 31342 13746
rect 35410 13694 35422 13746
rect 35474 13694 35486 13746
rect 36642 13694 36654 13746
rect 36706 13694 36718 13746
rect 15934 13682 15986 13694
rect 28366 13682 28418 13694
rect 34526 13682 34578 13694
rect 35982 13682 36034 13694
rect 40350 13682 40402 13694
rect 41246 13746 41298 13758
rect 42018 13694 42030 13746
rect 42082 13694 42094 13746
rect 41246 13682 41298 13694
rect 14254 13634 14306 13646
rect 24782 13634 24834 13646
rect 11666 13582 11678 13634
rect 11730 13582 11742 13634
rect 13794 13582 13806 13634
rect 13858 13582 13870 13634
rect 19842 13582 19854 13634
rect 19906 13582 19918 13634
rect 14254 13570 14306 13582
rect 24782 13570 24834 13582
rect 34302 13634 34354 13646
rect 41794 13582 41806 13634
rect 41858 13582 41870 13634
rect 43138 13582 43150 13634
rect 43202 13582 43214 13634
rect 34302 13570 34354 13582
rect 15598 13522 15650 13534
rect 15598 13458 15650 13470
rect 32174 13522 32226 13534
rect 32174 13458 32226 13470
rect 35422 13522 35474 13534
rect 35422 13458 35474 13470
rect 39678 13522 39730 13534
rect 39678 13458 39730 13470
rect 1344 13354 44576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 44576 13354
rect 1344 13268 44576 13302
rect 19406 13186 19458 13198
rect 36990 13186 37042 13198
rect 26674 13134 26686 13186
rect 26738 13134 26750 13186
rect 19406 13122 19458 13134
rect 36990 13122 37042 13134
rect 37438 13186 37490 13198
rect 37438 13122 37490 13134
rect 20190 13074 20242 13086
rect 15698 13022 15710 13074
rect 15762 13022 15774 13074
rect 17826 13022 17838 13074
rect 17890 13022 17902 13074
rect 19058 13022 19070 13074
rect 19122 13022 19134 13074
rect 20190 13010 20242 13022
rect 20638 13074 20690 13086
rect 22430 13074 22482 13086
rect 29374 13074 29426 13086
rect 21970 13022 21982 13074
rect 22034 13022 22046 13074
rect 26114 13022 26126 13074
rect 26178 13022 26190 13074
rect 20638 13010 20690 13022
rect 22430 13010 22482 13022
rect 29374 13010 29426 13022
rect 30046 13074 30098 13086
rect 30046 13010 30098 13022
rect 31166 13074 31218 13086
rect 31166 13010 31218 13022
rect 32062 13074 32114 13086
rect 37550 13074 37602 13086
rect 34290 13022 34302 13074
rect 34354 13022 34366 13074
rect 36418 13022 36430 13074
rect 36482 13022 36494 13074
rect 42354 13022 42366 13074
rect 42418 13022 42430 13074
rect 43698 13022 43710 13074
rect 43762 13022 43774 13074
rect 32062 13010 32114 13022
rect 37550 13010 37602 13022
rect 12798 12962 12850 12974
rect 18062 12962 18114 12974
rect 14354 12910 14366 12962
rect 14418 12910 14430 12962
rect 14914 12910 14926 12962
rect 14978 12910 14990 12962
rect 12798 12898 12850 12910
rect 18062 12898 18114 12910
rect 18398 12962 18450 12974
rect 18398 12898 18450 12910
rect 18734 12962 18786 12974
rect 27022 12962 27074 12974
rect 25778 12910 25790 12962
rect 25842 12910 25854 12962
rect 18734 12898 18786 12910
rect 27022 12898 27074 12910
rect 32622 12962 32674 12974
rect 32622 12898 32674 12910
rect 33182 12962 33234 12974
rect 38222 12962 38274 12974
rect 33618 12910 33630 12962
rect 33682 12910 33694 12962
rect 38658 12910 38670 12962
rect 38722 12910 38734 12962
rect 42130 12910 42142 12962
rect 42194 12910 42206 12962
rect 33182 12898 33234 12910
rect 38222 12898 38274 12910
rect 12462 12850 12514 12862
rect 12462 12786 12514 12798
rect 19182 12850 19234 12862
rect 19182 12786 19234 12798
rect 21646 12850 21698 12862
rect 21646 12786 21698 12798
rect 21870 12850 21922 12862
rect 21870 12786 21922 12798
rect 27246 12850 27298 12862
rect 27246 12786 27298 12798
rect 32958 12850 33010 12862
rect 32958 12786 33010 12798
rect 37102 12850 37154 12862
rect 37102 12786 37154 12798
rect 43038 12850 43090 12862
rect 43038 12786 43090 12798
rect 44158 12850 44210 12862
rect 44158 12786 44210 12798
rect 14590 12738 14642 12750
rect 14590 12674 14642 12686
rect 18286 12738 18338 12750
rect 18286 12674 18338 12686
rect 22878 12738 22930 12750
rect 22878 12674 22930 12686
rect 27694 12738 27746 12750
rect 27694 12674 27746 12686
rect 28142 12738 28194 12750
rect 28142 12674 28194 12686
rect 28590 12738 28642 12750
rect 28590 12674 28642 12686
rect 31502 12738 31554 12750
rect 31502 12674 31554 12686
rect 32846 12738 32898 12750
rect 41694 12738 41746 12750
rect 41122 12686 41134 12738
rect 41186 12686 41198 12738
rect 32846 12674 32898 12686
rect 41694 12674 41746 12686
rect 1344 12570 44576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 44576 12570
rect 1344 12484 44576 12518
rect 17502 12402 17554 12414
rect 17502 12338 17554 12350
rect 19406 12402 19458 12414
rect 19406 12338 19458 12350
rect 21758 12402 21810 12414
rect 21758 12338 21810 12350
rect 22990 12402 23042 12414
rect 22990 12338 23042 12350
rect 23662 12402 23714 12414
rect 23662 12338 23714 12350
rect 27022 12402 27074 12414
rect 27022 12338 27074 12350
rect 30270 12402 30322 12414
rect 30270 12338 30322 12350
rect 30606 12402 30658 12414
rect 30606 12338 30658 12350
rect 36766 12402 36818 12414
rect 36766 12338 36818 12350
rect 36990 12402 37042 12414
rect 36990 12338 37042 12350
rect 38782 12402 38834 12414
rect 38782 12338 38834 12350
rect 41134 12402 41186 12414
rect 41134 12338 41186 12350
rect 44270 12402 44322 12414
rect 44270 12338 44322 12350
rect 19854 12290 19906 12302
rect 22094 12290 22146 12302
rect 14690 12238 14702 12290
rect 14754 12238 14766 12290
rect 18050 12238 18062 12290
rect 18114 12238 18126 12290
rect 18386 12238 18398 12290
rect 18450 12238 18462 12290
rect 21410 12238 21422 12290
rect 21474 12238 21486 12290
rect 19854 12226 19906 12238
rect 22094 12226 22146 12238
rect 22430 12290 22482 12302
rect 22430 12226 22482 12238
rect 28142 12290 28194 12302
rect 30942 12290 30994 12302
rect 29138 12238 29150 12290
rect 29202 12238 29214 12290
rect 29698 12238 29710 12290
rect 29762 12238 29774 12290
rect 28142 12226 28194 12238
rect 30942 12226 30994 12238
rect 38894 12290 38946 12302
rect 38894 12226 38946 12238
rect 41470 12290 41522 12302
rect 41470 12226 41522 12238
rect 43262 12290 43314 12302
rect 43262 12226 43314 12238
rect 28590 12178 28642 12190
rect 14018 12126 14030 12178
rect 14082 12126 14094 12178
rect 19170 12126 19182 12178
rect 19234 12126 19246 12178
rect 27906 12126 27918 12178
rect 27970 12126 27982 12178
rect 28590 12114 28642 12126
rect 28926 12178 28978 12190
rect 28926 12114 28978 12126
rect 32062 12178 32114 12190
rect 32062 12114 32114 12126
rect 32286 12178 32338 12190
rect 32286 12114 32338 12126
rect 32622 12178 32674 12190
rect 36318 12178 36370 12190
rect 33058 12126 33070 12178
rect 33122 12126 33134 12178
rect 32622 12114 32674 12126
rect 36318 12114 36370 12126
rect 36542 12178 36594 12190
rect 42018 12126 42030 12178
rect 42082 12126 42094 12178
rect 43474 12126 43486 12178
rect 43538 12126 43550 12178
rect 36542 12114 36594 12126
rect 22878 12066 22930 12078
rect 16818 12014 16830 12066
rect 16882 12014 16894 12066
rect 22878 12002 22930 12014
rect 27470 12066 27522 12078
rect 27470 12002 27522 12014
rect 32398 12066 32450 12078
rect 36878 12066 36930 12078
rect 33842 12014 33854 12066
rect 33906 12014 33918 12066
rect 35970 12014 35982 12066
rect 36034 12014 36046 12066
rect 32398 12002 32450 12014
rect 36878 12002 36930 12014
rect 38110 12066 38162 12078
rect 42354 12014 42366 12066
rect 42418 12014 42430 12066
rect 38110 12002 38162 12014
rect 17838 11954 17890 11966
rect 17838 11890 17890 11902
rect 22766 11954 22818 11966
rect 38222 11954 38274 11966
rect 26898 11902 26910 11954
rect 26962 11951 26974 11954
rect 27458 11951 27470 11954
rect 26962 11905 27470 11951
rect 26962 11902 26974 11905
rect 27458 11902 27470 11905
rect 27522 11902 27534 11954
rect 42578 11902 42590 11954
rect 42642 11902 42654 11954
rect 22766 11890 22818 11902
rect 38222 11890 38274 11902
rect 1344 11786 44576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 44576 11786
rect 1344 11700 44576 11734
rect 21758 11618 21810 11630
rect 21758 11554 21810 11566
rect 22094 11618 22146 11630
rect 22094 11554 22146 11566
rect 27694 11618 27746 11630
rect 27694 11554 27746 11566
rect 38222 11618 38274 11630
rect 38222 11554 38274 11566
rect 13582 11506 13634 11518
rect 20750 11506 20802 11518
rect 31166 11506 31218 11518
rect 36430 11506 36482 11518
rect 16146 11454 16158 11506
rect 16210 11454 16222 11506
rect 18274 11454 18286 11506
rect 18338 11454 18350 11506
rect 25666 11454 25678 11506
rect 25730 11454 25742 11506
rect 33842 11454 33854 11506
rect 33906 11454 33918 11506
rect 35970 11454 35982 11506
rect 36034 11454 36046 11506
rect 13582 11442 13634 11454
rect 20750 11442 20802 11454
rect 31166 11442 31218 11454
rect 36430 11442 36482 11454
rect 38110 11506 38162 11518
rect 38110 11442 38162 11454
rect 29822 11394 29874 11406
rect 37102 11394 37154 11406
rect 19058 11342 19070 11394
rect 19122 11342 19134 11394
rect 22418 11342 22430 11394
rect 22482 11342 22494 11394
rect 22754 11342 22766 11394
rect 22818 11342 22830 11394
rect 32610 11342 32622 11394
rect 32674 11342 32686 11394
rect 33058 11342 33070 11394
rect 33122 11342 33134 11394
rect 29822 11330 29874 11342
rect 37102 11330 37154 11342
rect 37326 11394 37378 11406
rect 37326 11330 37378 11342
rect 37550 11394 37602 11406
rect 37550 11330 37602 11342
rect 37774 11394 37826 11406
rect 37774 11330 37826 11342
rect 38894 11394 38946 11406
rect 42590 11394 42642 11406
rect 39218 11342 39230 11394
rect 39282 11342 39294 11394
rect 38894 11330 38946 11342
rect 42590 11330 42642 11342
rect 12350 11282 12402 11294
rect 12350 11218 12402 11230
rect 21534 11282 21586 11294
rect 26574 11282 26626 11294
rect 23538 11230 23550 11282
rect 23602 11230 23614 11282
rect 21534 11218 21586 11230
rect 26574 11218 26626 11230
rect 27358 11282 27410 11294
rect 29486 11282 29538 11294
rect 28018 11230 28030 11282
rect 28082 11230 28094 11282
rect 28466 11230 28478 11282
rect 28530 11230 28542 11282
rect 27358 11218 27410 11230
rect 29486 11218 29538 11230
rect 30494 11282 30546 11294
rect 30494 11218 30546 11230
rect 30606 11282 30658 11294
rect 30606 11218 30658 11230
rect 12014 11170 12066 11182
rect 12014 11106 12066 11118
rect 12238 11170 12290 11182
rect 12238 11106 12290 11118
rect 12798 11170 12850 11182
rect 12798 11106 12850 11118
rect 21646 11170 21698 11182
rect 21646 11106 21698 11118
rect 22206 11170 22258 11182
rect 22206 11106 22258 11118
rect 26910 11170 26962 11182
rect 26910 11106 26962 11118
rect 29150 11170 29202 11182
rect 30830 11170 30882 11182
rect 30146 11118 30158 11170
rect 30210 11118 30222 11170
rect 29150 11106 29202 11118
rect 30830 11106 30882 11118
rect 32398 11170 32450 11182
rect 32398 11106 32450 11118
rect 36318 11170 36370 11182
rect 36318 11106 36370 11118
rect 37214 11170 37266 11182
rect 42366 11170 42418 11182
rect 41794 11118 41806 11170
rect 41858 11118 41870 11170
rect 37214 11106 37266 11118
rect 42366 11106 42418 11118
rect 42926 11170 42978 11182
rect 42926 11106 42978 11118
rect 1344 11002 44576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 44576 11002
rect 1344 10916 44576 10950
rect 13134 10834 13186 10846
rect 13134 10770 13186 10782
rect 15262 10834 15314 10846
rect 15262 10770 15314 10782
rect 15822 10834 15874 10846
rect 15822 10770 15874 10782
rect 23662 10834 23714 10846
rect 23662 10770 23714 10782
rect 31278 10834 31330 10846
rect 31278 10770 31330 10782
rect 33966 10834 34018 10846
rect 33966 10770 34018 10782
rect 34078 10834 34130 10846
rect 34078 10770 34130 10782
rect 35198 10834 35250 10846
rect 38334 10834 38386 10846
rect 36082 10782 36094 10834
rect 36146 10782 36158 10834
rect 35198 10770 35250 10782
rect 38334 10770 38386 10782
rect 38446 10834 38498 10846
rect 38446 10770 38498 10782
rect 41358 10834 41410 10846
rect 41358 10770 41410 10782
rect 11006 10722 11058 10734
rect 11006 10658 11058 10670
rect 11902 10722 11954 10734
rect 13806 10722 13858 10734
rect 12786 10670 12798 10722
rect 12850 10670 12862 10722
rect 11902 10658 11954 10670
rect 13806 10658 13858 10670
rect 15374 10722 15426 10734
rect 15374 10658 15426 10670
rect 21646 10722 21698 10734
rect 21646 10658 21698 10670
rect 22206 10722 22258 10734
rect 22206 10658 22258 10670
rect 23214 10722 23266 10734
rect 23214 10658 23266 10670
rect 24558 10722 24610 10734
rect 31054 10722 31106 10734
rect 28354 10670 28366 10722
rect 28418 10670 28430 10722
rect 24558 10658 24610 10670
rect 31054 10658 31106 10670
rect 31726 10722 31778 10734
rect 31726 10658 31778 10670
rect 35310 10722 35362 10734
rect 35310 10658 35362 10670
rect 35534 10722 35586 10734
rect 35970 10670 35982 10722
rect 36034 10670 36046 10722
rect 37426 10670 37438 10722
rect 37490 10670 37502 10722
rect 41010 10670 41022 10722
rect 41074 10670 41086 10722
rect 35534 10658 35586 10670
rect 11230 10610 11282 10622
rect 11230 10546 11282 10558
rect 11678 10610 11730 10622
rect 11678 10546 11730 10558
rect 12126 10610 12178 10622
rect 12126 10546 12178 10558
rect 12574 10610 12626 10622
rect 12574 10546 12626 10558
rect 14030 10610 14082 10622
rect 14030 10546 14082 10558
rect 14478 10610 14530 10622
rect 14478 10546 14530 10558
rect 15038 10610 15090 10622
rect 21870 10610 21922 10622
rect 21186 10558 21198 10610
rect 21250 10558 21262 10610
rect 15038 10546 15090 10558
rect 21870 10546 21922 10558
rect 22766 10610 22818 10622
rect 22766 10546 22818 10558
rect 22878 10610 22930 10622
rect 22878 10546 22930 10558
rect 23438 10610 23490 10622
rect 23438 10546 23490 10558
rect 23774 10610 23826 10622
rect 23774 10546 23826 10558
rect 23998 10610 24050 10622
rect 30830 10610 30882 10622
rect 27682 10558 27694 10610
rect 27746 10558 27758 10610
rect 23998 10546 24050 10558
rect 30830 10546 30882 10558
rect 34302 10610 34354 10622
rect 35086 10610 35138 10622
rect 36990 10610 37042 10622
rect 38110 10610 38162 10622
rect 34514 10558 34526 10610
rect 34578 10558 34590 10610
rect 34850 10558 34862 10610
rect 34914 10558 34926 10610
rect 35858 10558 35870 10610
rect 35922 10558 35934 10610
rect 37874 10558 37886 10610
rect 37938 10558 37950 10610
rect 34302 10546 34354 10558
rect 35086 10546 35138 10558
rect 36990 10546 37042 10558
rect 38110 10546 38162 10558
rect 11118 10498 11170 10510
rect 11118 10434 11170 10446
rect 12014 10498 12066 10510
rect 12014 10434 12066 10446
rect 13918 10498 13970 10510
rect 22094 10498 22146 10510
rect 18386 10446 18398 10498
rect 18450 10446 18462 10498
rect 20514 10446 20526 10498
rect 20578 10446 20590 10498
rect 13918 10434 13970 10446
rect 22094 10434 22146 10446
rect 23102 10498 23154 10510
rect 30942 10498 30994 10510
rect 30482 10446 30494 10498
rect 30546 10446 30558 10498
rect 23102 10434 23154 10446
rect 30942 10434 30994 10446
rect 31838 10498 31890 10510
rect 31838 10434 31890 10446
rect 34190 10498 34242 10510
rect 34190 10434 34242 10446
rect 38222 10498 38274 10510
rect 38222 10434 38274 10446
rect 41806 10498 41858 10510
rect 41806 10434 41858 10446
rect 24446 10386 24498 10398
rect 24446 10322 24498 10334
rect 41694 10386 41746 10398
rect 41694 10322 41746 10334
rect 1344 10218 44576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 44576 10218
rect 1344 10132 44576 10166
rect 18734 10050 18786 10062
rect 18734 9986 18786 9998
rect 37438 10050 37490 10062
rect 37438 9986 37490 9998
rect 37662 10050 37714 10062
rect 37662 9986 37714 9998
rect 18846 9938 18898 9950
rect 10098 9886 10110 9938
rect 10162 9886 10174 9938
rect 12226 9886 12238 9938
rect 12290 9886 12302 9938
rect 14242 9886 14254 9938
rect 14306 9886 14318 9938
rect 16370 9886 16382 9938
rect 16434 9886 16446 9938
rect 17938 9886 17950 9938
rect 18002 9886 18014 9938
rect 18846 9874 18898 9886
rect 21422 9938 21474 9950
rect 38334 9938 38386 9950
rect 23426 9886 23438 9938
rect 23490 9886 23502 9938
rect 25554 9886 25566 9938
rect 25618 9886 25630 9938
rect 29922 9886 29934 9938
rect 29986 9886 29998 9938
rect 32050 9886 32062 9938
rect 32114 9886 32126 9938
rect 38658 9886 38670 9938
rect 38722 9886 38734 9938
rect 44034 9886 44046 9938
rect 44098 9886 44110 9938
rect 21422 9874 21474 9886
rect 38334 9874 38386 9886
rect 12574 9826 12626 9838
rect 9426 9774 9438 9826
rect 9490 9774 9502 9826
rect 12574 9762 12626 9774
rect 12910 9826 12962 9838
rect 21534 9826 21586 9838
rect 13458 9774 13470 9826
rect 13522 9774 13534 9826
rect 17714 9774 17726 9826
rect 17778 9774 17790 9826
rect 12910 9762 12962 9774
rect 21534 9762 21586 9774
rect 21870 9826 21922 9838
rect 37214 9826 37266 9838
rect 22754 9774 22766 9826
rect 22818 9774 22830 9826
rect 29138 9774 29150 9826
rect 29202 9774 29214 9826
rect 34514 9774 34526 9826
rect 34578 9774 34590 9826
rect 35298 9774 35310 9826
rect 35362 9774 35374 9826
rect 35634 9774 35646 9826
rect 35698 9774 35710 9826
rect 21870 9762 21922 9774
rect 37214 9762 37266 9774
rect 38110 9826 38162 9838
rect 38882 9774 38894 9826
rect 38946 9774 38958 9826
rect 40674 9774 40686 9826
rect 40738 9774 40750 9826
rect 41234 9774 41246 9826
rect 41298 9774 41310 9826
rect 38110 9762 38162 9774
rect 12798 9714 12850 9726
rect 12798 9650 12850 9662
rect 18398 9714 18450 9726
rect 18398 9650 18450 9662
rect 20638 9714 20690 9726
rect 20638 9650 20690 9662
rect 21310 9714 21362 9726
rect 21310 9650 21362 9662
rect 34638 9714 34690 9726
rect 36990 9714 37042 9726
rect 35858 9662 35870 9714
rect 35922 9662 35934 9714
rect 43474 9662 43486 9714
rect 43538 9662 43550 9714
rect 34638 9650 34690 9662
rect 36990 9650 37042 9662
rect 20750 9602 20802 9614
rect 20750 9538 20802 9550
rect 32510 9602 32562 9614
rect 32510 9538 32562 9550
rect 1344 9434 44576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 44576 9434
rect 1344 9348 44576 9382
rect 15822 9266 15874 9278
rect 15822 9202 15874 9214
rect 23102 9266 23154 9278
rect 23102 9202 23154 9214
rect 25454 9266 25506 9278
rect 25454 9202 25506 9214
rect 33182 9266 33234 9278
rect 33182 9202 33234 9214
rect 33742 9266 33794 9278
rect 33742 9202 33794 9214
rect 34974 9266 35026 9278
rect 34974 9202 35026 9214
rect 35086 9266 35138 9278
rect 35086 9202 35138 9214
rect 35198 9266 35250 9278
rect 35198 9202 35250 9214
rect 38670 9266 38722 9278
rect 38670 9202 38722 9214
rect 43374 9266 43426 9278
rect 43374 9202 43426 9214
rect 44158 9266 44210 9278
rect 44158 9202 44210 9214
rect 24334 9154 24386 9166
rect 11666 9102 11678 9154
rect 11730 9102 11742 9154
rect 14018 9102 14030 9154
rect 14082 9102 14094 9154
rect 19394 9102 19406 9154
rect 19458 9102 19470 9154
rect 20626 9102 20638 9154
rect 20690 9102 20702 9154
rect 24334 9090 24386 9102
rect 25790 9154 25842 9166
rect 32174 9154 32226 9166
rect 27682 9102 27694 9154
rect 27746 9102 27758 9154
rect 30930 9102 30942 9154
rect 30994 9102 31006 9154
rect 31378 9102 31390 9154
rect 31442 9102 31454 9154
rect 25790 9090 25842 9102
rect 32174 9090 32226 9102
rect 33070 9154 33122 9166
rect 33070 9090 33122 9102
rect 36542 9154 36594 9166
rect 42478 9154 42530 9166
rect 37874 9102 37886 9154
rect 37938 9102 37950 9154
rect 36542 9090 36594 9102
rect 42478 9090 42530 9102
rect 13022 9042 13074 9054
rect 12450 8990 12462 9042
rect 12514 8990 12526 9042
rect 12786 8990 12798 9042
rect 12850 8990 12862 9042
rect 13022 8978 13074 8990
rect 13134 9042 13186 9054
rect 13134 8978 13186 8990
rect 13246 9042 13298 9054
rect 23214 9042 23266 9054
rect 25678 9042 25730 9054
rect 30606 9042 30658 9054
rect 13458 8990 13470 9042
rect 13522 8990 13534 9042
rect 14130 8990 14142 9042
rect 14194 8990 14206 9042
rect 14914 8990 14926 9042
rect 14978 8990 14990 9042
rect 15250 8990 15262 9042
rect 15314 8990 15326 9042
rect 18162 8990 18174 9042
rect 18226 8990 18238 9042
rect 18722 8990 18734 9042
rect 18786 8990 18798 9042
rect 19506 8990 19518 9042
rect 19570 8990 19582 9042
rect 19842 8990 19854 9042
rect 19906 8990 19918 9042
rect 25218 8990 25230 9042
rect 25282 8990 25294 9042
rect 26898 8990 26910 9042
rect 26962 8990 26974 9042
rect 13246 8978 13298 8990
rect 23214 8978 23266 8990
rect 25678 8978 25730 8990
rect 30606 8978 30658 8990
rect 31838 9042 31890 9054
rect 31838 8978 31890 8990
rect 33406 9042 33458 9054
rect 36318 9042 36370 9054
rect 38558 9042 38610 9054
rect 35858 8990 35870 9042
rect 35922 8990 35934 9042
rect 36642 8990 36654 9042
rect 36706 8990 36718 9042
rect 37202 8990 37214 9042
rect 37266 8990 37278 9042
rect 38322 8990 38334 9042
rect 38386 8990 38398 9042
rect 33406 8978 33458 8990
rect 36318 8978 36370 8990
rect 38558 8978 38610 8990
rect 38782 9042 38834 9054
rect 38994 8990 39006 9042
rect 39058 8990 39070 9042
rect 42690 8990 42702 9042
rect 42754 8990 42766 9042
rect 38782 8978 38834 8990
rect 15934 8930 15986 8942
rect 34750 8930 34802 8942
rect 9538 8878 9550 8930
rect 9602 8878 9614 8930
rect 22754 8878 22766 8930
rect 22818 8878 22830 8930
rect 25778 8878 25790 8930
rect 25842 8878 25854 8930
rect 29810 8878 29822 8930
rect 29874 8878 29886 8930
rect 15934 8866 15986 8878
rect 34750 8866 34802 8878
rect 39454 8930 39506 8942
rect 39454 8866 39506 8878
rect 41022 8930 41074 8942
rect 43698 8878 43710 8930
rect 43762 8878 43774 8930
rect 41022 8866 41074 8878
rect 15598 8818 15650 8830
rect 24222 8818 24274 8830
rect 18386 8766 18398 8818
rect 18450 8766 18462 8818
rect 15598 8754 15650 8766
rect 24222 8754 24274 8766
rect 30270 8818 30322 8830
rect 30270 8754 30322 8766
rect 34526 8818 34578 8830
rect 34526 8754 34578 8766
rect 39342 8818 39394 8830
rect 39342 8754 39394 8766
rect 40910 8818 40962 8830
rect 40910 8754 40962 8766
rect 1344 8650 44576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 44576 8650
rect 1344 8564 44576 8598
rect 12798 8482 12850 8494
rect 25678 8482 25730 8494
rect 17938 8430 17950 8482
rect 18002 8430 18014 8482
rect 42690 8430 42702 8482
rect 42754 8430 42766 8482
rect 12798 8418 12850 8430
rect 25678 8418 25730 8430
rect 11230 8370 11282 8382
rect 14030 8370 14082 8382
rect 29262 8370 29314 8382
rect 35758 8370 35810 8382
rect 12114 8318 12126 8370
rect 12178 8318 12190 8370
rect 18498 8318 18510 8370
rect 18562 8318 18574 8370
rect 20290 8318 20302 8370
rect 20354 8318 20366 8370
rect 21410 8318 21422 8370
rect 21474 8318 21486 8370
rect 22530 8318 22542 8370
rect 22594 8318 22606 8370
rect 34850 8318 34862 8370
rect 34914 8318 34926 8370
rect 42130 8318 42142 8370
rect 42194 8318 42206 8370
rect 42802 8318 42814 8370
rect 42866 8318 42878 8370
rect 11230 8306 11282 8318
rect 14030 8306 14082 8318
rect 29262 8306 29314 8318
rect 35758 8306 35810 8318
rect 11342 8258 11394 8270
rect 11342 8194 11394 8206
rect 11902 8258 11954 8270
rect 11902 8194 11954 8206
rect 12238 8258 12290 8270
rect 12238 8194 12290 8206
rect 12686 8258 12738 8270
rect 14142 8258 14194 8270
rect 17390 8258 17442 8270
rect 18846 8258 18898 8270
rect 13682 8206 13694 8258
rect 13746 8206 13758 8258
rect 16034 8206 16046 8258
rect 16098 8206 16110 8258
rect 17042 8206 17054 8258
rect 17106 8206 17118 8258
rect 17602 8206 17614 8258
rect 17666 8206 17678 8258
rect 12686 8194 12738 8206
rect 14142 8194 14194 8206
rect 17390 8194 17442 8206
rect 18846 8194 18898 8206
rect 19966 8258 20018 8270
rect 21758 8258 21810 8270
rect 20402 8206 20414 8258
rect 20466 8206 20478 8258
rect 21298 8206 21310 8258
rect 21362 8206 21374 8258
rect 19966 8194 20018 8206
rect 21758 8194 21810 8206
rect 22430 8258 22482 8270
rect 22430 8194 22482 8206
rect 22878 8258 22930 8270
rect 22878 8194 22930 8206
rect 25566 8258 25618 8270
rect 25566 8194 25618 8206
rect 29934 8258 29986 8270
rect 29934 8194 29986 8206
rect 30270 8258 30322 8270
rect 30270 8194 30322 8206
rect 30606 8258 30658 8270
rect 35198 8258 35250 8270
rect 32050 8206 32062 8258
rect 32114 8206 32126 8258
rect 30606 8194 30658 8206
rect 35198 8194 35250 8206
rect 35422 8258 35474 8270
rect 35422 8194 35474 8206
rect 35870 8258 35922 8270
rect 35870 8194 35922 8206
rect 38894 8258 38946 8270
rect 39330 8206 39342 8258
rect 39394 8206 39406 8258
rect 43138 8206 43150 8258
rect 43202 8206 43214 8258
rect 38894 8194 38946 8206
rect 10894 8146 10946 8158
rect 10894 8082 10946 8094
rect 11678 8146 11730 8158
rect 11678 8082 11730 8094
rect 14366 8146 14418 8158
rect 19070 8146 19122 8158
rect 15810 8094 15822 8146
rect 15874 8094 15886 8146
rect 14366 8082 14418 8094
rect 19070 8082 19122 8094
rect 19742 8146 19794 8158
rect 19742 8082 19794 8094
rect 21982 8146 22034 8158
rect 21982 8082 22034 8094
rect 22542 8146 22594 8158
rect 22542 8082 22594 8094
rect 31278 8146 31330 8158
rect 32722 8094 32734 8146
rect 32786 8094 32798 8146
rect 31278 8082 31330 8094
rect 10782 8034 10834 8046
rect 10782 7970 10834 7982
rect 12126 8034 12178 8046
rect 12126 7970 12178 7982
rect 13918 8034 13970 8046
rect 13918 7970 13970 7982
rect 18510 8034 18562 8046
rect 18510 7970 18562 7982
rect 18622 8034 18674 8046
rect 18622 7970 18674 7982
rect 20190 8034 20242 8046
rect 20190 7970 20242 7982
rect 21534 8034 21586 8046
rect 21534 7970 21586 7982
rect 22766 8034 22818 8046
rect 22766 7970 22818 7982
rect 29598 8034 29650 8046
rect 29598 7970 29650 7982
rect 30382 8034 30434 8046
rect 30382 7970 30434 7982
rect 30830 8034 30882 8046
rect 30830 7970 30882 7982
rect 30942 8034 30994 8046
rect 30942 7970 30994 7982
rect 31054 8034 31106 8046
rect 31054 7970 31106 7982
rect 35646 8034 35698 8046
rect 41794 7982 41806 8034
rect 41858 7982 41870 8034
rect 35646 7970 35698 7982
rect 1344 7866 44576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 44576 7866
rect 1344 7780 44576 7814
rect 19518 7698 19570 7710
rect 13682 7646 13694 7698
rect 13746 7646 13758 7698
rect 18834 7646 18846 7698
rect 18898 7646 18910 7698
rect 19518 7634 19570 7646
rect 19742 7698 19794 7710
rect 19742 7634 19794 7646
rect 22654 7698 22706 7710
rect 22654 7634 22706 7646
rect 24670 7698 24722 7710
rect 28814 7698 28866 7710
rect 28242 7646 28254 7698
rect 28306 7646 28318 7698
rect 24670 7634 24722 7646
rect 28814 7634 28866 7646
rect 32398 7698 32450 7710
rect 32398 7634 32450 7646
rect 33182 7698 33234 7710
rect 33182 7634 33234 7646
rect 33294 7698 33346 7710
rect 33294 7634 33346 7646
rect 34078 7698 34130 7710
rect 34078 7634 34130 7646
rect 35086 7698 35138 7710
rect 35086 7634 35138 7646
rect 35870 7698 35922 7710
rect 40910 7698 40962 7710
rect 39890 7646 39902 7698
rect 39954 7646 39966 7698
rect 35870 7634 35922 7646
rect 40910 7634 40962 7646
rect 43038 7698 43090 7710
rect 43038 7634 43090 7646
rect 24558 7586 24610 7598
rect 32622 7586 32674 7598
rect 17490 7534 17502 7586
rect 17554 7534 17566 7586
rect 18946 7534 18958 7586
rect 19010 7534 19022 7586
rect 29810 7534 29822 7586
rect 29874 7534 29886 7586
rect 24558 7522 24610 7534
rect 32622 7522 32674 7534
rect 33518 7586 33570 7598
rect 33518 7522 33570 7534
rect 35758 7586 35810 7598
rect 35758 7522 35810 7534
rect 10782 7474 10834 7486
rect 16830 7474 16882 7486
rect 11218 7422 11230 7474
rect 11282 7422 11294 7474
rect 10782 7410 10834 7422
rect 16830 7410 16882 7422
rect 17950 7474 18002 7486
rect 19630 7474 19682 7486
rect 18498 7422 18510 7474
rect 18562 7422 18574 7474
rect 17950 7410 18002 7422
rect 19630 7410 19682 7422
rect 19854 7474 19906 7486
rect 19854 7410 19906 7422
rect 19966 7474 20018 7486
rect 19966 7410 20018 7422
rect 22318 7474 22370 7486
rect 32286 7474 32338 7486
rect 25218 7422 25230 7474
rect 25282 7422 25294 7474
rect 25666 7422 25678 7474
rect 25730 7422 25742 7474
rect 29138 7422 29150 7474
rect 29202 7422 29214 7474
rect 22318 7410 22370 7422
rect 32286 7410 32338 7422
rect 33070 7474 33122 7486
rect 33070 7410 33122 7422
rect 34862 7474 34914 7486
rect 34862 7410 34914 7422
rect 34974 7474 35026 7486
rect 34974 7410 35026 7422
rect 35198 7474 35250 7486
rect 42702 7474 42754 7486
rect 35410 7422 35422 7474
rect 35474 7422 35486 7474
rect 36866 7422 36878 7474
rect 36930 7422 36942 7474
rect 37426 7422 37438 7474
rect 37490 7422 37502 7474
rect 42242 7422 42254 7474
rect 42306 7422 42318 7474
rect 43250 7422 43262 7474
rect 43314 7422 43326 7474
rect 35198 7410 35250 7422
rect 42702 7410 42754 7422
rect 16718 7362 16770 7374
rect 14018 7310 14030 7362
rect 14082 7310 14094 7362
rect 16718 7298 16770 7310
rect 22766 7362 22818 7374
rect 33966 7362 34018 7374
rect 31938 7310 31950 7362
rect 32002 7310 32014 7362
rect 22766 7298 22818 7310
rect 33966 7298 34018 7310
rect 41022 7362 41074 7374
rect 42018 7310 42030 7362
rect 42082 7310 42094 7362
rect 41022 7298 41074 7310
rect 22206 7250 22258 7262
rect 22206 7186 22258 7198
rect 40462 7250 40514 7262
rect 40462 7186 40514 7198
rect 1344 7082 44576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 44576 7082
rect 1344 6996 44576 7030
rect 16830 6914 16882 6926
rect 16830 6850 16882 6862
rect 24894 6914 24946 6926
rect 24894 6850 24946 6862
rect 43374 6914 43426 6926
rect 43374 6850 43426 6862
rect 28578 6750 28590 6802
rect 28642 6750 28654 6802
rect 30818 6750 30830 6802
rect 30882 6750 30894 6802
rect 32946 6750 32958 6802
rect 33010 6750 33022 6802
rect 36194 6750 36206 6802
rect 36258 6750 36270 6802
rect 38658 6750 38670 6802
rect 38722 6750 38734 6802
rect 8878 6690 8930 6702
rect 12350 6690 12402 6702
rect 9314 6638 9326 6690
rect 9378 6638 9390 6690
rect 8878 6626 8930 6638
rect 12350 6626 12402 6638
rect 12574 6690 12626 6702
rect 12574 6626 12626 6638
rect 12686 6690 12738 6702
rect 20302 6690 20354 6702
rect 19954 6638 19966 6690
rect 20018 6638 20030 6690
rect 12686 6626 12738 6638
rect 20302 6626 20354 6638
rect 21422 6690 21474 6702
rect 36990 6690 37042 6702
rect 21858 6638 21870 6690
rect 21922 6638 21934 6690
rect 25106 6638 25118 6690
rect 25170 6638 25182 6690
rect 25554 6638 25566 6690
rect 25618 6638 25630 6690
rect 30034 6638 30046 6690
rect 30098 6638 30110 6690
rect 33282 6638 33294 6690
rect 33346 6638 33358 6690
rect 38882 6638 38894 6690
rect 38946 6638 38958 6690
rect 39778 6638 39790 6690
rect 39842 6638 39854 6690
rect 40338 6638 40350 6690
rect 40402 6638 40414 6690
rect 21422 6626 21474 6638
rect 36990 6626 37042 6638
rect 13806 6578 13858 6590
rect 13806 6514 13858 6526
rect 14142 6578 14194 6590
rect 14142 6514 14194 6526
rect 14478 6578 14530 6590
rect 14478 6514 14530 6526
rect 15262 6578 15314 6590
rect 15262 6514 15314 6526
rect 16606 6578 16658 6590
rect 37102 6578 37154 6590
rect 34066 6526 34078 6578
rect 34130 6526 34142 6578
rect 16606 6514 16658 6526
rect 37102 6514 37154 6526
rect 37438 6578 37490 6590
rect 37438 6514 37490 6526
rect 39454 6578 39506 6590
rect 43598 6578 43650 6590
rect 42578 6526 42590 6578
rect 42642 6526 42654 6578
rect 39454 6514 39506 6526
rect 43598 6514 43650 6526
rect 43934 6578 43986 6590
rect 43934 6514 43986 6526
rect 14814 6466 14866 6478
rect 11778 6414 11790 6466
rect 11842 6414 11854 6466
rect 14814 6402 14866 6414
rect 15150 6466 15202 6478
rect 15150 6402 15202 6414
rect 16494 6466 16546 6478
rect 37550 6466 37602 6478
rect 17602 6414 17614 6466
rect 17666 6414 17678 6466
rect 24322 6414 24334 6466
rect 24386 6414 24398 6466
rect 28130 6414 28142 6466
rect 28194 6414 28206 6466
rect 16494 6402 16546 6414
rect 37550 6402 37602 6414
rect 1344 6298 44576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 44576 6298
rect 1344 6212 44576 6246
rect 12238 6130 12290 6142
rect 12238 6066 12290 6078
rect 13134 6130 13186 6142
rect 18174 6130 18226 6142
rect 16370 6078 16382 6130
rect 16434 6078 16446 6130
rect 13134 6066 13186 6078
rect 18174 6066 18226 6078
rect 18846 6130 18898 6142
rect 18846 6066 18898 6078
rect 23774 6130 23826 6142
rect 23774 6066 23826 6078
rect 26910 6130 26962 6142
rect 26910 6066 26962 6078
rect 28478 6130 28530 6142
rect 28478 6066 28530 6078
rect 29150 6130 29202 6142
rect 29150 6066 29202 6078
rect 32174 6130 32226 6142
rect 32174 6066 32226 6078
rect 32622 6130 32674 6142
rect 32622 6066 32674 6078
rect 33070 6130 33122 6142
rect 33070 6066 33122 6078
rect 33182 6130 33234 6142
rect 33182 6066 33234 6078
rect 33294 6130 33346 6142
rect 33294 6066 33346 6078
rect 34190 6130 34242 6142
rect 41470 6130 41522 6142
rect 37650 6078 37662 6130
rect 37714 6078 37726 6130
rect 34190 6066 34242 6078
rect 41470 6066 41522 6078
rect 43598 6130 43650 6142
rect 43598 6066 43650 6078
rect 43822 6130 43874 6142
rect 43822 6066 43874 6078
rect 17726 6018 17778 6030
rect 25230 6018 25282 6030
rect 22978 5966 22990 6018
rect 23042 5966 23054 6018
rect 17726 5954 17778 5966
rect 25230 5954 25282 5966
rect 31278 6018 31330 6030
rect 31278 5954 31330 5966
rect 31614 6018 31666 6030
rect 31614 5954 31666 5966
rect 34302 6018 34354 6030
rect 34302 5954 34354 5966
rect 42926 6018 42978 6030
rect 42926 5954 42978 5966
rect 44158 6018 44210 6030
rect 44158 5954 44210 5966
rect 17838 5906 17890 5918
rect 27246 5906 27298 5918
rect 34750 5906 34802 5918
rect 38670 5906 38722 5918
rect 40910 5906 40962 5918
rect 12450 5854 12462 5906
rect 12514 5854 12526 5906
rect 13346 5854 13358 5906
rect 13410 5854 13422 5906
rect 13906 5854 13918 5906
rect 13970 5854 13982 5906
rect 18386 5854 18398 5906
rect 18450 5854 18462 5906
rect 20178 5854 20190 5906
rect 20242 5854 20254 5906
rect 20738 5854 20750 5906
rect 20802 5854 20814 5906
rect 24434 5854 24446 5906
rect 24498 5854 24510 5906
rect 28018 5854 28030 5906
rect 28082 5854 28094 5906
rect 28690 5854 28702 5906
rect 28754 5854 28766 5906
rect 29362 5854 29374 5906
rect 29426 5854 29438 5906
rect 33618 5854 33630 5906
rect 33682 5854 33694 5906
rect 35186 5854 35198 5906
rect 35250 5854 35262 5906
rect 38882 5854 38894 5906
rect 38946 5854 38958 5906
rect 42242 5854 42254 5906
rect 42306 5854 42318 5906
rect 17838 5842 17890 5854
rect 27246 5842 27298 5854
rect 34750 5842 34802 5854
rect 38670 5842 38722 5854
rect 40910 5842 40962 5854
rect 23998 5794 24050 5806
rect 16706 5742 16718 5794
rect 16770 5742 16782 5794
rect 19282 5742 19294 5794
rect 19346 5742 19358 5794
rect 27682 5742 27694 5794
rect 27746 5742 27758 5794
rect 37986 5742 37998 5794
rect 38050 5742 38062 5794
rect 42130 5742 42142 5794
rect 42194 5742 42206 5794
rect 23998 5730 24050 5742
rect 25342 5682 25394 5694
rect 38546 5630 38558 5682
rect 38610 5630 38622 5682
rect 25342 5618 25394 5630
rect 1344 5514 44576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 44576 5514
rect 1344 5428 44576 5462
rect 20862 5346 20914 5358
rect 12338 5294 12350 5346
rect 12402 5294 12414 5346
rect 14130 5294 14142 5346
rect 14194 5294 14206 5346
rect 20862 5282 20914 5294
rect 22430 5346 22482 5358
rect 29362 5294 29374 5346
rect 29426 5294 29438 5346
rect 22430 5282 22482 5294
rect 21646 5234 21698 5246
rect 12562 5182 12574 5234
rect 12626 5182 12638 5234
rect 14242 5182 14254 5234
rect 14306 5182 14318 5234
rect 28130 5182 28142 5234
rect 28194 5182 28206 5234
rect 29474 5182 29486 5234
rect 29538 5182 29550 5234
rect 31042 5182 31054 5234
rect 31106 5182 31118 5234
rect 33058 5182 33070 5234
rect 33122 5182 33134 5234
rect 40338 5182 40350 5234
rect 40402 5182 40414 5234
rect 41458 5182 41470 5234
rect 41522 5182 41534 5234
rect 21646 5170 21698 5182
rect 16382 5122 16434 5134
rect 12674 5070 12686 5122
rect 12738 5070 12750 5122
rect 14914 5070 14926 5122
rect 14978 5070 14990 5122
rect 15698 5070 15710 5122
rect 15762 5070 15774 5122
rect 16382 5058 16434 5070
rect 17390 5122 17442 5134
rect 22206 5122 22258 5134
rect 25902 5122 25954 5134
rect 17826 5070 17838 5122
rect 17890 5070 17902 5122
rect 25442 5070 25454 5122
rect 25506 5070 25518 5122
rect 17390 5058 17442 5070
rect 22206 5058 22258 5070
rect 25902 5058 25954 5070
rect 27470 5122 27522 5134
rect 30606 5122 30658 5134
rect 37102 5122 37154 5134
rect 42142 5122 42194 5134
rect 28354 5070 28366 5122
rect 28418 5070 28430 5122
rect 30034 5070 30046 5122
rect 30098 5070 30110 5122
rect 35970 5070 35982 5122
rect 36034 5070 36046 5122
rect 36418 5070 36430 5122
rect 36482 5070 36494 5122
rect 37538 5070 37550 5122
rect 37602 5070 37614 5122
rect 41234 5070 41246 5122
rect 41298 5070 41310 5122
rect 42690 5070 42702 5122
rect 42754 5070 42766 5122
rect 27470 5058 27522 5070
rect 30606 5058 30658 5070
rect 37102 5058 37154 5070
rect 42142 5058 42194 5070
rect 16606 5010 16658 5022
rect 16606 4946 16658 4958
rect 42478 4898 42530 4910
rect 20290 4846 20302 4898
rect 20354 4846 20366 4898
rect 23202 4846 23214 4898
rect 23266 4846 23278 4898
rect 33618 4846 33630 4898
rect 33682 4846 33694 4898
rect 39778 4846 39790 4898
rect 39842 4846 39854 4898
rect 42478 4834 42530 4846
rect 1344 4730 44576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 44576 4730
rect 1344 4644 44576 4678
rect 16494 4562 16546 4574
rect 14802 4510 14814 4562
rect 14866 4510 14878 4562
rect 16494 4498 16546 4510
rect 17950 4562 18002 4574
rect 17950 4498 18002 4510
rect 25230 4562 25282 4574
rect 37774 4562 37826 4574
rect 37202 4510 37214 4562
rect 37266 4510 37278 4562
rect 25230 4498 25282 4510
rect 37774 4498 37826 4510
rect 39790 4562 39842 4574
rect 39790 4498 39842 4510
rect 41582 4562 41634 4574
rect 41582 4498 41634 4510
rect 19070 4450 19122 4462
rect 19070 4386 19122 4398
rect 39454 4450 39506 4462
rect 39454 4386 39506 4398
rect 41694 4450 41746 4462
rect 41694 4386 41746 4398
rect 12126 4338 12178 4350
rect 17390 4338 17442 4350
rect 24670 4338 24722 4350
rect 34302 4338 34354 4350
rect 37998 4338 38050 4350
rect 12450 4286 12462 4338
rect 12514 4286 12526 4338
rect 16706 4286 16718 4338
rect 16770 4286 16782 4338
rect 19506 4286 19518 4338
rect 19570 4286 19582 4338
rect 21522 4286 21534 4338
rect 21586 4286 21598 4338
rect 22306 4286 22318 4338
rect 22370 4286 22382 4338
rect 23762 4286 23774 4338
rect 23826 4286 23838 4338
rect 25442 4286 25454 4338
rect 25506 4286 25518 4338
rect 28578 4286 28590 4338
rect 28642 4286 28654 4338
rect 30818 4286 30830 4338
rect 30882 4286 30894 4338
rect 34738 4286 34750 4338
rect 34802 4286 34814 4338
rect 38658 4286 38670 4338
rect 38722 4286 38734 4338
rect 12126 4274 12178 4286
rect 17390 4274 17442 4286
rect 24670 4274 24722 4286
rect 34302 4274 34354 4286
rect 37998 4274 38050 4286
rect 29486 4226 29538 4238
rect 15362 4174 15374 4226
rect 15426 4174 15438 4226
rect 19842 4174 19854 4226
rect 19906 4174 19918 4226
rect 21410 4174 21422 4226
rect 21474 4174 21486 4226
rect 22978 4174 22990 4226
rect 23042 4174 23054 4226
rect 24322 4174 24334 4226
rect 24386 4174 24398 4226
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 29486 4162 29538 4174
rect 29934 4226 29986 4238
rect 41022 4226 41074 4238
rect 30482 4174 30494 4226
rect 30546 4174 30558 4226
rect 38434 4174 38446 4226
rect 38498 4174 38510 4226
rect 29934 4162 29986 4174
rect 41022 4162 41074 4174
rect 44270 4226 44322 4238
rect 44270 4162 44322 4174
rect 21186 4062 21198 4114
rect 21250 4062 21262 4114
rect 23090 4062 23102 4114
rect 23154 4062 23166 4114
rect 28690 4062 28702 4114
rect 28754 4062 28766 4114
rect 1344 3946 44576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 44576 3946
rect 1344 3860 44576 3894
rect 35086 3778 35138 3790
rect 14466 3726 14478 3778
rect 14530 3726 14542 3778
rect 35086 3714 35138 3726
rect 35198 3666 35250 3678
rect 14242 3614 14254 3666
rect 14306 3614 14318 3666
rect 35198 3602 35250 3614
rect 37886 3554 37938 3566
rect 14018 3502 14030 3554
rect 14082 3502 14094 3554
rect 21298 3502 21310 3554
rect 21362 3502 21374 3554
rect 23090 3502 23102 3554
rect 23154 3502 23166 3554
rect 37886 3490 37938 3502
rect 38558 3554 38610 3566
rect 38558 3490 38610 3502
rect 21086 3442 21138 3454
rect 21086 3378 21138 3390
rect 22878 3442 22930 3454
rect 22878 3378 22930 3390
rect 37550 3442 37602 3454
rect 37550 3378 37602 3390
rect 38222 3442 38274 3454
rect 38222 3378 38274 3390
rect 43822 3442 43874 3454
rect 43822 3378 43874 3390
rect 44158 3442 44210 3454
rect 44158 3378 44210 3390
rect 1344 3162 44576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 44576 3162
rect 1344 3076 44576 3110
<< via1 >>
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 32846 42030 32898 42082
rect 34078 42030 34130 42082
rect 43598 42030 43650 42082
rect 43710 42030 43762 42082
rect 33070 41918 33122 41970
rect 33854 41918 33906 41970
rect 34190 41918 34242 41970
rect 43038 41918 43090 41970
rect 32510 41806 32562 41858
rect 41918 41806 41970 41858
rect 43710 41694 43762 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 34638 41246 34690 41298
rect 40910 41246 40962 41298
rect 44158 41246 44210 41298
rect 29934 41134 29986 41186
rect 30158 41134 30210 41186
rect 31838 41134 31890 41186
rect 35534 41134 35586 41186
rect 38110 41134 38162 41186
rect 41246 41134 41298 41186
rect 32510 41022 32562 41074
rect 36094 41022 36146 41074
rect 38782 41022 38834 41074
rect 42030 41022 42082 41074
rect 29598 40910 29650 40962
rect 34862 40910 34914 40962
rect 34974 40910 35026 40962
rect 35198 40910 35250 40962
rect 35870 40910 35922 40962
rect 35982 40910 36034 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 32510 40574 32562 40626
rect 38222 40574 38274 40626
rect 39118 40574 39170 40626
rect 39342 40574 39394 40626
rect 31838 40462 31890 40514
rect 33966 40462 34018 40514
rect 36542 40462 36594 40514
rect 39566 40462 39618 40514
rect 39678 40462 39730 40514
rect 40238 40462 40290 40514
rect 40350 40462 40402 40514
rect 26910 40350 26962 40402
rect 30046 40350 30098 40402
rect 30270 40350 30322 40402
rect 30718 40350 30770 40402
rect 31614 40350 31666 40402
rect 32174 40350 32226 40402
rect 33070 40350 33122 40402
rect 33518 40350 33570 40402
rect 33742 40350 33794 40402
rect 37326 40350 37378 40402
rect 39006 40350 39058 40402
rect 39902 40350 39954 40402
rect 40910 40350 40962 40402
rect 27582 40238 27634 40290
rect 29710 40238 29762 40290
rect 30158 40238 30210 40290
rect 34078 40238 34130 40290
rect 34414 40238 34466 40290
rect 38110 40238 38162 40290
rect 38670 40238 38722 40290
rect 41694 40238 41746 40290
rect 43822 40238 43874 40290
rect 38558 40126 38610 40178
rect 40238 40126 40290 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 27694 39790 27746 39842
rect 37102 39790 37154 39842
rect 26798 39678 26850 39730
rect 27582 39678 27634 39730
rect 28590 39678 28642 39730
rect 29934 39678 29986 39730
rect 32062 39678 32114 39730
rect 35310 39678 35362 39730
rect 36094 39678 36146 39730
rect 38334 39678 38386 39730
rect 40462 39678 40514 39730
rect 41134 39678 41186 39730
rect 26686 39566 26738 39618
rect 28366 39566 28418 39618
rect 29262 39566 29314 39618
rect 32510 39566 32562 39618
rect 35646 39566 35698 39618
rect 36990 39566 37042 39618
rect 37550 39566 37602 39618
rect 43934 39566 43986 39618
rect 27022 39454 27074 39506
rect 33182 39454 33234 39506
rect 35870 39454 35922 39506
rect 36206 39454 36258 39506
rect 43262 39454 43314 39506
rect 27470 39342 27522 39394
rect 28030 39342 28082 39394
rect 37102 39342 37154 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 30382 39006 30434 39058
rect 30830 39006 30882 39058
rect 31950 39006 32002 39058
rect 36318 39006 36370 39058
rect 38670 39006 38722 39058
rect 39790 39006 39842 39058
rect 41246 39006 41298 39058
rect 43150 39006 43202 39058
rect 30494 38894 30546 38946
rect 31278 38894 31330 38946
rect 31502 38894 31554 38946
rect 36430 38894 36482 38946
rect 38222 38894 38274 38946
rect 38782 38894 38834 38946
rect 39678 38894 39730 38946
rect 27246 38782 27298 38834
rect 30606 38782 30658 38834
rect 32510 38782 32562 38834
rect 33070 38782 33122 38834
rect 37886 38782 37938 38834
rect 38558 38782 38610 38834
rect 39230 38782 39282 38834
rect 40014 38782 40066 38834
rect 41022 38782 41074 38834
rect 44158 38782 44210 38834
rect 27918 38670 27970 38722
rect 30046 38670 30098 38722
rect 31614 38670 31666 38722
rect 32286 38670 32338 38722
rect 33854 38670 33906 38722
rect 35982 38670 36034 38722
rect 39678 38670 39730 38722
rect 37998 38558 38050 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 43150 38222 43202 38274
rect 29262 38110 29314 38162
rect 30158 38110 30210 38162
rect 33182 38110 33234 38162
rect 34414 38110 34466 38162
rect 29038 37998 29090 38050
rect 29486 37998 29538 38050
rect 29710 37998 29762 38050
rect 30046 37998 30098 38050
rect 30718 37998 30770 38050
rect 33294 37998 33346 38050
rect 34078 37998 34130 38050
rect 35086 37998 35138 38050
rect 37214 37998 37266 38050
rect 40126 37998 40178 38050
rect 40574 37998 40626 38050
rect 40910 37998 40962 38050
rect 41246 37998 41298 38050
rect 41582 37998 41634 38050
rect 43598 37998 43650 38050
rect 43934 37998 43986 38050
rect 30270 37886 30322 37938
rect 33630 37886 33682 37938
rect 35422 37886 35474 37938
rect 36990 37886 37042 37938
rect 40462 37886 40514 37938
rect 40798 37886 40850 37938
rect 41358 37886 41410 37938
rect 41806 37886 41858 37938
rect 42478 37886 42530 37938
rect 43038 37886 43090 37938
rect 43150 37886 43202 37938
rect 43710 37886 43762 37938
rect 31838 37774 31890 37826
rect 33070 37774 33122 37826
rect 40238 37774 40290 37826
rect 42142 37774 42194 37826
rect 42590 37774 42642 37826
rect 42814 37774 42866 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 29934 37438 29986 37490
rect 33742 37438 33794 37490
rect 39118 37438 39170 37490
rect 26238 37326 26290 37378
rect 27806 37326 27858 37378
rect 29822 37326 29874 37378
rect 33630 37326 33682 37378
rect 36990 37326 37042 37378
rect 38446 37326 38498 37378
rect 38782 37326 38834 37378
rect 41134 37326 41186 37378
rect 26126 37214 26178 37266
rect 26910 37214 26962 37266
rect 27246 37214 27298 37266
rect 28030 37214 28082 37266
rect 30158 37214 30210 37266
rect 33966 37214 34018 37266
rect 36766 37214 36818 37266
rect 37662 37214 37714 37266
rect 38222 37214 38274 37266
rect 39454 37214 39506 37266
rect 41022 37214 41074 37266
rect 41358 37214 41410 37266
rect 41582 37214 41634 37266
rect 25230 37102 25282 37154
rect 38334 37102 38386 37154
rect 39566 37102 39618 37154
rect 25342 36990 25394 37042
rect 27134 36990 27186 37042
rect 37214 36990 37266 37042
rect 37550 36990 37602 37042
rect 37998 36990 38050 37042
rect 43486 36990 43538 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 7310 36542 7362 36594
rect 34862 36542 34914 36594
rect 38670 36542 38722 36594
rect 40798 36542 40850 36594
rect 41134 36542 41186 36594
rect 10110 36430 10162 36482
rect 15598 36430 15650 36482
rect 16046 36430 16098 36482
rect 25902 36430 25954 36482
rect 26462 36430 26514 36482
rect 27134 36430 27186 36482
rect 31950 36430 32002 36482
rect 37886 36430 37938 36482
rect 43934 36430 43986 36482
rect 9438 36318 9490 36370
rect 26910 36318 26962 36370
rect 27470 36318 27522 36370
rect 28030 36318 28082 36370
rect 32734 36318 32786 36370
rect 43262 36318 43314 36370
rect 18286 36206 18338 36258
rect 19070 36206 19122 36258
rect 19406 36206 19458 36258
rect 23550 36206 23602 36258
rect 27246 36206 27298 36258
rect 27358 36206 27410 36258
rect 27918 36206 27970 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 10446 35870 10498 35922
rect 17726 35870 17778 35922
rect 35982 35870 36034 35922
rect 39342 35870 39394 35922
rect 40014 35870 40066 35922
rect 15822 35758 15874 35810
rect 16158 35758 16210 35810
rect 16494 35758 16546 35810
rect 17502 35758 17554 35810
rect 18286 35758 18338 35810
rect 18622 35758 18674 35810
rect 19294 35758 19346 35810
rect 23550 35758 23602 35810
rect 31838 35758 31890 35810
rect 35534 35758 35586 35810
rect 36766 35758 36818 35810
rect 43038 35758 43090 35810
rect 10782 35646 10834 35698
rect 16718 35646 16770 35698
rect 17390 35646 17442 35698
rect 17950 35646 18002 35698
rect 18846 35646 18898 35698
rect 19518 35646 19570 35698
rect 20302 35646 20354 35698
rect 24110 35646 24162 35698
rect 24222 35646 24274 35698
rect 24446 35646 24498 35698
rect 24670 35646 24722 35698
rect 25454 35646 25506 35698
rect 26014 35646 26066 35698
rect 29038 35646 29090 35698
rect 29374 35646 29426 35698
rect 29598 35646 29650 35698
rect 32174 35646 32226 35698
rect 32958 35646 33010 35698
rect 33406 35646 33458 35698
rect 33630 35646 33682 35698
rect 35758 35646 35810 35698
rect 36318 35646 36370 35698
rect 37438 35646 37490 35698
rect 37662 35646 37714 35698
rect 38782 35646 38834 35698
rect 39006 35646 39058 35698
rect 39566 35646 39618 35698
rect 40238 35646 40290 35698
rect 43822 35646 43874 35698
rect 20974 35534 21026 35586
rect 23102 35534 23154 35586
rect 24334 35534 24386 35586
rect 28366 35534 28418 35586
rect 28702 35534 28754 35586
rect 28814 35534 28866 35586
rect 33182 35534 33234 35586
rect 35422 35534 35474 35586
rect 40910 35534 40962 35586
rect 23438 35422 23490 35474
rect 29710 35422 29762 35474
rect 36430 35422 36482 35474
rect 37102 35422 37154 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 29374 35086 29426 35138
rect 38334 35086 38386 35138
rect 39790 35086 39842 35138
rect 9326 34974 9378 35026
rect 11454 34974 11506 35026
rect 24894 34974 24946 35026
rect 26126 34974 26178 35026
rect 27358 34974 27410 35026
rect 31054 34974 31106 35026
rect 32286 34974 32338 35026
rect 34414 34974 34466 35026
rect 41918 34974 41970 35026
rect 44046 34974 44098 35026
rect 8654 34862 8706 34914
rect 16158 34862 16210 34914
rect 16830 34862 16882 34914
rect 18958 34862 19010 34914
rect 21982 34862 22034 34914
rect 22542 34862 22594 34914
rect 25230 34862 25282 34914
rect 27022 34862 27074 34914
rect 27470 34862 27522 34914
rect 29150 34862 29202 34914
rect 29598 34862 29650 34914
rect 31614 34862 31666 34914
rect 35310 34862 35362 34914
rect 35422 34862 35474 34914
rect 35534 34862 35586 34914
rect 36094 34862 36146 34914
rect 36206 34862 36258 34914
rect 38334 34862 38386 34914
rect 40014 34862 40066 34914
rect 40798 34862 40850 34914
rect 41246 34862 41298 34914
rect 15822 34750 15874 34802
rect 15934 34750 15986 34802
rect 20414 34750 20466 34802
rect 20526 34750 20578 34802
rect 25342 34750 25394 34802
rect 26462 34750 26514 34802
rect 28142 34750 28194 34802
rect 29934 34750 29986 34802
rect 31166 34750 31218 34802
rect 35870 34750 35922 34802
rect 36990 34750 37042 34802
rect 37662 34750 37714 34802
rect 38670 34750 38722 34802
rect 40462 34750 40514 34802
rect 15598 34638 15650 34690
rect 19966 34638 20018 34690
rect 20190 34638 20242 34690
rect 25566 34638 25618 34690
rect 25902 34638 25954 34690
rect 26014 34638 26066 34690
rect 26238 34638 26290 34690
rect 29486 34638 29538 34690
rect 30942 34638 30994 34690
rect 37326 34638 37378 34690
rect 37998 34638 38050 34690
rect 39454 34638 39506 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 16270 34302 16322 34354
rect 20190 34302 20242 34354
rect 20974 34302 21026 34354
rect 24558 34302 24610 34354
rect 26462 34302 26514 34354
rect 30942 34302 30994 34354
rect 39678 34302 39730 34354
rect 40350 34302 40402 34354
rect 41806 34302 41858 34354
rect 43262 34302 43314 34354
rect 43486 34302 43538 34354
rect 8206 34190 8258 34242
rect 8654 34190 8706 34242
rect 11230 34190 11282 34242
rect 24446 34190 24498 34242
rect 25790 34190 25842 34242
rect 27358 34190 27410 34242
rect 30382 34190 30434 34242
rect 31054 34190 31106 34242
rect 32286 34190 32338 34242
rect 32510 34190 32562 34242
rect 36654 34190 36706 34242
rect 36990 34190 37042 34242
rect 37774 34190 37826 34242
rect 39342 34190 39394 34242
rect 40014 34190 40066 34242
rect 40910 34190 40962 34242
rect 41246 34190 41298 34242
rect 42590 34190 42642 34242
rect 43150 34190 43202 34242
rect 7982 34078 8034 34130
rect 8990 34078 9042 34130
rect 9886 34078 9938 34130
rect 10558 34078 10610 34130
rect 11454 34078 11506 34130
rect 12686 34078 12738 34130
rect 13134 34078 13186 34130
rect 15374 34078 15426 34130
rect 17278 34078 17330 34130
rect 17950 34078 18002 34130
rect 21198 34078 21250 34130
rect 21982 34078 22034 34130
rect 24782 34078 24834 34130
rect 25678 34078 25730 34130
rect 26238 34078 26290 34130
rect 28254 34078 28306 34130
rect 28926 34078 28978 34130
rect 29486 34078 29538 34130
rect 30606 34078 30658 34130
rect 31278 34078 31330 34130
rect 31950 34078 32002 34130
rect 33070 34078 33122 34130
rect 36430 34078 36482 34130
rect 36542 34078 36594 34130
rect 37214 34078 37266 34130
rect 42142 34078 42194 34130
rect 10334 33966 10386 34018
rect 24110 33966 24162 34018
rect 25454 33966 25506 34018
rect 26798 33966 26850 34018
rect 29934 33966 29986 34018
rect 32062 33966 32114 34018
rect 33854 33966 33906 34018
rect 35982 33966 36034 34018
rect 42478 33966 42530 34018
rect 43822 33966 43874 34018
rect 37326 33854 37378 33906
rect 37662 33854 37714 33906
rect 42814 33854 42866 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 14590 33518 14642 33570
rect 35422 33518 35474 33570
rect 41022 33518 41074 33570
rect 8430 33406 8482 33458
rect 10558 33406 10610 33458
rect 22094 33406 22146 33458
rect 24222 33406 24274 33458
rect 27358 33406 27410 33458
rect 34526 33406 34578 33458
rect 7758 33294 7810 33346
rect 15598 33294 15650 33346
rect 17726 33294 17778 33346
rect 18174 33294 18226 33346
rect 18622 33294 18674 33346
rect 18958 33294 19010 33346
rect 21310 33294 21362 33346
rect 25790 33294 25842 33346
rect 27022 33294 27074 33346
rect 29262 33294 29314 33346
rect 29710 33294 29762 33346
rect 31614 33294 31666 33346
rect 35534 33294 35586 33346
rect 36094 33294 36146 33346
rect 36430 33294 36482 33346
rect 37102 33294 37154 33346
rect 38446 33294 38498 33346
rect 39902 33294 39954 33346
rect 40238 33294 40290 33346
rect 44046 33294 44098 33346
rect 6974 33182 7026 33234
rect 7310 33182 7362 33234
rect 18734 33182 18786 33234
rect 25902 33182 25954 33234
rect 26910 33182 26962 33234
rect 30158 33182 30210 33234
rect 32398 33182 32450 33234
rect 35870 33182 35922 33234
rect 37662 33182 37714 33234
rect 37998 33182 38050 33234
rect 38670 33182 38722 33234
rect 38782 33182 38834 33234
rect 40462 33182 40514 33234
rect 40574 33182 40626 33234
rect 24670 33070 24722 33122
rect 25006 33070 25058 33122
rect 36206 33070 36258 33122
rect 37326 33070 37378 33122
rect 39566 33070 39618 33122
rect 43150 33070 43202 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 14030 32734 14082 32786
rect 14702 32734 14754 32786
rect 15934 32734 15986 32786
rect 17950 32734 18002 32786
rect 24670 32734 24722 32786
rect 25790 32734 25842 32786
rect 26126 32734 26178 32786
rect 27694 32734 27746 32786
rect 28030 32734 28082 32786
rect 28926 32734 28978 32786
rect 29598 32734 29650 32786
rect 32398 32734 32450 32786
rect 36878 32734 36930 32786
rect 37662 32734 37714 32786
rect 37998 32734 38050 32786
rect 39678 32734 39730 32786
rect 40350 32734 40402 32786
rect 42926 32734 42978 32786
rect 8206 32622 8258 32674
rect 9550 32622 9602 32674
rect 14926 32622 14978 32674
rect 15598 32622 15650 32674
rect 16158 32622 16210 32674
rect 24334 32622 24386 32674
rect 26350 32622 26402 32674
rect 26910 32622 26962 32674
rect 28478 32622 28530 32674
rect 29038 32622 29090 32674
rect 29374 32622 29426 32674
rect 32510 32622 32562 32674
rect 33854 32622 33906 32674
rect 35982 32622 36034 32674
rect 36206 32622 36258 32674
rect 36430 32622 36482 32674
rect 36766 32622 36818 32674
rect 38782 32622 38834 32674
rect 38894 32622 38946 32674
rect 40014 32622 40066 32674
rect 43374 32622 43426 32674
rect 8878 32510 8930 32562
rect 9998 32510 10050 32562
rect 10446 32510 10498 32562
rect 10894 32510 10946 32562
rect 11566 32510 11618 32562
rect 14590 32510 14642 32562
rect 15038 32510 15090 32562
rect 15486 32510 15538 32562
rect 15822 32510 15874 32562
rect 16270 32510 16322 32562
rect 18286 32510 18338 32562
rect 20190 32510 20242 32562
rect 25902 32510 25954 32562
rect 26686 32510 26738 32562
rect 27022 32510 27074 32562
rect 27246 32510 27298 32562
rect 28814 32510 28866 32562
rect 32174 32510 32226 32562
rect 33182 32510 33234 32562
rect 33518 32510 33570 32562
rect 35198 32510 35250 32562
rect 35646 32510 35698 32562
rect 36318 32510 36370 32562
rect 37102 32510 37154 32562
rect 37438 32510 37490 32562
rect 39118 32510 39170 32562
rect 39342 32510 39394 32562
rect 41022 32510 41074 32562
rect 41358 32510 41410 32562
rect 41806 32510 41858 32562
rect 42030 32510 42082 32562
rect 42478 32510 42530 32562
rect 43598 32510 43650 32562
rect 6078 32398 6130 32450
rect 20862 32398 20914 32450
rect 22990 32398 23042 32450
rect 26014 32398 26066 32450
rect 27918 32398 27970 32450
rect 33406 32398 33458 32450
rect 34974 32398 35026 32450
rect 42254 32398 42306 32450
rect 29710 32286 29762 32338
rect 34638 32286 34690 32338
rect 35534 32286 35586 32338
rect 41134 32286 41186 32338
rect 41470 32286 41522 32338
rect 42702 32286 42754 32338
rect 43038 32286 43090 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 26910 31950 26962 32002
rect 31838 31950 31890 32002
rect 39678 31950 39730 32002
rect 7982 31838 8034 31890
rect 10110 31838 10162 31890
rect 17166 31838 17218 31890
rect 31054 31838 31106 31890
rect 33518 31838 33570 31890
rect 35646 31838 35698 31890
rect 37774 31838 37826 31890
rect 7198 31726 7250 31778
rect 11454 31726 11506 31778
rect 13470 31726 13522 31778
rect 14030 31726 14082 31778
rect 16158 31726 16210 31778
rect 23438 31726 23490 31778
rect 23886 31726 23938 31778
rect 27358 31726 27410 31778
rect 28030 31726 28082 31778
rect 31278 31726 31330 31778
rect 32734 31726 32786 31778
rect 39118 31726 39170 31778
rect 39342 31726 39394 31778
rect 40350 31726 40402 31778
rect 44046 31726 44098 31778
rect 17502 31614 17554 31666
rect 27806 31614 27858 31666
rect 37326 31614 37378 31666
rect 37438 31614 37490 31666
rect 38670 31614 38722 31666
rect 38782 31614 38834 31666
rect 40014 31614 40066 31666
rect 40574 31614 40626 31666
rect 41246 31614 41298 31666
rect 11118 31502 11170 31554
rect 17838 31502 17890 31554
rect 18286 31502 18338 31554
rect 26350 31502 26402 31554
rect 27134 31502 27186 31554
rect 32398 31502 32450 31554
rect 36990 31502 37042 31554
rect 37214 31502 37266 31554
rect 38446 31502 38498 31554
rect 40238 31502 40290 31554
rect 41022 31502 41074 31554
rect 41134 31502 41186 31554
rect 43150 31502 43202 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 13918 31166 13970 31218
rect 14478 31166 14530 31218
rect 14814 31166 14866 31218
rect 16382 31166 16434 31218
rect 20078 31166 20130 31218
rect 24222 31166 24274 31218
rect 27022 31166 27074 31218
rect 27918 31166 27970 31218
rect 31726 31166 31778 31218
rect 38894 31166 38946 31218
rect 40350 31166 40402 31218
rect 8318 31054 8370 31106
rect 14926 31054 14978 31106
rect 20526 31054 20578 31106
rect 25678 31054 25730 31106
rect 26014 31054 26066 31106
rect 26686 31054 26738 31106
rect 30270 31054 30322 31106
rect 30942 31054 30994 31106
rect 33070 31054 33122 31106
rect 35086 31054 35138 31106
rect 35422 31054 35474 31106
rect 39118 31054 39170 31106
rect 39678 31054 39730 31106
rect 39902 31054 39954 31106
rect 43038 31054 43090 31106
rect 8654 30942 8706 30994
rect 9550 30942 9602 30994
rect 9998 30942 10050 30994
rect 10782 30942 10834 30994
rect 11454 30942 11506 30994
rect 14590 30942 14642 30994
rect 16718 30942 16770 30994
rect 19854 30942 19906 30994
rect 24558 30942 24610 30994
rect 30606 30942 30658 30994
rect 31278 30942 31330 30994
rect 31726 30942 31778 30994
rect 32510 30942 32562 30994
rect 33294 30942 33346 30994
rect 35758 30942 35810 30994
rect 39230 30942 39282 30994
rect 39790 30942 39842 30994
rect 43710 30942 43762 30994
rect 10334 30830 10386 30882
rect 20974 30830 21026 30882
rect 21422 30830 21474 30882
rect 27582 30830 27634 30882
rect 36542 30830 36594 30882
rect 38670 30830 38722 30882
rect 40910 30830 40962 30882
rect 20414 30718 20466 30770
rect 21310 30718 21362 30770
rect 27246 30718 27298 30770
rect 28030 30718 28082 30770
rect 31502 30718 31554 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 27022 30382 27074 30434
rect 33742 30382 33794 30434
rect 17054 30270 17106 30322
rect 20750 30270 20802 30322
rect 30494 30270 30546 30322
rect 31950 30270 32002 30322
rect 33406 30270 33458 30322
rect 39342 30270 39394 30322
rect 13806 30158 13858 30210
rect 14254 30158 14306 30210
rect 17838 30158 17890 30210
rect 18622 30158 18674 30210
rect 23550 30158 23602 30210
rect 23998 30158 24050 30210
rect 27470 30158 27522 30210
rect 30606 30158 30658 30210
rect 32286 30158 32338 30210
rect 32958 30158 33010 30210
rect 34302 30158 34354 30210
rect 36990 30158 37042 30210
rect 37214 30158 37266 30210
rect 37550 30158 37602 30210
rect 37998 30158 38050 30210
rect 41470 30158 41522 30210
rect 42142 30158 42194 30210
rect 42590 30158 42642 30210
rect 42814 30158 42866 30210
rect 43486 30158 43538 30210
rect 21646 30046 21698 30098
rect 28142 30046 28194 30098
rect 29598 30046 29650 30098
rect 29934 30046 29986 30098
rect 31278 30046 31330 30098
rect 34078 30046 34130 30098
rect 35086 30046 35138 30098
rect 37102 30046 37154 30098
rect 38222 30046 38274 30098
rect 16494 29934 16546 29986
rect 21310 29934 21362 29986
rect 26462 29934 26514 29986
rect 27246 29934 27298 29986
rect 27806 29934 27858 29986
rect 28030 29934 28082 29986
rect 32734 29934 32786 29986
rect 33630 29934 33682 29986
rect 34750 29934 34802 29986
rect 38782 29934 38834 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 13246 29598 13298 29650
rect 15038 29598 15090 29650
rect 16382 29598 16434 29650
rect 24334 29598 24386 29650
rect 25342 29598 25394 29650
rect 29934 29598 29986 29650
rect 30606 29598 30658 29650
rect 34190 29598 34242 29650
rect 8206 29486 8258 29538
rect 15150 29486 15202 29538
rect 16270 29486 16322 29538
rect 17502 29486 17554 29538
rect 18286 29486 18338 29538
rect 20638 29486 20690 29538
rect 23662 29486 23714 29538
rect 26238 29486 26290 29538
rect 27582 29486 27634 29538
rect 27918 29486 27970 29538
rect 28702 29486 28754 29538
rect 32510 29486 32562 29538
rect 33070 29486 33122 29538
rect 35422 29486 35474 29538
rect 40014 29486 40066 29538
rect 41694 29486 41746 29538
rect 8878 29374 8930 29426
rect 9550 29374 9602 29426
rect 10110 29374 10162 29426
rect 12238 29374 12290 29426
rect 17838 29374 17890 29426
rect 19854 29374 19906 29426
rect 23998 29374 24050 29426
rect 24670 29374 24722 29426
rect 25678 29374 25730 29426
rect 26462 29374 26514 29426
rect 27022 29374 27074 29426
rect 27358 29374 27410 29426
rect 28814 29374 28866 29426
rect 29262 29374 29314 29426
rect 29710 29374 29762 29426
rect 30270 29374 30322 29426
rect 30494 29374 30546 29426
rect 30718 29374 30770 29426
rect 30830 29374 30882 29426
rect 31950 29374 32002 29426
rect 33406 29374 33458 29426
rect 34750 29374 34802 29426
rect 40238 29374 40290 29426
rect 40910 29374 40962 29426
rect 6078 29262 6130 29314
rect 13918 29262 13970 29314
rect 16830 29262 16882 29314
rect 22766 29262 22818 29314
rect 33182 29262 33234 29314
rect 33966 29262 34018 29314
rect 34302 29262 34354 29314
rect 37550 29262 37602 29314
rect 43822 29262 43874 29314
rect 14030 29150 14082 29202
rect 16718 29150 16770 29202
rect 18398 29150 18450 29202
rect 28702 29150 28754 29202
rect 32398 29150 32450 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 30718 28814 30770 28866
rect 8318 28702 8370 28754
rect 10446 28702 10498 28754
rect 19182 28702 19234 28754
rect 30942 28702 30994 28754
rect 33070 28702 33122 28754
rect 41918 28702 41970 28754
rect 44046 28702 44098 28754
rect 7646 28590 7698 28642
rect 15934 28590 15986 28642
rect 16382 28590 16434 28642
rect 20638 28590 20690 28642
rect 24782 28590 24834 28642
rect 25006 28590 25058 28642
rect 25566 28590 25618 28642
rect 28702 28590 28754 28642
rect 29710 28590 29762 28642
rect 30270 28590 30322 28642
rect 33742 28590 33794 28642
rect 34302 28590 34354 28642
rect 41246 28590 41298 28642
rect 18622 28478 18674 28530
rect 29822 28478 29874 28530
rect 30158 28478 30210 28530
rect 20302 28366 20354 28418
rect 24446 28366 24498 28418
rect 28030 28366 28082 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 13022 28030 13074 28082
rect 24670 28030 24722 28082
rect 26014 28030 26066 28082
rect 28030 28030 28082 28082
rect 28254 28030 28306 28082
rect 13806 27918 13858 27970
rect 17390 27918 17442 27970
rect 17502 27918 17554 27970
rect 18174 27918 18226 27970
rect 21422 27918 21474 27970
rect 25230 27918 25282 27970
rect 25902 27918 25954 27970
rect 27470 27918 27522 27970
rect 28366 27918 28418 27970
rect 29150 27918 29202 27970
rect 43822 27918 43874 27970
rect 11006 27806 11058 27858
rect 16046 27806 16098 27858
rect 16606 27806 16658 27858
rect 18734 27806 18786 27858
rect 19182 27806 19234 27858
rect 24446 27806 24498 27858
rect 25566 27806 25618 27858
rect 26574 27806 26626 27858
rect 26910 27806 26962 27858
rect 27358 27806 27410 27858
rect 29598 27806 29650 27858
rect 44158 27806 44210 27858
rect 11118 27694 11170 27746
rect 11566 27694 11618 27746
rect 12014 27694 12066 27746
rect 21982 27694 22034 27746
rect 23998 27694 24050 27746
rect 29262 27694 29314 27746
rect 30382 27694 30434 27746
rect 32510 27694 32562 27746
rect 43150 27694 43202 27746
rect 43598 27694 43650 27746
rect 11902 27582 11954 27634
rect 18286 27582 18338 27634
rect 26014 27582 26066 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 15822 27246 15874 27298
rect 20190 27246 20242 27298
rect 21422 27246 21474 27298
rect 27806 27246 27858 27298
rect 9214 27134 9266 27186
rect 19630 27134 19682 27186
rect 20302 27134 20354 27186
rect 29598 27134 29650 27186
rect 35086 27134 35138 27186
rect 37102 27134 37154 27186
rect 44158 27134 44210 27186
rect 9662 27022 9714 27074
rect 10110 27022 10162 27074
rect 11006 27022 11058 27074
rect 11230 27022 11282 27074
rect 12462 27022 12514 27074
rect 16270 27022 16322 27074
rect 16606 27022 16658 27074
rect 24334 27022 24386 27074
rect 24782 27022 24834 27074
rect 32398 27022 32450 27074
rect 41022 27022 41074 27074
rect 41806 27022 41858 27074
rect 10558 26910 10610 26962
rect 11902 26910 11954 26962
rect 12238 26910 12290 26962
rect 15374 26910 15426 26962
rect 15710 26910 15762 26962
rect 18958 26910 19010 26962
rect 21310 26910 21362 26962
rect 27022 26910 27074 26962
rect 31726 26910 31778 26962
rect 34750 26910 34802 26962
rect 35646 26910 35698 26962
rect 36094 26910 36146 26962
rect 38558 26910 38610 26962
rect 39230 26910 39282 26962
rect 40798 26910 40850 26962
rect 35982 26798 36034 26850
rect 38222 26798 38274 26850
rect 38894 26798 38946 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 13134 26462 13186 26514
rect 13918 26462 13970 26514
rect 19070 26462 19122 26514
rect 25902 26462 25954 26514
rect 30942 26462 30994 26514
rect 34190 26462 34242 26514
rect 37550 26462 37602 26514
rect 44158 26462 44210 26514
rect 23550 26350 23602 26402
rect 26574 26350 26626 26402
rect 27022 26350 27074 26402
rect 30830 26350 30882 26402
rect 8542 26238 8594 26290
rect 8990 26238 9042 26290
rect 10110 26238 10162 26290
rect 10670 26238 10722 26290
rect 14142 26238 14194 26290
rect 16830 26238 16882 26290
rect 19294 26238 19346 26290
rect 20862 26238 20914 26290
rect 21310 26238 21362 26290
rect 26238 26238 26290 26290
rect 34638 26238 34690 26290
rect 34974 26238 35026 26290
rect 39454 26238 39506 26290
rect 41022 26238 41074 26290
rect 41806 26238 41858 26290
rect 9662 26126 9714 26178
rect 13470 26126 13522 26178
rect 17502 26126 17554 26178
rect 19854 26126 19906 26178
rect 20302 26126 20354 26178
rect 24110 26126 24162 26178
rect 27582 26126 27634 26178
rect 34078 26126 34130 26178
rect 37886 26126 37938 26178
rect 38894 26126 38946 26178
rect 9774 26014 9826 26066
rect 17390 26014 17442 26066
rect 19742 26014 19794 26066
rect 39230 26014 39282 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 19742 25678 19794 25730
rect 22542 25678 22594 25730
rect 23998 25678 24050 25730
rect 37550 25678 37602 25730
rect 38670 25678 38722 25730
rect 8318 25566 8370 25618
rect 9550 25566 9602 25618
rect 21422 25566 21474 25618
rect 22430 25566 22482 25618
rect 24110 25566 24162 25618
rect 28030 25566 28082 25618
rect 37886 25566 37938 25618
rect 41470 25566 41522 25618
rect 7310 25454 7362 25506
rect 7870 25454 7922 25506
rect 12350 25454 12402 25506
rect 12798 25454 12850 25506
rect 16158 25454 16210 25506
rect 16718 25454 16770 25506
rect 25678 25454 25730 25506
rect 26350 25454 26402 25506
rect 33070 25454 33122 25506
rect 33518 25454 33570 25506
rect 37438 25454 37490 25506
rect 38782 25454 38834 25506
rect 39454 25454 39506 25506
rect 10110 25342 10162 25394
rect 15710 25342 15762 25394
rect 19966 25342 20018 25394
rect 25118 25342 25170 25394
rect 42254 25342 42306 25394
rect 15822 25230 15874 25282
rect 19182 25230 19234 25282
rect 20302 25230 20354 25282
rect 21310 25230 21362 25282
rect 25454 25230 25506 25282
rect 28590 25230 28642 25282
rect 29262 25230 29314 25282
rect 35870 25230 35922 25282
rect 36542 25230 36594 25282
rect 41358 25230 41410 25282
rect 41918 25230 41970 25282
rect 44158 25230 44210 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 6974 24894 7026 24946
rect 7758 24894 7810 24946
rect 10334 24894 10386 24946
rect 10894 24894 10946 24946
rect 21310 24894 21362 24946
rect 21982 24894 22034 24946
rect 37998 24894 38050 24946
rect 17950 24782 18002 24834
rect 22542 24782 22594 24834
rect 25230 24782 25282 24834
rect 27246 24782 27298 24834
rect 27806 24782 27858 24834
rect 43038 24782 43090 24834
rect 8094 24670 8146 24722
rect 13358 24670 13410 24722
rect 13806 24670 13858 24722
rect 18062 24670 18114 24722
rect 18510 24670 18562 24722
rect 18846 24670 18898 24722
rect 25566 24670 25618 24722
rect 26126 24670 26178 24722
rect 27134 24670 27186 24722
rect 29038 24670 29090 24722
rect 34078 24670 34130 24722
rect 35086 24670 35138 24722
rect 35534 24670 35586 24722
rect 41470 24670 41522 24722
rect 42702 24670 42754 24722
rect 7198 24558 7250 24610
rect 8654 24558 8706 24610
rect 26462 24558 26514 24610
rect 29710 24558 29762 24610
rect 31838 24558 31890 24610
rect 32174 24558 32226 24610
rect 33742 24558 33794 24610
rect 34638 24558 34690 24610
rect 38334 24558 38386 24610
rect 41694 24558 41746 24610
rect 42254 24558 42306 24610
rect 22430 24446 22482 24498
rect 32286 24446 32338 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 19406 24110 19458 24162
rect 19742 24110 19794 24162
rect 8766 23998 8818 24050
rect 15486 23998 15538 24050
rect 24782 23998 24834 24050
rect 26910 23998 26962 24050
rect 29262 23998 29314 24050
rect 32958 23998 33010 24050
rect 33294 23998 33346 24050
rect 44046 23998 44098 24050
rect 7198 23886 7250 23938
rect 7758 23886 7810 23938
rect 8542 23886 8594 23938
rect 12462 23886 12514 23938
rect 18286 23886 18338 23938
rect 18846 23886 18898 23938
rect 24110 23886 24162 23938
rect 29486 23886 29538 23938
rect 29598 23886 29650 23938
rect 30046 23886 30098 23938
rect 34974 23886 35026 23938
rect 35198 23886 35250 23938
rect 35422 23886 35474 23938
rect 37550 23886 37602 23938
rect 40686 23886 40738 23938
rect 41246 23886 41298 23938
rect 7870 23774 7922 23826
rect 9214 23774 9266 23826
rect 9550 23774 9602 23826
rect 9886 23774 9938 23826
rect 16046 23774 16098 23826
rect 19294 23774 19346 23826
rect 19854 23774 19906 23826
rect 29150 23774 29202 23826
rect 30830 23774 30882 23826
rect 36318 23774 36370 23826
rect 37214 23774 37266 23826
rect 43486 23774 43538 23826
rect 6190 23662 6242 23714
rect 6526 23662 6578 23714
rect 12798 23662 12850 23714
rect 20302 23662 20354 23714
rect 28142 23662 28194 23714
rect 33406 23662 33458 23714
rect 35310 23662 35362 23714
rect 35534 23662 35586 23714
rect 36206 23662 36258 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 13582 23326 13634 23378
rect 21534 23326 21586 23378
rect 30830 23326 30882 23378
rect 31614 23326 31666 23378
rect 35534 23326 35586 23378
rect 39790 23326 39842 23378
rect 8654 23214 8706 23266
rect 20190 23214 20242 23266
rect 20862 23214 20914 23266
rect 21198 23214 21250 23266
rect 31054 23214 31106 23266
rect 35086 23214 35138 23266
rect 36542 23214 36594 23266
rect 36990 23214 37042 23266
rect 37886 23214 37938 23266
rect 42478 23214 42530 23266
rect 43822 23214 43874 23266
rect 6078 23102 6130 23154
rect 6414 23102 6466 23154
rect 7198 23102 7250 23154
rect 7758 23102 7810 23154
rect 7870 23102 7922 23154
rect 8318 23102 8370 23154
rect 10782 23102 10834 23154
rect 11230 23102 11282 23154
rect 17838 23102 17890 23154
rect 18398 23102 18450 23154
rect 19182 23102 19234 23154
rect 19518 23102 19570 23154
rect 20526 23102 20578 23154
rect 21758 23102 21810 23154
rect 25342 23102 25394 23154
rect 28478 23102 28530 23154
rect 28702 23102 28754 23154
rect 28926 23102 28978 23154
rect 29038 23102 29090 23154
rect 30382 23102 30434 23154
rect 30606 23102 30658 23154
rect 31166 23102 31218 23154
rect 31838 23102 31890 23154
rect 32398 23102 32450 23154
rect 35310 23102 35362 23154
rect 35982 23102 36034 23154
rect 36318 23102 36370 23154
rect 36766 23102 36818 23154
rect 37774 23102 37826 23154
rect 38894 23102 38946 23154
rect 41582 23102 41634 23154
rect 42814 23102 42866 23154
rect 43262 23102 43314 23154
rect 44158 23102 44210 23154
rect 5518 22990 5570 23042
rect 14142 22990 14194 23042
rect 26014 22990 26066 23042
rect 28142 22990 28194 23042
rect 28814 22990 28866 23042
rect 29710 22990 29762 23042
rect 34974 22990 35026 23042
rect 36430 22990 36482 23042
rect 38446 22990 38498 23042
rect 40350 22990 40402 23042
rect 41694 22990 41746 23042
rect 18510 22878 18562 22930
rect 30046 22878 30098 22930
rect 30382 22878 30434 22930
rect 35870 22878 35922 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 10446 22542 10498 22594
rect 11790 22542 11842 22594
rect 18846 22542 18898 22594
rect 19294 22542 19346 22594
rect 34974 22542 35026 22594
rect 38558 22542 38610 22594
rect 12798 22430 12850 22482
rect 15262 22430 15314 22482
rect 19294 22430 19346 22482
rect 23998 22430 24050 22482
rect 29598 22430 29650 22482
rect 33070 22430 33122 22482
rect 33966 22430 34018 22482
rect 42366 22430 42418 22482
rect 44270 22430 44322 22482
rect 4846 22318 4898 22370
rect 5966 22318 6018 22370
rect 6526 22318 6578 22370
rect 6974 22318 7026 22370
rect 7422 22318 7474 22370
rect 10894 22318 10946 22370
rect 12350 22318 12402 22370
rect 12686 22318 12738 22370
rect 13582 22318 13634 22370
rect 18174 22318 18226 22370
rect 20414 22318 20466 22370
rect 21758 22318 21810 22370
rect 23774 22318 23826 22370
rect 25566 22318 25618 22370
rect 26686 22318 26738 22370
rect 27134 22318 27186 22370
rect 28254 22318 28306 22370
rect 30270 22318 30322 22370
rect 33742 22318 33794 22370
rect 34190 22318 34242 22370
rect 35198 22318 35250 22370
rect 35422 22318 35474 22370
rect 35646 22318 35698 22370
rect 36990 22318 37042 22370
rect 37438 22318 37490 22370
rect 39118 22318 39170 22370
rect 39454 22318 39506 22370
rect 9662 22206 9714 22258
rect 11678 22206 11730 22258
rect 12462 22206 12514 22258
rect 12798 22206 12850 22258
rect 17390 22206 17442 22258
rect 22094 22206 22146 22258
rect 22542 22206 22594 22258
rect 24110 22206 24162 22258
rect 25790 22206 25842 22258
rect 27470 22206 27522 22258
rect 28590 22206 28642 22258
rect 29486 22206 29538 22258
rect 30942 22206 30994 22258
rect 34414 22206 34466 22258
rect 37214 22206 37266 22258
rect 38670 22206 38722 22258
rect 5070 22094 5122 22146
rect 10670 22094 10722 22146
rect 13694 22094 13746 22146
rect 13806 22094 13858 22146
rect 13918 22094 13970 22146
rect 14030 22094 14082 22146
rect 19742 22094 19794 22146
rect 20190 22094 20242 22146
rect 21422 22094 21474 22146
rect 23102 22094 23154 22146
rect 26350 22094 26402 22146
rect 29710 22094 29762 22146
rect 34302 22094 34354 22146
rect 35086 22094 35138 22146
rect 37326 22094 37378 22146
rect 37550 22094 37602 22146
rect 41918 22094 41970 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 11006 21758 11058 21810
rect 12910 21758 12962 21810
rect 15486 21758 15538 21810
rect 17502 21758 17554 21810
rect 18846 21758 18898 21810
rect 30942 21758 30994 21810
rect 36094 21758 36146 21810
rect 39790 21758 39842 21810
rect 6638 21646 6690 21698
rect 7646 21646 7698 21698
rect 10558 21646 10610 21698
rect 14478 21646 14530 21698
rect 15822 21646 15874 21698
rect 15934 21646 15986 21698
rect 16494 21646 16546 21698
rect 17726 21646 17778 21698
rect 19630 21646 19682 21698
rect 28590 21646 28642 21698
rect 34414 21646 34466 21698
rect 34974 21646 35026 21698
rect 36542 21646 36594 21698
rect 3950 21534 4002 21586
rect 4398 21534 4450 21586
rect 7758 21534 7810 21586
rect 11342 21534 11394 21586
rect 11566 21534 11618 21586
rect 11790 21534 11842 21586
rect 12014 21534 12066 21586
rect 13134 21534 13186 21586
rect 13358 21534 13410 21586
rect 14142 21534 14194 21586
rect 14254 21534 14306 21586
rect 14702 21534 14754 21586
rect 16382 21534 16434 21586
rect 16942 21534 16994 21586
rect 17278 21534 17330 21586
rect 17950 21534 18002 21586
rect 18734 21534 18786 21586
rect 19406 21534 19458 21586
rect 19966 21534 20018 21586
rect 25342 21534 25394 21586
rect 28478 21534 28530 21586
rect 29150 21534 29202 21586
rect 31278 21534 31330 21586
rect 31726 21534 31778 21586
rect 33966 21534 34018 21586
rect 34190 21534 34242 21586
rect 34638 21534 34690 21586
rect 35422 21534 35474 21586
rect 36430 21534 36482 21586
rect 36654 21534 36706 21586
rect 36878 21534 36930 21586
rect 37102 21534 37154 21586
rect 41918 21534 41970 21586
rect 7198 21422 7250 21474
rect 10894 21422 10946 21474
rect 11902 21422 11954 21474
rect 13470 21422 13522 21474
rect 14366 21422 14418 21474
rect 15374 21422 15426 21474
rect 16718 21422 16770 21474
rect 20750 21422 20802 21474
rect 22878 21422 22930 21474
rect 26014 21422 26066 21474
rect 28142 21422 28194 21474
rect 29598 21422 29650 21474
rect 40238 21422 40290 21474
rect 41694 21422 41746 21474
rect 10446 21310 10498 21362
rect 12462 21310 12514 21362
rect 12574 21310 12626 21362
rect 18622 21310 18674 21362
rect 28590 21310 28642 21362
rect 29150 21310 29202 21362
rect 29598 21310 29650 21362
rect 34078 21310 34130 21362
rect 35198 21310 35250 21362
rect 35646 21310 35698 21362
rect 42254 21310 42306 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 13694 20974 13746 21026
rect 19294 20974 19346 21026
rect 21534 20974 21586 21026
rect 26350 20974 26402 21026
rect 31502 20974 31554 21026
rect 31838 20974 31890 21026
rect 35870 20974 35922 21026
rect 4398 20862 4450 20914
rect 5966 20862 6018 20914
rect 15374 20862 15426 20914
rect 17502 20862 17554 20914
rect 19182 20862 19234 20914
rect 27918 20862 27970 20914
rect 33966 20862 34018 20914
rect 35310 20862 35362 20914
rect 35982 20862 36034 20914
rect 37102 20862 37154 20914
rect 41470 20862 41522 20914
rect 42366 20862 42418 20914
rect 6078 20750 6130 20802
rect 11566 20750 11618 20802
rect 12014 20750 12066 20802
rect 13918 20750 13970 20802
rect 14142 20750 14194 20802
rect 18174 20750 18226 20802
rect 18958 20750 19010 20802
rect 20526 20750 20578 20802
rect 21870 20750 21922 20802
rect 25342 20750 25394 20802
rect 26014 20750 26066 20802
rect 27134 20750 27186 20802
rect 27806 20750 27858 20802
rect 29822 20750 29874 20802
rect 30046 20750 30098 20802
rect 30606 20750 30658 20802
rect 32286 20750 32338 20802
rect 33070 20750 33122 20802
rect 33854 20750 33906 20802
rect 34750 20750 34802 20802
rect 34974 20750 35026 20802
rect 38110 20750 38162 20802
rect 38670 20750 38722 20802
rect 42926 20750 42978 20802
rect 43486 20750 43538 20802
rect 5070 20638 5122 20690
rect 5630 20638 5682 20690
rect 9214 20638 9266 20690
rect 13470 20638 13522 20690
rect 14590 20638 14642 20690
rect 19742 20638 19794 20690
rect 20078 20638 20130 20690
rect 20750 20638 20802 20690
rect 22094 20638 22146 20690
rect 22654 20638 22706 20690
rect 23214 20638 23266 20690
rect 26910 20638 26962 20690
rect 28142 20638 28194 20690
rect 29262 20638 29314 20690
rect 29486 20638 29538 20690
rect 30494 20638 30546 20690
rect 32398 20638 32450 20690
rect 34190 20638 34242 20690
rect 34414 20638 34466 20690
rect 35198 20638 35250 20690
rect 37214 20638 37266 20690
rect 37662 20638 37714 20690
rect 4286 20526 4338 20578
rect 4734 20526 4786 20578
rect 8430 20526 8482 20578
rect 25566 20526 25618 20578
rect 29598 20526 29650 20578
rect 30270 20526 30322 20578
rect 33406 20526 33458 20578
rect 33966 20526 34018 20578
rect 35422 20526 35474 20578
rect 36430 20526 36482 20578
rect 37102 20526 37154 20578
rect 37438 20526 37490 20578
rect 41134 20526 41186 20578
rect 43262 20526 43314 20578
rect 44270 20526 44322 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 4846 20190 4898 20242
rect 11454 20190 11506 20242
rect 14478 20190 14530 20242
rect 26574 20190 26626 20242
rect 35534 20190 35586 20242
rect 39118 20190 39170 20242
rect 5630 20078 5682 20130
rect 11342 20078 11394 20130
rect 12350 20078 12402 20130
rect 12574 20078 12626 20130
rect 12686 20078 12738 20130
rect 12910 20078 12962 20130
rect 14254 20078 14306 20130
rect 17838 20078 17890 20130
rect 19182 20078 19234 20130
rect 20638 20078 20690 20130
rect 25902 20078 25954 20130
rect 26798 20078 26850 20130
rect 27918 20078 27970 20130
rect 29262 20078 29314 20130
rect 31726 20078 31778 20130
rect 32062 20078 32114 20130
rect 32510 20078 32562 20130
rect 33070 20078 33122 20130
rect 34190 20078 34242 20130
rect 40014 20078 40066 20130
rect 40350 20078 40402 20130
rect 40910 20078 40962 20130
rect 43822 20078 43874 20130
rect 2046 19966 2098 20018
rect 2606 19966 2658 20018
rect 12014 19966 12066 20018
rect 12126 19966 12178 20018
rect 13358 19966 13410 20018
rect 14590 19966 14642 20018
rect 14702 19966 14754 20018
rect 14814 19966 14866 20018
rect 17614 19966 17666 20018
rect 18286 19966 18338 20018
rect 19406 19966 19458 20018
rect 19966 19966 20018 20018
rect 25790 19966 25842 20018
rect 26126 19966 26178 20018
rect 27022 19966 27074 20018
rect 27582 19966 27634 20018
rect 28590 19966 28642 20018
rect 33406 19966 33458 20018
rect 33966 19966 34018 20018
rect 34638 19966 34690 20018
rect 35198 19966 35250 20018
rect 35422 19966 35474 20018
rect 35646 19966 35698 20018
rect 35982 19966 36034 20018
rect 36542 19966 36594 20018
rect 39678 19966 39730 20018
rect 41806 19966 41858 20018
rect 42814 19966 42866 20018
rect 44158 19966 44210 20018
rect 13806 19854 13858 19906
rect 15262 19854 15314 19906
rect 22766 19854 22818 19906
rect 31390 19854 31442 19906
rect 32398 19854 32450 19906
rect 34414 19854 34466 19906
rect 34974 19854 35026 19906
rect 41694 19854 41746 19906
rect 42590 19854 42642 19906
rect 15374 19742 15426 19794
rect 18622 19742 18674 19794
rect 42702 19742 42754 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 27134 19406 27186 19458
rect 28254 19406 28306 19458
rect 32846 19406 32898 19458
rect 36990 19406 37042 19458
rect 6526 19294 6578 19346
rect 12238 19294 12290 19346
rect 14142 19294 14194 19346
rect 18174 19294 18226 19346
rect 20302 19294 20354 19346
rect 22094 19294 22146 19346
rect 28366 19294 28418 19346
rect 29934 19294 29986 19346
rect 32062 19294 32114 19346
rect 33966 19294 34018 19346
rect 36094 19294 36146 19346
rect 37102 19294 37154 19346
rect 44046 19294 44098 19346
rect 3278 19182 3330 19234
rect 4622 19182 4674 19234
rect 4958 19182 5010 19234
rect 5070 19182 5122 19234
rect 5966 19182 6018 19234
rect 6862 19182 6914 19234
rect 11902 19182 11954 19234
rect 17054 19182 17106 19234
rect 17390 19182 17442 19234
rect 22318 19182 22370 19234
rect 27246 19182 27298 19234
rect 29150 19182 29202 19234
rect 32846 19182 32898 19234
rect 33294 19182 33346 19234
rect 40686 19182 40738 19234
rect 41134 19182 41186 19234
rect 3166 19070 3218 19122
rect 7422 19070 7474 19122
rect 12126 19070 12178 19122
rect 16270 19070 16322 19122
rect 21982 19070 22034 19122
rect 27918 19070 27970 19122
rect 32510 19070 32562 19122
rect 40238 19070 40290 19122
rect 5630 18958 5682 19010
rect 12350 18958 12402 19010
rect 12462 18958 12514 19010
rect 20750 18958 20802 19010
rect 27134 18958 27186 19010
rect 27582 18958 27634 19010
rect 28478 18958 28530 19010
rect 40350 18958 40402 19010
rect 43486 18958 43538 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 1598 18622 1650 18674
rect 2382 18622 2434 18674
rect 15710 18622 15762 18674
rect 15822 18622 15874 18674
rect 43374 18622 43426 18674
rect 7646 18510 7698 18562
rect 8318 18510 8370 18562
rect 10446 18510 10498 18562
rect 10670 18510 10722 18562
rect 15038 18510 15090 18562
rect 15598 18510 15650 18562
rect 17502 18510 17554 18562
rect 17614 18510 17666 18562
rect 18286 18510 18338 18562
rect 24110 18510 24162 18562
rect 25230 18510 25282 18562
rect 28366 18510 28418 18562
rect 29486 18510 29538 18562
rect 29934 18510 29986 18562
rect 32398 18510 32450 18562
rect 33406 18510 33458 18562
rect 35870 18510 35922 18562
rect 36654 18510 36706 18562
rect 41246 18510 41298 18562
rect 4734 18398 4786 18450
rect 5182 18398 5234 18450
rect 6638 18398 6690 18450
rect 7198 18398 7250 18450
rect 7870 18398 7922 18450
rect 8542 18398 8594 18450
rect 10894 18398 10946 18450
rect 11118 18398 11170 18450
rect 11678 18398 11730 18450
rect 12574 18398 12626 18450
rect 13694 18398 13746 18450
rect 14478 18398 14530 18450
rect 14814 18398 14866 18450
rect 16270 18398 16322 18450
rect 17278 18398 17330 18450
rect 18622 18398 18674 18450
rect 20638 18398 20690 18450
rect 21198 18398 21250 18450
rect 24446 18398 24498 18450
rect 25454 18398 25506 18450
rect 26462 18398 26514 18450
rect 26910 18398 26962 18450
rect 28254 18398 28306 18450
rect 29262 18398 29314 18450
rect 30158 18398 30210 18450
rect 31054 18398 31106 18450
rect 31166 18398 31218 18450
rect 31838 18398 31890 18450
rect 32174 18398 32226 18450
rect 33070 18398 33122 18450
rect 34078 18398 34130 18450
rect 34302 18398 34354 18450
rect 34638 18398 34690 18450
rect 34862 18398 34914 18450
rect 35310 18398 35362 18450
rect 35534 18398 35586 18450
rect 36206 18398 36258 18450
rect 36542 18398 36594 18450
rect 40014 18398 40066 18450
rect 42030 18398 42082 18450
rect 42702 18398 42754 18450
rect 43038 18398 43090 18450
rect 6414 18286 6466 18338
rect 10558 18286 10610 18338
rect 11454 18286 11506 18338
rect 11902 18286 11954 18338
rect 14926 18286 14978 18338
rect 21758 18286 21810 18338
rect 26350 18286 26402 18338
rect 27918 18286 27970 18338
rect 28926 18286 28978 18338
rect 29598 18286 29650 18338
rect 30718 18286 30770 18338
rect 32510 18286 32562 18338
rect 34526 18286 34578 18338
rect 35086 18286 35138 18338
rect 37102 18286 37154 18338
rect 40126 18286 40178 18338
rect 42254 18286 42306 18338
rect 12126 18174 12178 18226
rect 13806 18174 13858 18226
rect 20974 18174 21026 18226
rect 26126 18174 26178 18226
rect 41134 18174 41186 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 9774 17838 9826 17890
rect 11454 17838 11506 17890
rect 27694 17838 27746 17890
rect 37102 17838 37154 17890
rect 5966 17726 6018 17778
rect 9662 17726 9714 17778
rect 11678 17726 11730 17778
rect 12014 17726 12066 17778
rect 13470 17726 13522 17778
rect 15598 17726 15650 17778
rect 22318 17726 22370 17778
rect 23438 17726 23490 17778
rect 24670 17726 24722 17778
rect 26798 17726 26850 17778
rect 28142 17726 28194 17778
rect 36430 17726 36482 17778
rect 37550 17726 37602 17778
rect 42142 17726 42194 17778
rect 8878 17614 8930 17666
rect 9326 17614 9378 17666
rect 10334 17614 10386 17666
rect 16270 17614 16322 17666
rect 16606 17614 16658 17666
rect 16942 17614 16994 17666
rect 19182 17614 19234 17666
rect 19854 17614 19906 17666
rect 20302 17614 20354 17666
rect 20526 17614 20578 17666
rect 20862 17614 20914 17666
rect 21534 17614 21586 17666
rect 21870 17614 21922 17666
rect 23998 17614 24050 17666
rect 27134 17614 27186 17666
rect 27358 17614 27410 17666
rect 32286 17614 32338 17666
rect 33070 17614 33122 17666
rect 33518 17614 33570 17666
rect 38894 17614 38946 17666
rect 39342 17614 39394 17666
rect 42590 17614 42642 17666
rect 6526 17502 6578 17554
rect 18846 17502 18898 17554
rect 19518 17502 19570 17554
rect 21310 17502 21362 17554
rect 22206 17502 22258 17554
rect 22430 17502 22482 17554
rect 22990 17502 23042 17554
rect 28030 17502 28082 17554
rect 34302 17502 34354 17554
rect 36990 17502 37042 17554
rect 10110 17390 10162 17442
rect 11902 17390 11954 17442
rect 12126 17390 12178 17442
rect 16830 17390 16882 17442
rect 17502 17390 17554 17442
rect 17838 17390 17890 17442
rect 20526 17390 20578 17442
rect 21422 17390 21474 17442
rect 22878 17390 22930 17442
rect 28254 17390 28306 17442
rect 29374 17390 29426 17442
rect 32510 17390 32562 17442
rect 32846 17390 32898 17442
rect 37438 17390 37490 17442
rect 41806 17390 41858 17442
rect 42926 17390 42978 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 6078 17054 6130 17106
rect 18286 17054 18338 17106
rect 18510 17054 18562 17106
rect 23886 17054 23938 17106
rect 25342 17054 25394 17106
rect 27806 17054 27858 17106
rect 30830 17054 30882 17106
rect 39790 17054 39842 17106
rect 40350 17054 40402 17106
rect 41918 17054 41970 17106
rect 43822 17054 43874 17106
rect 13134 16942 13186 16994
rect 23438 16942 23490 16994
rect 26462 16942 26514 16994
rect 28254 16942 28306 16994
rect 34190 16942 34242 16994
rect 5294 16830 5346 16882
rect 8318 16830 8370 16882
rect 8990 16830 9042 16882
rect 9998 16830 10050 16882
rect 10670 16830 10722 16882
rect 13358 16830 13410 16882
rect 14030 16830 14082 16882
rect 19070 16830 19122 16882
rect 19406 16830 19458 16882
rect 22878 16830 22930 16882
rect 23998 16830 24050 16882
rect 24782 16830 24834 16882
rect 25678 16830 25730 16882
rect 26350 16830 26402 16882
rect 27470 16830 27522 16882
rect 28478 16830 28530 16882
rect 29934 16830 29986 16882
rect 33406 16830 33458 16882
rect 36766 16830 36818 16882
rect 37326 16830 37378 16882
rect 42142 16830 42194 16882
rect 43598 16830 43650 16882
rect 44158 16830 44210 16882
rect 12798 16718 12850 16770
rect 14702 16718 14754 16770
rect 16830 16718 16882 16770
rect 20190 16718 20242 16770
rect 22318 16718 22370 16770
rect 23102 16718 23154 16770
rect 27806 16718 27858 16770
rect 29486 16718 29538 16770
rect 36318 16718 36370 16770
rect 23886 16606 23938 16658
rect 28814 16606 28866 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 7198 16270 7250 16322
rect 9886 16270 9938 16322
rect 12798 16270 12850 16322
rect 15934 16270 15986 16322
rect 26910 16270 26962 16322
rect 29150 16270 29202 16322
rect 33966 16270 34018 16322
rect 34302 16270 34354 16322
rect 7086 16158 7138 16210
rect 9102 16158 9154 16210
rect 10446 16158 10498 16210
rect 11230 16158 11282 16210
rect 12462 16158 12514 16210
rect 17278 16158 17330 16210
rect 18846 16158 18898 16210
rect 19966 16158 20018 16210
rect 21758 16158 21810 16210
rect 23438 16158 23490 16210
rect 29710 16158 29762 16210
rect 33070 16158 33122 16210
rect 43934 16158 43986 16210
rect 10110 16046 10162 16098
rect 10334 16046 10386 16098
rect 15150 16046 15202 16098
rect 16606 16046 16658 16098
rect 19070 16046 19122 16098
rect 19742 16046 19794 16098
rect 20078 16046 20130 16098
rect 20750 16046 20802 16098
rect 21310 16046 21362 16098
rect 21646 16046 21698 16098
rect 21870 16046 21922 16098
rect 23102 16046 23154 16098
rect 23886 16046 23938 16098
rect 25342 16046 25394 16098
rect 25790 16046 25842 16098
rect 27918 16046 27970 16098
rect 28478 16046 28530 16098
rect 29486 16046 29538 16098
rect 31950 16046 32002 16098
rect 32510 16046 32562 16098
rect 34302 16046 34354 16098
rect 39342 16046 39394 16098
rect 40014 16046 40066 16098
rect 40686 16046 40738 16098
rect 41134 16046 41186 16098
rect 9550 15934 9602 15986
rect 11790 15934 11842 15986
rect 12238 15934 12290 15986
rect 14142 15934 14194 15986
rect 14478 15934 14530 15986
rect 14814 15934 14866 15986
rect 16718 15934 16770 15986
rect 22206 15934 22258 15986
rect 24894 15934 24946 15986
rect 30046 15934 30098 15986
rect 40238 15934 40290 15986
rect 43374 15934 43426 15986
rect 9438 15822 9490 15874
rect 10558 15822 10610 15874
rect 11118 15822 11170 15874
rect 13470 15822 13522 15874
rect 13806 15822 13858 15874
rect 15598 15822 15650 15874
rect 17726 15822 17778 15874
rect 19406 15822 19458 15874
rect 20526 15822 20578 15874
rect 20638 15822 20690 15874
rect 22542 15822 22594 15874
rect 24446 15822 24498 15874
rect 28366 15822 28418 15874
rect 30382 15822 30434 15874
rect 30718 15822 30770 15874
rect 31054 15822 31106 15874
rect 31614 15822 31666 15874
rect 32286 15822 32338 15874
rect 38782 15822 38834 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 8766 15486 8818 15538
rect 13134 15486 13186 15538
rect 14142 15486 14194 15538
rect 14590 15486 14642 15538
rect 15150 15486 15202 15538
rect 19070 15486 19122 15538
rect 27022 15486 27074 15538
rect 30046 15486 30098 15538
rect 30606 15486 30658 15538
rect 32398 15486 32450 15538
rect 40910 15486 40962 15538
rect 8990 15374 9042 15426
rect 13358 15374 13410 15426
rect 15486 15374 15538 15426
rect 19518 15374 19570 15426
rect 24334 15374 24386 15426
rect 25230 15374 25282 15426
rect 25454 15374 25506 15426
rect 25678 15374 25730 15426
rect 26350 15374 26402 15426
rect 26798 15374 26850 15426
rect 27582 15374 27634 15426
rect 28142 15374 28194 15426
rect 28590 15374 28642 15426
rect 30382 15374 30434 15426
rect 31390 15374 31442 15426
rect 39902 15374 39954 15426
rect 8430 15262 8482 15314
rect 8878 15262 8930 15314
rect 9662 15262 9714 15314
rect 12686 15262 12738 15314
rect 19294 15262 19346 15314
rect 19630 15262 19682 15314
rect 19966 15262 20018 15314
rect 20750 15262 20802 15314
rect 24222 15262 24274 15314
rect 26126 15262 26178 15314
rect 27694 15262 27746 15314
rect 28478 15262 28530 15314
rect 31278 15262 31330 15314
rect 39678 15262 39730 15314
rect 41134 15262 41186 15314
rect 42478 15262 42530 15314
rect 43486 15262 43538 15314
rect 10334 15150 10386 15202
rect 12462 15150 12514 15202
rect 13246 15150 13298 15202
rect 22878 15150 22930 15202
rect 23662 15150 23714 15202
rect 29486 15150 29538 15202
rect 30494 15150 30546 15202
rect 39230 15150 39282 15202
rect 42030 15150 42082 15202
rect 43038 15150 43090 15202
rect 23326 15038 23378 15090
rect 25790 15038 25842 15090
rect 28590 15038 28642 15090
rect 32062 15038 32114 15090
rect 41918 15038 41970 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 13582 14702 13634 14754
rect 21310 14702 21362 14754
rect 26574 14702 26626 14754
rect 9774 14590 9826 14642
rect 11902 14590 11954 14642
rect 14254 14590 14306 14642
rect 21422 14590 21474 14642
rect 21870 14590 21922 14642
rect 25454 14590 25506 14642
rect 28254 14590 28306 14642
rect 31950 14590 32002 14642
rect 34078 14590 34130 14642
rect 34750 14590 34802 14642
rect 9102 14478 9154 14530
rect 12238 14478 12290 14530
rect 12574 14478 12626 14530
rect 13694 14478 13746 14530
rect 15150 14478 15202 14530
rect 18734 14478 18786 14530
rect 19182 14478 19234 14530
rect 19518 14478 19570 14530
rect 20078 14478 20130 14530
rect 20526 14478 20578 14530
rect 21646 14478 21698 14530
rect 22654 14478 22706 14530
rect 25790 14478 25842 14530
rect 26014 14478 26066 14530
rect 27806 14478 27858 14530
rect 28142 14478 28194 14530
rect 29150 14478 29202 14530
rect 30606 14478 30658 14530
rect 30942 14478 30994 14530
rect 31166 14478 31218 14530
rect 40798 14478 40850 14530
rect 41246 14478 41298 14530
rect 15486 14366 15538 14418
rect 15710 14366 15762 14418
rect 16718 14366 16770 14418
rect 20750 14366 20802 14418
rect 23326 14366 23378 14418
rect 26126 14366 26178 14418
rect 29262 14366 29314 14418
rect 30606 14366 30658 14418
rect 41806 14478 41858 14530
rect 42030 14478 42082 14530
rect 34414 14366 34466 14418
rect 34638 14366 34690 14418
rect 41582 14366 41634 14418
rect 12350 14254 12402 14306
rect 13022 14254 13074 14306
rect 13582 14254 13634 14306
rect 14814 14254 14866 14306
rect 16382 14254 16434 14306
rect 17166 14254 17218 14306
rect 18174 14254 18226 14306
rect 18622 14254 18674 14306
rect 18846 14254 18898 14306
rect 18958 14254 19010 14306
rect 21982 14254 22034 14306
rect 22206 14254 22258 14306
rect 28030 14254 28082 14306
rect 30270 14254 30322 14306
rect 30494 14254 30546 14306
rect 35758 14254 35810 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 17502 13918 17554 13970
rect 18734 13918 18786 13970
rect 19406 13918 19458 13970
rect 23102 13918 23154 13970
rect 25342 13918 25394 13970
rect 26238 13918 26290 13970
rect 27134 13918 27186 13970
rect 27358 13918 27410 13970
rect 28702 13918 28754 13970
rect 30830 13918 30882 13970
rect 39118 13918 39170 13970
rect 40014 13918 40066 13970
rect 42702 13918 42754 13970
rect 16606 13806 16658 13858
rect 18958 13806 19010 13858
rect 19070 13806 19122 13858
rect 20302 13806 20354 13858
rect 26574 13806 26626 13858
rect 27022 13806 27074 13858
rect 29150 13806 29202 13858
rect 30494 13806 30546 13858
rect 31502 13806 31554 13858
rect 31838 13806 31890 13858
rect 32062 13806 32114 13858
rect 33070 13806 33122 13858
rect 33406 13806 33458 13858
rect 34190 13806 34242 13858
rect 34750 13806 34802 13858
rect 35086 13806 35138 13858
rect 10894 13694 10946 13746
rect 15934 13694 15986 13746
rect 16494 13694 16546 13746
rect 20414 13694 20466 13746
rect 20862 13694 20914 13746
rect 22878 13694 22930 13746
rect 25566 13694 25618 13746
rect 26462 13694 26514 13746
rect 28366 13694 28418 13746
rect 28590 13694 28642 13746
rect 31278 13694 31330 13746
rect 34526 13694 34578 13746
rect 35422 13694 35474 13746
rect 35982 13694 36034 13746
rect 36654 13694 36706 13746
rect 40350 13694 40402 13746
rect 41246 13694 41298 13746
rect 42030 13694 42082 13746
rect 11678 13582 11730 13634
rect 13806 13582 13858 13634
rect 14254 13582 14306 13634
rect 19854 13582 19906 13634
rect 24782 13582 24834 13634
rect 34302 13582 34354 13634
rect 41806 13582 41858 13634
rect 43150 13582 43202 13634
rect 15598 13470 15650 13522
rect 32174 13470 32226 13522
rect 35422 13470 35474 13522
rect 39678 13470 39730 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19406 13134 19458 13186
rect 26686 13134 26738 13186
rect 36990 13134 37042 13186
rect 37438 13134 37490 13186
rect 15710 13022 15762 13074
rect 17838 13022 17890 13074
rect 19070 13022 19122 13074
rect 20190 13022 20242 13074
rect 20638 13022 20690 13074
rect 21982 13022 22034 13074
rect 22430 13022 22482 13074
rect 26126 13022 26178 13074
rect 29374 13022 29426 13074
rect 30046 13022 30098 13074
rect 31166 13022 31218 13074
rect 32062 13022 32114 13074
rect 34302 13022 34354 13074
rect 36430 13022 36482 13074
rect 37550 13022 37602 13074
rect 42366 13022 42418 13074
rect 43710 13022 43762 13074
rect 12798 12910 12850 12962
rect 14366 12910 14418 12962
rect 14926 12910 14978 12962
rect 18062 12910 18114 12962
rect 18398 12910 18450 12962
rect 18734 12910 18786 12962
rect 25790 12910 25842 12962
rect 27022 12910 27074 12962
rect 32622 12910 32674 12962
rect 33182 12910 33234 12962
rect 33630 12910 33682 12962
rect 38222 12910 38274 12962
rect 38670 12910 38722 12962
rect 42142 12910 42194 12962
rect 12462 12798 12514 12850
rect 19182 12798 19234 12850
rect 21646 12798 21698 12850
rect 21870 12798 21922 12850
rect 27246 12798 27298 12850
rect 32958 12798 33010 12850
rect 37102 12798 37154 12850
rect 43038 12798 43090 12850
rect 44158 12798 44210 12850
rect 14590 12686 14642 12738
rect 18286 12686 18338 12738
rect 22878 12686 22930 12738
rect 27694 12686 27746 12738
rect 28142 12686 28194 12738
rect 28590 12686 28642 12738
rect 31502 12686 31554 12738
rect 32846 12686 32898 12738
rect 41134 12686 41186 12738
rect 41694 12686 41746 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 17502 12350 17554 12402
rect 19406 12350 19458 12402
rect 21758 12350 21810 12402
rect 22990 12350 23042 12402
rect 23662 12350 23714 12402
rect 27022 12350 27074 12402
rect 30270 12350 30322 12402
rect 30606 12350 30658 12402
rect 36766 12350 36818 12402
rect 36990 12350 37042 12402
rect 38782 12350 38834 12402
rect 41134 12350 41186 12402
rect 44270 12350 44322 12402
rect 14702 12238 14754 12290
rect 18062 12238 18114 12290
rect 18398 12238 18450 12290
rect 19854 12238 19906 12290
rect 21422 12238 21474 12290
rect 22094 12238 22146 12290
rect 22430 12238 22482 12290
rect 28142 12238 28194 12290
rect 29150 12238 29202 12290
rect 29710 12238 29762 12290
rect 30942 12238 30994 12290
rect 38894 12238 38946 12290
rect 41470 12238 41522 12290
rect 43262 12238 43314 12290
rect 14030 12126 14082 12178
rect 19182 12126 19234 12178
rect 27918 12126 27970 12178
rect 28590 12126 28642 12178
rect 28926 12126 28978 12178
rect 32062 12126 32114 12178
rect 32286 12126 32338 12178
rect 32622 12126 32674 12178
rect 33070 12126 33122 12178
rect 36318 12126 36370 12178
rect 36542 12126 36594 12178
rect 42030 12126 42082 12178
rect 43486 12126 43538 12178
rect 16830 12014 16882 12066
rect 22878 12014 22930 12066
rect 27470 12014 27522 12066
rect 32398 12014 32450 12066
rect 33854 12014 33906 12066
rect 35982 12014 36034 12066
rect 36878 12014 36930 12066
rect 38110 12014 38162 12066
rect 42366 12014 42418 12066
rect 17838 11902 17890 11954
rect 22766 11902 22818 11954
rect 26910 11902 26962 11954
rect 27470 11902 27522 11954
rect 38222 11902 38274 11954
rect 42590 11902 42642 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 21758 11566 21810 11618
rect 22094 11566 22146 11618
rect 27694 11566 27746 11618
rect 38222 11566 38274 11618
rect 13582 11454 13634 11506
rect 16158 11454 16210 11506
rect 18286 11454 18338 11506
rect 20750 11454 20802 11506
rect 25678 11454 25730 11506
rect 31166 11454 31218 11506
rect 33854 11454 33906 11506
rect 35982 11454 36034 11506
rect 36430 11454 36482 11506
rect 38110 11454 38162 11506
rect 19070 11342 19122 11394
rect 22430 11342 22482 11394
rect 22766 11342 22818 11394
rect 29822 11342 29874 11394
rect 32622 11342 32674 11394
rect 33070 11342 33122 11394
rect 37102 11342 37154 11394
rect 37326 11342 37378 11394
rect 37550 11342 37602 11394
rect 37774 11342 37826 11394
rect 38894 11342 38946 11394
rect 39230 11342 39282 11394
rect 42590 11342 42642 11394
rect 12350 11230 12402 11282
rect 21534 11230 21586 11282
rect 23550 11230 23602 11282
rect 26574 11230 26626 11282
rect 27358 11230 27410 11282
rect 28030 11230 28082 11282
rect 28478 11230 28530 11282
rect 29486 11230 29538 11282
rect 30494 11230 30546 11282
rect 30606 11230 30658 11282
rect 12014 11118 12066 11170
rect 12238 11118 12290 11170
rect 12798 11118 12850 11170
rect 21646 11118 21698 11170
rect 22206 11118 22258 11170
rect 26910 11118 26962 11170
rect 29150 11118 29202 11170
rect 30158 11118 30210 11170
rect 30830 11118 30882 11170
rect 32398 11118 32450 11170
rect 36318 11118 36370 11170
rect 37214 11118 37266 11170
rect 41806 11118 41858 11170
rect 42366 11118 42418 11170
rect 42926 11118 42978 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 13134 10782 13186 10834
rect 15262 10782 15314 10834
rect 15822 10782 15874 10834
rect 23662 10782 23714 10834
rect 31278 10782 31330 10834
rect 33966 10782 34018 10834
rect 34078 10782 34130 10834
rect 35198 10782 35250 10834
rect 36094 10782 36146 10834
rect 38334 10782 38386 10834
rect 38446 10782 38498 10834
rect 41358 10782 41410 10834
rect 11006 10670 11058 10722
rect 11902 10670 11954 10722
rect 12798 10670 12850 10722
rect 13806 10670 13858 10722
rect 15374 10670 15426 10722
rect 21646 10670 21698 10722
rect 22206 10670 22258 10722
rect 23214 10670 23266 10722
rect 24558 10670 24610 10722
rect 28366 10670 28418 10722
rect 31054 10670 31106 10722
rect 31726 10670 31778 10722
rect 35310 10670 35362 10722
rect 35534 10670 35586 10722
rect 35982 10670 36034 10722
rect 37438 10670 37490 10722
rect 41022 10670 41074 10722
rect 11230 10558 11282 10610
rect 11678 10558 11730 10610
rect 12126 10558 12178 10610
rect 12574 10558 12626 10610
rect 14030 10558 14082 10610
rect 14478 10558 14530 10610
rect 15038 10558 15090 10610
rect 21198 10558 21250 10610
rect 21870 10558 21922 10610
rect 22766 10558 22818 10610
rect 22878 10558 22930 10610
rect 23438 10558 23490 10610
rect 23774 10558 23826 10610
rect 23998 10558 24050 10610
rect 27694 10558 27746 10610
rect 30830 10558 30882 10610
rect 34302 10558 34354 10610
rect 34526 10558 34578 10610
rect 34862 10558 34914 10610
rect 35086 10558 35138 10610
rect 35870 10558 35922 10610
rect 36990 10558 37042 10610
rect 37886 10558 37938 10610
rect 38110 10558 38162 10610
rect 11118 10446 11170 10498
rect 12014 10446 12066 10498
rect 13918 10446 13970 10498
rect 18398 10446 18450 10498
rect 20526 10446 20578 10498
rect 22094 10446 22146 10498
rect 23102 10446 23154 10498
rect 30494 10446 30546 10498
rect 30942 10446 30994 10498
rect 31838 10446 31890 10498
rect 34190 10446 34242 10498
rect 38222 10446 38274 10498
rect 41806 10446 41858 10498
rect 24446 10334 24498 10386
rect 41694 10334 41746 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 18734 9998 18786 10050
rect 37438 9998 37490 10050
rect 37662 9998 37714 10050
rect 10110 9886 10162 9938
rect 12238 9886 12290 9938
rect 14254 9886 14306 9938
rect 16382 9886 16434 9938
rect 17950 9886 18002 9938
rect 18846 9886 18898 9938
rect 21422 9886 21474 9938
rect 23438 9886 23490 9938
rect 25566 9886 25618 9938
rect 29934 9886 29986 9938
rect 32062 9886 32114 9938
rect 38334 9886 38386 9938
rect 38670 9886 38722 9938
rect 44046 9886 44098 9938
rect 9438 9774 9490 9826
rect 12574 9774 12626 9826
rect 12910 9774 12962 9826
rect 13470 9774 13522 9826
rect 17726 9774 17778 9826
rect 21534 9774 21586 9826
rect 21870 9774 21922 9826
rect 22766 9774 22818 9826
rect 29150 9774 29202 9826
rect 34526 9774 34578 9826
rect 35310 9774 35362 9826
rect 35646 9774 35698 9826
rect 37214 9774 37266 9826
rect 38110 9774 38162 9826
rect 38894 9774 38946 9826
rect 40686 9774 40738 9826
rect 41246 9774 41298 9826
rect 12798 9662 12850 9714
rect 18398 9662 18450 9714
rect 20638 9662 20690 9714
rect 21310 9662 21362 9714
rect 34638 9662 34690 9714
rect 35870 9662 35922 9714
rect 36990 9662 37042 9714
rect 43486 9662 43538 9714
rect 20750 9550 20802 9602
rect 32510 9550 32562 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 15822 9214 15874 9266
rect 23102 9214 23154 9266
rect 25454 9214 25506 9266
rect 33182 9214 33234 9266
rect 33742 9214 33794 9266
rect 34974 9214 35026 9266
rect 35086 9214 35138 9266
rect 35198 9214 35250 9266
rect 38670 9214 38722 9266
rect 43374 9214 43426 9266
rect 44158 9214 44210 9266
rect 11678 9102 11730 9154
rect 14030 9102 14082 9154
rect 19406 9102 19458 9154
rect 20638 9102 20690 9154
rect 24334 9102 24386 9154
rect 25790 9102 25842 9154
rect 27694 9102 27746 9154
rect 30942 9102 30994 9154
rect 31390 9102 31442 9154
rect 32174 9102 32226 9154
rect 33070 9102 33122 9154
rect 36542 9102 36594 9154
rect 37886 9102 37938 9154
rect 42478 9102 42530 9154
rect 12462 8990 12514 9042
rect 12798 8990 12850 9042
rect 13022 8990 13074 9042
rect 13134 8990 13186 9042
rect 13246 8990 13298 9042
rect 13470 8990 13522 9042
rect 14142 8990 14194 9042
rect 14926 8990 14978 9042
rect 15262 8990 15314 9042
rect 18174 8990 18226 9042
rect 18734 8990 18786 9042
rect 19518 8990 19570 9042
rect 19854 8990 19906 9042
rect 23214 8990 23266 9042
rect 25230 8990 25282 9042
rect 25678 8990 25730 9042
rect 26910 8990 26962 9042
rect 30606 8990 30658 9042
rect 31838 8990 31890 9042
rect 33406 8990 33458 9042
rect 35870 8990 35922 9042
rect 36318 8990 36370 9042
rect 36654 8990 36706 9042
rect 37214 8990 37266 9042
rect 38334 8990 38386 9042
rect 38558 8990 38610 9042
rect 38782 8990 38834 9042
rect 39006 8990 39058 9042
rect 42702 8990 42754 9042
rect 9550 8878 9602 8930
rect 15934 8878 15986 8930
rect 22766 8878 22818 8930
rect 25790 8878 25842 8930
rect 29822 8878 29874 8930
rect 34750 8878 34802 8930
rect 39454 8878 39506 8930
rect 41022 8878 41074 8930
rect 43710 8878 43762 8930
rect 15598 8766 15650 8818
rect 18398 8766 18450 8818
rect 24222 8766 24274 8818
rect 30270 8766 30322 8818
rect 34526 8766 34578 8818
rect 39342 8766 39394 8818
rect 40910 8766 40962 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 12798 8430 12850 8482
rect 17950 8430 18002 8482
rect 25678 8430 25730 8482
rect 42702 8430 42754 8482
rect 11230 8318 11282 8370
rect 12126 8318 12178 8370
rect 14030 8318 14082 8370
rect 18510 8318 18562 8370
rect 20302 8318 20354 8370
rect 21422 8318 21474 8370
rect 22542 8318 22594 8370
rect 29262 8318 29314 8370
rect 34862 8318 34914 8370
rect 35758 8318 35810 8370
rect 42142 8318 42194 8370
rect 42814 8318 42866 8370
rect 11342 8206 11394 8258
rect 11902 8206 11954 8258
rect 12238 8206 12290 8258
rect 12686 8206 12738 8258
rect 13694 8206 13746 8258
rect 14142 8206 14194 8258
rect 16046 8206 16098 8258
rect 17054 8206 17106 8258
rect 17390 8206 17442 8258
rect 17614 8206 17666 8258
rect 18846 8206 18898 8258
rect 19966 8206 20018 8258
rect 20414 8206 20466 8258
rect 21310 8206 21362 8258
rect 21758 8206 21810 8258
rect 22430 8206 22482 8258
rect 22878 8206 22930 8258
rect 25566 8206 25618 8258
rect 29934 8206 29986 8258
rect 30270 8206 30322 8258
rect 30606 8206 30658 8258
rect 32062 8206 32114 8258
rect 35198 8206 35250 8258
rect 35422 8206 35474 8258
rect 35870 8206 35922 8258
rect 38894 8206 38946 8258
rect 39342 8206 39394 8258
rect 43150 8206 43202 8258
rect 10894 8094 10946 8146
rect 11678 8094 11730 8146
rect 14366 8094 14418 8146
rect 15822 8094 15874 8146
rect 19070 8094 19122 8146
rect 19742 8094 19794 8146
rect 21982 8094 22034 8146
rect 22542 8094 22594 8146
rect 31278 8094 31330 8146
rect 32734 8094 32786 8146
rect 10782 7982 10834 8034
rect 12126 7982 12178 8034
rect 13918 7982 13970 8034
rect 18510 7982 18562 8034
rect 18622 7982 18674 8034
rect 20190 7982 20242 8034
rect 21534 7982 21586 8034
rect 22766 7982 22818 8034
rect 29598 7982 29650 8034
rect 30382 7982 30434 8034
rect 30830 7982 30882 8034
rect 30942 7982 30994 8034
rect 31054 7982 31106 8034
rect 35646 7982 35698 8034
rect 41806 7982 41858 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 13694 7646 13746 7698
rect 18846 7646 18898 7698
rect 19518 7646 19570 7698
rect 19742 7646 19794 7698
rect 22654 7646 22706 7698
rect 24670 7646 24722 7698
rect 28254 7646 28306 7698
rect 28814 7646 28866 7698
rect 32398 7646 32450 7698
rect 33182 7646 33234 7698
rect 33294 7646 33346 7698
rect 34078 7646 34130 7698
rect 35086 7646 35138 7698
rect 35870 7646 35922 7698
rect 39902 7646 39954 7698
rect 40910 7646 40962 7698
rect 43038 7646 43090 7698
rect 17502 7534 17554 7586
rect 18958 7534 19010 7586
rect 24558 7534 24610 7586
rect 29822 7534 29874 7586
rect 32622 7534 32674 7586
rect 33518 7534 33570 7586
rect 35758 7534 35810 7586
rect 10782 7422 10834 7474
rect 11230 7422 11282 7474
rect 16830 7422 16882 7474
rect 17950 7422 18002 7474
rect 18510 7422 18562 7474
rect 19630 7422 19682 7474
rect 19854 7422 19906 7474
rect 19966 7422 20018 7474
rect 22318 7422 22370 7474
rect 25230 7422 25282 7474
rect 25678 7422 25730 7474
rect 29150 7422 29202 7474
rect 32286 7422 32338 7474
rect 33070 7422 33122 7474
rect 34862 7422 34914 7474
rect 34974 7422 35026 7474
rect 35198 7422 35250 7474
rect 35422 7422 35474 7474
rect 36878 7422 36930 7474
rect 37438 7422 37490 7474
rect 42254 7422 42306 7474
rect 42702 7422 42754 7474
rect 43262 7422 43314 7474
rect 14030 7310 14082 7362
rect 16718 7310 16770 7362
rect 22766 7310 22818 7362
rect 31950 7310 32002 7362
rect 33966 7310 34018 7362
rect 41022 7310 41074 7362
rect 42030 7310 42082 7362
rect 22206 7198 22258 7250
rect 40462 7198 40514 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 16830 6862 16882 6914
rect 24894 6862 24946 6914
rect 43374 6862 43426 6914
rect 28590 6750 28642 6802
rect 30830 6750 30882 6802
rect 32958 6750 33010 6802
rect 36206 6750 36258 6802
rect 38670 6750 38722 6802
rect 8878 6638 8930 6690
rect 9326 6638 9378 6690
rect 12350 6638 12402 6690
rect 12574 6638 12626 6690
rect 12686 6638 12738 6690
rect 19966 6638 20018 6690
rect 20302 6638 20354 6690
rect 21422 6638 21474 6690
rect 21870 6638 21922 6690
rect 25118 6638 25170 6690
rect 25566 6638 25618 6690
rect 30046 6638 30098 6690
rect 33294 6638 33346 6690
rect 36990 6638 37042 6690
rect 38894 6638 38946 6690
rect 39790 6638 39842 6690
rect 40350 6638 40402 6690
rect 13806 6526 13858 6578
rect 14142 6526 14194 6578
rect 14478 6526 14530 6578
rect 15262 6526 15314 6578
rect 16606 6526 16658 6578
rect 34078 6526 34130 6578
rect 37102 6526 37154 6578
rect 37438 6526 37490 6578
rect 39454 6526 39506 6578
rect 42590 6526 42642 6578
rect 43598 6526 43650 6578
rect 43934 6526 43986 6578
rect 11790 6414 11842 6466
rect 14814 6414 14866 6466
rect 15150 6414 15202 6466
rect 16494 6414 16546 6466
rect 17614 6414 17666 6466
rect 24334 6414 24386 6466
rect 28142 6414 28194 6466
rect 37550 6414 37602 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 12238 6078 12290 6130
rect 13134 6078 13186 6130
rect 16382 6078 16434 6130
rect 18174 6078 18226 6130
rect 18846 6078 18898 6130
rect 23774 6078 23826 6130
rect 26910 6078 26962 6130
rect 28478 6078 28530 6130
rect 29150 6078 29202 6130
rect 32174 6078 32226 6130
rect 32622 6078 32674 6130
rect 33070 6078 33122 6130
rect 33182 6078 33234 6130
rect 33294 6078 33346 6130
rect 34190 6078 34242 6130
rect 37662 6078 37714 6130
rect 41470 6078 41522 6130
rect 43598 6078 43650 6130
rect 43822 6078 43874 6130
rect 17726 5966 17778 6018
rect 22990 5966 23042 6018
rect 25230 5966 25282 6018
rect 31278 5966 31330 6018
rect 31614 5966 31666 6018
rect 34302 5966 34354 6018
rect 42926 5966 42978 6018
rect 44158 5966 44210 6018
rect 12462 5854 12514 5906
rect 13358 5854 13410 5906
rect 13918 5854 13970 5906
rect 17838 5854 17890 5906
rect 18398 5854 18450 5906
rect 20190 5854 20242 5906
rect 20750 5854 20802 5906
rect 24446 5854 24498 5906
rect 27246 5854 27298 5906
rect 28030 5854 28082 5906
rect 28702 5854 28754 5906
rect 29374 5854 29426 5906
rect 33630 5854 33682 5906
rect 34750 5854 34802 5906
rect 35198 5854 35250 5906
rect 38670 5854 38722 5906
rect 38894 5854 38946 5906
rect 40910 5854 40962 5906
rect 42254 5854 42306 5906
rect 16718 5742 16770 5794
rect 19294 5742 19346 5794
rect 23998 5742 24050 5794
rect 27694 5742 27746 5794
rect 37998 5742 38050 5794
rect 42142 5742 42194 5794
rect 25342 5630 25394 5682
rect 38558 5630 38610 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 12350 5294 12402 5346
rect 14142 5294 14194 5346
rect 20862 5294 20914 5346
rect 22430 5294 22482 5346
rect 29374 5294 29426 5346
rect 12574 5182 12626 5234
rect 14254 5182 14306 5234
rect 21646 5182 21698 5234
rect 28142 5182 28194 5234
rect 29486 5182 29538 5234
rect 31054 5182 31106 5234
rect 33070 5182 33122 5234
rect 40350 5182 40402 5234
rect 41470 5182 41522 5234
rect 12686 5070 12738 5122
rect 14926 5070 14978 5122
rect 15710 5070 15762 5122
rect 16382 5070 16434 5122
rect 17390 5070 17442 5122
rect 17838 5070 17890 5122
rect 22206 5070 22258 5122
rect 25454 5070 25506 5122
rect 25902 5070 25954 5122
rect 27470 5070 27522 5122
rect 28366 5070 28418 5122
rect 30046 5070 30098 5122
rect 30606 5070 30658 5122
rect 35982 5070 36034 5122
rect 36430 5070 36482 5122
rect 37102 5070 37154 5122
rect 37550 5070 37602 5122
rect 41246 5070 41298 5122
rect 42142 5070 42194 5122
rect 42702 5070 42754 5122
rect 16606 4958 16658 5010
rect 20302 4846 20354 4898
rect 23214 4846 23266 4898
rect 33630 4846 33682 4898
rect 39790 4846 39842 4898
rect 42478 4846 42530 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 14814 4510 14866 4562
rect 16494 4510 16546 4562
rect 17950 4510 18002 4562
rect 25230 4510 25282 4562
rect 37214 4510 37266 4562
rect 37774 4510 37826 4562
rect 39790 4510 39842 4562
rect 41582 4510 41634 4562
rect 19070 4398 19122 4450
rect 39454 4398 39506 4450
rect 41694 4398 41746 4450
rect 12126 4286 12178 4338
rect 12462 4286 12514 4338
rect 16718 4286 16770 4338
rect 17390 4286 17442 4338
rect 19518 4286 19570 4338
rect 21534 4286 21586 4338
rect 22318 4286 22370 4338
rect 23774 4286 23826 4338
rect 24670 4286 24722 4338
rect 25454 4286 25506 4338
rect 28590 4286 28642 4338
rect 30830 4286 30882 4338
rect 34302 4286 34354 4338
rect 34750 4286 34802 4338
rect 37998 4286 38050 4338
rect 38670 4286 38722 4338
rect 15374 4174 15426 4226
rect 19854 4174 19906 4226
rect 21422 4174 21474 4226
rect 22990 4174 23042 4226
rect 24334 4174 24386 4226
rect 28142 4174 28194 4226
rect 29486 4174 29538 4226
rect 29934 4174 29986 4226
rect 30494 4174 30546 4226
rect 38446 4174 38498 4226
rect 41022 4174 41074 4226
rect 44270 4174 44322 4226
rect 21198 4062 21250 4114
rect 23102 4062 23154 4114
rect 28702 4062 28754 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 14478 3726 14530 3778
rect 35086 3726 35138 3778
rect 14254 3614 14306 3666
rect 35198 3614 35250 3666
rect 14030 3502 14082 3554
rect 21310 3502 21362 3554
rect 23102 3502 23154 3554
rect 37886 3502 37938 3554
rect 38558 3502 38610 3554
rect 21086 3390 21138 3442
rect 22878 3390 22930 3442
rect 37550 3390 37602 3442
rect 38222 3390 38274 3442
rect 43822 3390 43874 3442
rect 44158 3390 44210 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 41916 43092 41972 43102
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 32844 42084 32900 42094
rect 32844 41990 32900 42028
rect 34076 42084 34132 42094
rect 34076 41990 34132 42028
rect 40348 42084 40404 42094
rect 31612 41972 31668 41982
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 29932 41188 29988 41198
rect 29932 41094 29988 41132
rect 30156 41186 30212 41198
rect 30156 41134 30158 41186
rect 30210 41134 30212 41186
rect 29596 40964 29652 40974
rect 29596 40962 29876 40964
rect 29596 40910 29598 40962
rect 29650 40910 29876 40962
rect 29596 40908 29876 40910
rect 29596 40898 29652 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 26908 40516 26964 40526
rect 26908 40402 26964 40460
rect 26908 40350 26910 40402
rect 26962 40350 26964 40402
rect 26908 40338 26964 40350
rect 27244 40516 27300 40526
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 26796 39732 26852 39742
rect 26796 39638 26852 39676
rect 26684 39620 26740 39630
rect 26684 39526 26740 39564
rect 27020 39506 27076 39518
rect 27020 39454 27022 39506
rect 27074 39454 27076 39506
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 27020 38612 27076 39454
rect 27244 38834 27300 40460
rect 29260 40516 29316 40526
rect 28588 40404 28644 40414
rect 27580 40290 27636 40302
rect 27580 40238 27582 40290
rect 27634 40238 27636 40290
rect 27580 39730 27636 40238
rect 27692 40292 27748 40302
rect 27692 39842 27748 40236
rect 27692 39790 27694 39842
rect 27746 39790 27748 39842
rect 27692 39778 27748 39790
rect 27580 39678 27582 39730
rect 27634 39678 27636 39730
rect 27580 39666 27636 39678
rect 28588 39730 28644 40348
rect 28588 39678 28590 39730
rect 28642 39678 28644 39730
rect 28588 39666 28644 39678
rect 28364 39620 28420 39630
rect 28364 39526 28420 39564
rect 29260 39618 29316 40460
rect 29708 40404 29764 40414
rect 29820 40404 29876 40908
rect 30156 40628 30212 41134
rect 31276 41188 31332 41198
rect 30156 40572 30436 40628
rect 30044 40404 30100 40414
rect 29820 40402 30100 40404
rect 29820 40350 30046 40402
rect 30098 40350 30100 40402
rect 29820 40348 30100 40350
rect 29708 40290 29764 40348
rect 29708 40238 29710 40290
rect 29762 40238 29764 40290
rect 29708 40226 29764 40238
rect 29932 39732 29988 39742
rect 29932 39638 29988 39676
rect 29260 39566 29262 39618
rect 29314 39566 29316 39618
rect 29260 39554 29316 39566
rect 30044 39620 30100 40348
rect 30268 40404 30324 40414
rect 30268 40310 30324 40348
rect 30156 40292 30212 40302
rect 30156 40198 30212 40236
rect 30044 39554 30100 39564
rect 30380 39732 30436 40572
rect 30716 40404 30772 40414
rect 31276 40404 31332 41132
rect 30716 40402 30884 40404
rect 30716 40350 30718 40402
rect 30770 40350 30884 40402
rect 30716 40348 30884 40350
rect 30716 40338 30772 40348
rect 27468 39396 27524 39406
rect 28028 39396 28084 39406
rect 27468 39394 28028 39396
rect 27468 39342 27470 39394
rect 27522 39342 28028 39394
rect 27468 39340 28028 39342
rect 27468 39330 27524 39340
rect 28028 39302 28084 39340
rect 29036 39396 29092 39406
rect 27244 38782 27246 38834
rect 27298 38782 27300 38834
rect 27244 38770 27300 38782
rect 27020 38546 27076 38556
rect 27916 38722 27972 38734
rect 27916 38670 27918 38722
rect 27970 38670 27972 38722
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 27916 38164 27972 38670
rect 27916 38098 27972 38108
rect 29036 38724 29092 39340
rect 30156 39284 30212 39294
rect 30380 39284 30436 39676
rect 29820 39060 29876 39070
rect 29708 38948 29764 38958
rect 29036 38050 29092 38668
rect 29484 38836 29540 38846
rect 29260 38164 29316 38174
rect 29260 38070 29316 38108
rect 29036 37998 29038 38050
rect 29090 37998 29092 38050
rect 29036 37986 29092 37998
rect 29484 38050 29540 38780
rect 29484 37998 29486 38050
rect 29538 37998 29540 38050
rect 29484 37986 29540 37998
rect 29708 38050 29764 38892
rect 29708 37998 29710 38050
rect 29762 37998 29764 38050
rect 29708 37986 29764 37998
rect 29820 38724 29876 39004
rect 30044 38836 30100 38846
rect 30044 38722 30100 38780
rect 30044 38670 30046 38722
rect 30098 38670 30100 38722
rect 30044 38668 30100 38670
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 26236 37378 26292 37390
rect 26236 37326 26238 37378
rect 26290 37326 26292 37378
rect 26124 37266 26180 37278
rect 26124 37214 26126 37266
rect 26178 37214 26180 37266
rect 25228 37154 25284 37166
rect 25228 37102 25230 37154
rect 25282 37102 25284 37154
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 7308 36594 7364 36606
rect 7308 36542 7310 36594
rect 7362 36542 7364 36594
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 7308 35028 7364 36542
rect 10108 36482 10164 36494
rect 10108 36430 10110 36482
rect 10162 36430 10164 36482
rect 9436 36372 9492 36382
rect 9436 36278 9492 36316
rect 7308 34962 7364 34972
rect 9324 35028 9380 35038
rect 9324 34934 9380 34972
rect 8652 34916 8708 34926
rect 8652 34914 8820 34916
rect 8652 34862 8654 34914
rect 8706 34862 8820 34914
rect 8652 34860 8820 34862
rect 8652 34850 8708 34860
rect 8204 34242 8260 34254
rect 8652 34244 8708 34254
rect 8204 34190 8206 34242
rect 8258 34190 8260 34242
rect 7980 34130 8036 34142
rect 7980 34078 7982 34130
rect 8034 34078 8036 34130
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 6972 33460 7028 33470
rect 6972 33234 7028 33404
rect 7756 33460 7812 33470
rect 7756 33346 7812 33404
rect 7756 33294 7758 33346
rect 7810 33294 7812 33346
rect 7756 33282 7812 33294
rect 6972 33182 6974 33234
rect 7026 33182 7028 33234
rect 6076 32450 6132 32462
rect 6076 32398 6078 32450
rect 6130 32398 6132 32450
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 6076 31892 6132 32398
rect 6972 31948 7028 33182
rect 7308 33236 7364 33246
rect 7308 33142 7364 33180
rect 7980 32676 8036 34078
rect 7980 32610 8036 32620
rect 8204 32674 8260 34190
rect 8428 34242 8708 34244
rect 8428 34190 8654 34242
rect 8706 34190 8708 34242
rect 8428 34188 8708 34190
rect 8428 33458 8484 34188
rect 8652 34178 8708 34188
rect 8428 33406 8430 33458
rect 8482 33406 8484 33458
rect 8428 33394 8484 33406
rect 8764 33460 8820 34860
rect 8988 34132 9044 34142
rect 9884 34132 9940 34142
rect 8988 34130 9940 34132
rect 8988 34078 8990 34130
rect 9042 34078 9886 34130
rect 9938 34078 9940 34130
rect 8988 34076 9940 34078
rect 8988 34066 9044 34076
rect 9884 34066 9940 34076
rect 8876 33460 8932 33470
rect 8764 33404 8876 33460
rect 8204 32622 8206 32674
rect 8258 32622 8260 32674
rect 8204 32610 8260 32622
rect 8876 32562 8932 33404
rect 10108 33236 10164 36430
rect 15596 36482 15652 36494
rect 15596 36430 15598 36482
rect 15650 36430 15652 36482
rect 10444 36372 10500 36382
rect 10444 35924 10500 36316
rect 10332 35922 10500 35924
rect 10332 35870 10446 35922
rect 10498 35870 10500 35922
rect 10332 35868 10500 35870
rect 10332 34020 10388 35868
rect 10444 35858 10500 35868
rect 15596 35812 15652 36430
rect 16044 36484 16100 36494
rect 16044 36482 16324 36484
rect 16044 36430 16046 36482
rect 16098 36430 16324 36482
rect 16044 36428 16324 36430
rect 16044 36418 16100 36428
rect 15820 35812 15876 35822
rect 15596 35810 15876 35812
rect 15596 35758 15822 35810
rect 15874 35758 15876 35810
rect 15596 35756 15876 35758
rect 10780 35700 10836 35710
rect 15820 35700 15876 35756
rect 16156 35812 16212 35822
rect 16156 35718 16212 35756
rect 15820 35644 16100 35700
rect 10780 35606 10836 35644
rect 15820 35252 15876 35262
rect 11452 35028 11508 35038
rect 10556 35026 11508 35028
rect 10556 34974 11454 35026
rect 11506 34974 11508 35026
rect 10556 34972 11508 34974
rect 10556 34130 10612 34972
rect 11452 34962 11508 34972
rect 14588 34916 14644 34926
rect 11452 34356 11508 34366
rect 10556 34078 10558 34130
rect 10610 34078 10612 34130
rect 10556 34066 10612 34078
rect 11228 34242 11284 34254
rect 11228 34190 11230 34242
rect 11282 34190 11284 34242
rect 10108 33170 10164 33180
rect 10220 34018 10388 34020
rect 10220 33966 10334 34018
rect 10386 33966 10388 34018
rect 10220 33964 10388 33966
rect 10220 33012 10276 33964
rect 10332 33954 10388 33964
rect 9996 32956 10276 33012
rect 10556 33458 10612 33470
rect 10556 33406 10558 33458
rect 10610 33406 10612 33458
rect 9548 32676 9604 32686
rect 9548 32582 9604 32620
rect 8876 32510 8878 32562
rect 8930 32510 8932 32562
rect 8876 32498 8932 32510
rect 9996 32562 10052 32956
rect 9996 32510 9998 32562
rect 10050 32510 10052 32562
rect 6972 31892 7252 31948
rect 6076 31826 6132 31836
rect 7196 31778 7252 31892
rect 7980 31892 8036 31902
rect 7980 31798 8036 31836
rect 7196 31726 7198 31778
rect 7250 31726 7252 31778
rect 7196 31714 7252 31726
rect 8316 31106 8372 31118
rect 8316 31054 8318 31106
rect 8370 31054 8372 31106
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 8204 29540 8260 29550
rect 8316 29540 8372 31054
rect 8652 30996 8708 31006
rect 9548 30996 9604 31006
rect 8652 30994 9604 30996
rect 8652 30942 8654 30994
rect 8706 30942 9550 30994
rect 9602 30942 9604 30994
rect 8652 30940 9604 30942
rect 8652 30930 8708 30940
rect 9548 30930 9604 30940
rect 9996 30994 10052 32510
rect 10444 32564 10500 32574
rect 10556 32564 10612 33406
rect 10444 32562 10612 32564
rect 10444 32510 10446 32562
rect 10498 32510 10612 32562
rect 10444 32508 10612 32510
rect 10892 33236 10948 33246
rect 11228 33236 11284 34190
rect 10948 33180 11284 33236
rect 11452 34130 11508 34300
rect 11452 34078 11454 34130
rect 11506 34078 11508 34130
rect 10892 32562 10948 33180
rect 10892 32510 10894 32562
rect 10946 32510 10948 32562
rect 10444 32498 10500 32508
rect 10892 32498 10948 32510
rect 9996 30942 9998 30994
rect 10050 30942 10052 30994
rect 9996 30930 10052 30942
rect 10108 31890 10164 31902
rect 10108 31838 10110 31890
rect 10162 31838 10164 31890
rect 10108 30884 10164 31838
rect 11452 31778 11508 34078
rect 12684 34132 12740 34142
rect 12684 34038 12740 34076
rect 13132 34130 13188 34142
rect 13132 34078 13134 34130
rect 13186 34078 13188 34130
rect 11564 32562 11620 32574
rect 11564 32510 11566 32562
rect 11618 32510 11620 32562
rect 11564 32340 11620 32510
rect 13132 32564 13188 34078
rect 13132 32498 13188 32508
rect 13468 34132 13524 34142
rect 11564 32274 11620 32284
rect 11452 31726 11454 31778
rect 11506 31726 11508 31778
rect 11452 31714 11508 31726
rect 13468 31778 13524 34076
rect 14588 33570 14644 34860
rect 15820 34802 15876 35196
rect 16044 34916 16100 35644
rect 16156 34916 16212 34926
rect 16044 34914 16212 34916
rect 16044 34862 16158 34914
rect 16210 34862 16212 34914
rect 16044 34860 16212 34862
rect 16156 34850 16212 34860
rect 15820 34750 15822 34802
rect 15874 34750 15876 34802
rect 15820 34738 15876 34750
rect 15932 34804 15988 34814
rect 15932 34710 15988 34748
rect 15596 34690 15652 34702
rect 15596 34638 15598 34690
rect 15650 34638 15652 34690
rect 15372 34132 15428 34142
rect 15372 34130 15540 34132
rect 15372 34078 15374 34130
rect 15426 34078 15540 34130
rect 15372 34076 15540 34078
rect 15372 34066 15428 34076
rect 14588 33518 14590 33570
rect 14642 33518 14644 33570
rect 14588 33506 14644 33518
rect 15484 33124 15540 34076
rect 15596 33346 15652 34638
rect 16268 34354 16324 36428
rect 18284 36260 18340 36270
rect 17724 36258 18340 36260
rect 17724 36206 18286 36258
rect 18338 36206 18340 36258
rect 17724 36204 18340 36206
rect 17724 35922 17780 36204
rect 18284 36194 18340 36204
rect 19068 36258 19124 36270
rect 19068 36206 19070 36258
rect 19122 36206 19124 36258
rect 17724 35870 17726 35922
rect 17778 35870 17780 35922
rect 17724 35858 17780 35870
rect 17948 35924 18004 35934
rect 19068 35924 19124 36206
rect 16268 34302 16270 34354
rect 16322 34302 16324 34354
rect 16268 34290 16324 34302
rect 16492 35810 16548 35822
rect 16492 35758 16494 35810
rect 16546 35758 16548 35810
rect 16492 34132 16548 35758
rect 16716 35812 16772 35822
rect 16716 35698 16772 35756
rect 17500 35810 17556 35822
rect 17500 35758 17502 35810
rect 17554 35758 17556 35810
rect 16716 35646 16718 35698
rect 16770 35646 16772 35698
rect 16716 35634 16772 35646
rect 17388 35698 17444 35710
rect 17388 35646 17390 35698
rect 17442 35646 17444 35698
rect 16828 34916 16884 34926
rect 16828 34822 16884 34860
rect 17388 34804 17444 35646
rect 17500 35252 17556 35758
rect 17948 35700 18004 35868
rect 18732 35868 19124 35924
rect 19404 36258 19460 36270
rect 19404 36206 19406 36258
rect 19458 36206 19460 36258
rect 19404 35924 19460 36206
rect 23548 36260 23604 36270
rect 23548 36258 23716 36260
rect 23548 36206 23550 36258
rect 23602 36206 23716 36258
rect 23548 36204 23716 36206
rect 23548 36194 23604 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 17500 35186 17556 35196
rect 17836 35698 18004 35700
rect 17836 35646 17950 35698
rect 18002 35646 18004 35698
rect 17836 35644 18004 35646
rect 16492 34066 16548 34076
rect 17276 34132 17332 34142
rect 17276 34038 17332 34076
rect 15596 33294 15598 33346
rect 15650 33294 15652 33346
rect 15596 33282 15652 33294
rect 17388 33348 17444 34748
rect 17388 33282 17444 33292
rect 17724 34132 17780 34142
rect 17724 33346 17780 34076
rect 17724 33294 17726 33346
rect 17778 33294 17780 33346
rect 17724 33282 17780 33294
rect 15484 33068 15988 33124
rect 14028 32788 14084 32798
rect 14700 32788 14756 32798
rect 14028 32786 14756 32788
rect 14028 32734 14030 32786
rect 14082 32734 14702 32786
rect 14754 32734 14756 32786
rect 14028 32732 14756 32734
rect 14028 32722 14084 32732
rect 14700 32722 14756 32732
rect 15932 32786 15988 33068
rect 15932 32734 15934 32786
rect 15986 32734 15988 32786
rect 15932 32722 15988 32734
rect 14924 32676 14980 32686
rect 14812 32620 14924 32676
rect 14588 32564 14644 32574
rect 14588 32470 14644 32508
rect 13468 31726 13470 31778
rect 13522 31726 13524 31778
rect 13468 31714 13524 31726
rect 14028 31780 14084 31790
rect 14028 31778 14532 31780
rect 14028 31726 14030 31778
rect 14082 31726 14532 31778
rect 14028 31724 14532 31726
rect 14028 31714 14084 31724
rect 11116 31554 11172 31566
rect 11116 31502 11118 31554
rect 11170 31502 11172 31554
rect 10780 30996 10836 31006
rect 11116 30996 11172 31502
rect 13916 31220 13972 31230
rect 13916 31218 14420 31220
rect 13916 31166 13918 31218
rect 13970 31166 14420 31218
rect 13916 31164 14420 31166
rect 13916 31154 13972 31164
rect 10780 30994 11172 30996
rect 10780 30942 10782 30994
rect 10834 30942 11172 30994
rect 10780 30940 11172 30942
rect 11452 30994 11508 31006
rect 11452 30942 11454 30994
rect 11506 30942 11508 30994
rect 10332 30884 10388 30894
rect 10108 30882 10388 30884
rect 10108 30830 10334 30882
rect 10386 30830 10388 30882
rect 10108 30828 10388 30830
rect 10332 30818 10388 30828
rect 8204 29538 8372 29540
rect 8204 29486 8206 29538
rect 8258 29486 8372 29538
rect 8204 29484 8372 29486
rect 8204 29474 8260 29484
rect 8876 29428 8932 29438
rect 6076 29314 6132 29326
rect 6076 29262 6078 29314
rect 6130 29262 6132 29314
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 6076 28756 6132 29262
rect 6076 28690 6132 28700
rect 8316 28756 8372 28766
rect 8316 28662 8372 28700
rect 7644 28644 7700 28654
rect 7644 28550 7700 28588
rect 8876 28644 8932 29372
rect 9548 29428 9604 29438
rect 9548 29334 9604 29372
rect 10108 29428 10164 29438
rect 10780 29428 10836 30940
rect 11452 29652 11508 30942
rect 14364 30996 14420 31164
rect 14476 31218 14532 31724
rect 14476 31166 14478 31218
rect 14530 31166 14532 31218
rect 14476 31154 14532 31166
rect 14812 31218 14868 32620
rect 14924 32582 14980 32620
rect 15596 32676 15652 32686
rect 15596 32582 15652 32620
rect 16156 32676 16212 32686
rect 16156 32582 16212 32620
rect 17500 32676 17556 32686
rect 15036 32564 15092 32574
rect 15484 32564 15540 32574
rect 15036 32562 15540 32564
rect 15036 32510 15038 32562
rect 15090 32510 15486 32562
rect 15538 32510 15540 32562
rect 15036 32508 15540 32510
rect 15036 31948 15092 32508
rect 15484 32498 15540 32508
rect 15820 32562 15876 32574
rect 15820 32510 15822 32562
rect 15874 32510 15876 32562
rect 14812 31166 14814 31218
rect 14866 31166 14868 31218
rect 14812 31154 14868 31166
rect 14924 31892 15092 31948
rect 15820 31948 15876 32510
rect 16268 32562 16324 32574
rect 16268 32510 16270 32562
rect 16322 32510 16324 32562
rect 15820 31892 16212 31948
rect 14924 31106 14980 31892
rect 15036 31826 15092 31836
rect 16156 31778 16212 31892
rect 16268 31892 16324 32510
rect 17164 32340 17220 32350
rect 16324 31836 16436 31892
rect 16268 31826 16324 31836
rect 16156 31726 16158 31778
rect 16210 31726 16212 31778
rect 16156 31714 16212 31726
rect 16380 31218 16436 31836
rect 17164 31890 17220 32284
rect 17164 31838 17166 31890
rect 17218 31838 17220 31890
rect 17164 31826 17220 31838
rect 17500 31666 17556 32620
rect 17500 31614 17502 31666
rect 17554 31614 17556 31666
rect 17500 31602 17556 31614
rect 17836 31556 17892 35644
rect 17948 35634 18004 35644
rect 18284 35810 18340 35822
rect 18284 35758 18286 35810
rect 18338 35758 18340 35810
rect 18284 35252 18340 35758
rect 18620 35812 18676 35822
rect 18620 35718 18676 35756
rect 18732 35588 18788 35868
rect 19404 35858 19460 35868
rect 19292 35810 19348 35822
rect 19292 35758 19294 35810
rect 19346 35758 19348 35810
rect 18284 34804 18340 35196
rect 18284 34738 18340 34748
rect 18620 35532 18788 35588
rect 18844 35700 18900 35710
rect 19292 35700 19348 35758
rect 23548 35812 23604 35822
rect 23548 35718 23604 35756
rect 18844 35698 19348 35700
rect 18844 35646 18846 35698
rect 18898 35646 19348 35698
rect 18844 35644 19348 35646
rect 19516 35698 19572 35710
rect 19516 35646 19518 35698
rect 19570 35646 19572 35698
rect 17948 34692 18004 34702
rect 17948 34130 18004 34636
rect 17948 34078 17950 34130
rect 18002 34078 18004 34130
rect 17948 34066 18004 34078
rect 18620 34132 18676 35532
rect 18620 34066 18676 34076
rect 18732 34804 18788 34814
rect 18172 34020 18228 34030
rect 17948 33348 18004 33358
rect 17948 32786 18004 33292
rect 18172 33346 18228 33964
rect 18172 33294 18174 33346
rect 18226 33294 18228 33346
rect 18172 33282 18228 33294
rect 18620 33348 18676 33358
rect 18620 33254 18676 33292
rect 18732 33234 18788 34748
rect 18844 34356 18900 35644
rect 18844 34290 18900 34300
rect 18956 34914 19012 34926
rect 18956 34862 18958 34914
rect 19010 34862 19012 34914
rect 18956 33346 19012 34862
rect 18956 33294 18958 33346
rect 19010 33294 19012 33346
rect 18956 33282 19012 33294
rect 18732 33182 18734 33234
rect 18786 33182 18788 33234
rect 18732 33170 18788 33182
rect 17948 32734 17950 32786
rect 18002 32734 18004 32786
rect 17948 32722 18004 32734
rect 18284 32562 18340 32574
rect 18284 32510 18286 32562
rect 18338 32510 18340 32562
rect 18284 31948 18340 32510
rect 19516 31948 19572 35646
rect 20300 35700 20356 35710
rect 23660 35700 23716 36204
rect 24220 36036 24276 36046
rect 23772 35700 23828 35710
rect 20300 35698 20916 35700
rect 20300 35646 20302 35698
rect 20354 35646 20916 35698
rect 20300 35644 20916 35646
rect 23660 35644 23772 35700
rect 19964 34692 20020 34730
rect 19964 34626 20020 34636
rect 20188 34690 20244 34702
rect 20188 34638 20190 34690
rect 20242 34638 20244 34690
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20188 34354 20244 34638
rect 20188 34302 20190 34354
rect 20242 34302 20244 34354
rect 20188 34290 20244 34302
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 18284 31892 18452 31948
rect 17836 31462 17892 31500
rect 18284 31556 18340 31566
rect 18284 31462 18340 31500
rect 16380 31166 16382 31218
rect 16434 31166 16436 31218
rect 16380 31154 16436 31166
rect 14924 31054 14926 31106
rect 14978 31054 14980 31106
rect 14924 31042 14980 31054
rect 14588 30996 14644 31006
rect 14364 30994 14644 30996
rect 14364 30942 14590 30994
rect 14642 30942 14644 30994
rect 14364 30940 14644 30942
rect 14588 30930 14644 30940
rect 16716 30996 16772 31006
rect 16716 30902 16772 30940
rect 18396 30996 18452 31892
rect 15148 30324 15204 30334
rect 13804 30212 13860 30222
rect 14252 30212 14308 30222
rect 13804 30210 13972 30212
rect 13804 30158 13806 30210
rect 13858 30158 13972 30210
rect 13804 30156 13972 30158
rect 13804 30146 13860 30156
rect 11452 29586 11508 29596
rect 13244 29652 13300 29662
rect 13244 29558 13300 29596
rect 10108 29426 10500 29428
rect 10108 29374 10110 29426
rect 10162 29374 10500 29426
rect 10108 29372 10500 29374
rect 10108 29362 10164 29372
rect 10444 28754 10500 29372
rect 10780 29362 10836 29372
rect 12236 29426 12292 29438
rect 12236 29374 12238 29426
rect 12290 29374 12292 29426
rect 10444 28702 10446 28754
rect 10498 28702 10500 28754
rect 10444 28690 10500 28702
rect 8876 28578 8932 28588
rect 11116 27972 11172 27982
rect 12236 27972 12292 29374
rect 13020 29316 13076 29326
rect 13020 28082 13076 29260
rect 13916 29316 13972 30156
rect 14252 30210 15092 30212
rect 14252 30158 14254 30210
rect 14306 30158 15092 30210
rect 14252 30156 15092 30158
rect 14252 30146 14308 30156
rect 15036 29650 15092 30156
rect 15036 29598 15038 29650
rect 15090 29598 15092 29650
rect 15036 29586 15092 29598
rect 15148 29538 15204 30268
rect 15148 29486 15150 29538
rect 15202 29486 15204 29538
rect 15148 29474 15204 29486
rect 15932 30324 15988 30334
rect 13916 29222 13972 29260
rect 14028 29202 14084 29214
rect 14028 29150 14030 29202
rect 14082 29150 14084 29202
rect 14028 28532 14084 29150
rect 15932 28642 15988 30268
rect 17052 30324 17108 30334
rect 17052 30230 17108 30268
rect 17836 30212 17892 30222
rect 17612 30156 17836 30212
rect 16492 29986 16548 29998
rect 16492 29934 16494 29986
rect 16546 29934 16548 29986
rect 16380 29652 16436 29662
rect 16492 29652 16548 29934
rect 16380 29650 16548 29652
rect 16380 29598 16382 29650
rect 16434 29598 16548 29650
rect 16380 29596 16548 29598
rect 16380 29586 16436 29596
rect 16268 29540 16324 29550
rect 16268 29446 16324 29484
rect 17500 29540 17556 29550
rect 16828 29316 16884 29326
rect 16828 29222 16884 29260
rect 16716 29204 16772 29214
rect 15932 28590 15934 28642
rect 15986 28590 15988 28642
rect 15932 28578 15988 28590
rect 16380 29202 16772 29204
rect 16380 29150 16718 29202
rect 16770 29150 16772 29202
rect 16380 29148 16772 29150
rect 16380 28642 16436 29148
rect 16716 29138 16772 29148
rect 16380 28590 16382 28642
rect 16434 28590 16436 28642
rect 16380 28578 16436 28590
rect 14028 28466 14084 28476
rect 16044 28532 16100 28542
rect 13020 28030 13022 28082
rect 13074 28030 13076 28082
rect 13020 28018 13076 28030
rect 11004 27916 11116 27972
rect 11172 27916 11284 27972
rect 11004 27858 11060 27916
rect 11116 27906 11172 27916
rect 11004 27806 11006 27858
rect 11058 27806 11060 27858
rect 11004 27794 11060 27806
rect 11116 27746 11172 27758
rect 11116 27694 11118 27746
rect 11170 27694 11172 27746
rect 10780 27636 10836 27646
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 8540 27300 8596 27310
rect 8540 26292 8596 27244
rect 9212 27300 9268 27310
rect 8988 27188 9044 27198
rect 8316 26290 8596 26292
rect 8316 26238 8542 26290
rect 8594 26238 8596 26290
rect 8316 26236 8596 26238
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 8316 25620 8372 26236
rect 8540 26226 8596 26236
rect 8764 27076 8820 27086
rect 7868 25618 8372 25620
rect 7868 25566 8318 25618
rect 8370 25566 8372 25618
rect 7868 25564 8372 25566
rect 7308 25506 7364 25518
rect 7868 25508 7924 25564
rect 8316 25554 8372 25564
rect 7308 25454 7310 25506
rect 7362 25454 7364 25506
rect 6972 25284 7028 25294
rect 6972 24946 7028 25228
rect 6972 24894 6974 24946
rect 7026 24894 7028 24946
rect 6972 24882 7028 24894
rect 7196 24610 7252 24622
rect 7196 24558 7198 24610
rect 7250 24558 7252 24610
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 7196 24164 7252 24558
rect 6860 24108 7196 24164
rect 6188 23714 6244 23726
rect 6188 23662 6190 23714
rect 6242 23662 6244 23714
rect 6076 23154 6132 23166
rect 6076 23102 6078 23154
rect 6130 23102 6132 23154
rect 5516 23042 5572 23054
rect 5516 22990 5518 23042
rect 5570 22990 5572 23042
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4844 22372 4900 22382
rect 4844 22278 4900 22316
rect 5516 22372 5572 22990
rect 6076 23044 6132 23102
rect 6188 23156 6244 23662
rect 6524 23714 6580 23726
rect 6524 23662 6526 23714
rect 6578 23662 6580 23714
rect 6412 23156 6468 23166
rect 6188 23100 6412 23156
rect 6412 23062 6468 23100
rect 5516 22306 5572 22316
rect 5964 22370 6020 22382
rect 5964 22318 5966 22370
rect 6018 22318 6020 22370
rect 5068 22146 5124 22158
rect 5068 22094 5070 22146
rect 5122 22094 5124 22146
rect 5068 21700 5124 22094
rect 5292 21700 5348 21710
rect 5068 21644 5292 21700
rect 5292 21634 5348 21644
rect 3948 21588 4004 21598
rect 4396 21588 4452 21598
rect 3948 21586 4340 21588
rect 3948 21534 3950 21586
rect 4002 21534 4340 21586
rect 3948 21532 4340 21534
rect 3948 21522 4004 21532
rect 4284 20916 4340 21532
rect 4396 21494 4452 21532
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4396 20916 4452 20926
rect 4284 20914 4452 20916
rect 4284 20862 4398 20914
rect 4450 20862 4452 20914
rect 4284 20860 4452 20862
rect 4284 20578 4340 20590
rect 4284 20526 4286 20578
rect 4338 20526 4340 20578
rect 2044 20018 2100 20030
rect 2044 19966 2046 20018
rect 2098 19966 2100 20018
rect 2044 19124 2100 19966
rect 2604 20018 2660 20030
rect 2604 19966 2606 20018
rect 2658 19966 2660 20018
rect 2604 19908 2660 19966
rect 2604 19842 2660 19852
rect 4284 19908 4340 20526
rect 4396 20132 4452 20860
rect 5964 20914 6020 22318
rect 5964 20862 5966 20914
rect 6018 20862 6020 20914
rect 5068 20692 5124 20702
rect 5628 20692 5684 20702
rect 5068 20690 5684 20692
rect 5068 20638 5070 20690
rect 5122 20638 5630 20690
rect 5682 20638 5684 20690
rect 5068 20636 5684 20638
rect 5068 20626 5124 20636
rect 5628 20626 5684 20636
rect 4732 20580 4788 20590
rect 4732 20578 4900 20580
rect 4732 20526 4734 20578
rect 4786 20526 4900 20578
rect 4732 20524 4900 20526
rect 4732 20514 4788 20524
rect 4844 20242 4900 20524
rect 4844 20190 4846 20242
rect 4898 20190 4900 20242
rect 4844 20178 4900 20190
rect 5964 20188 6020 20862
rect 6076 20802 6132 22988
rect 6524 22484 6580 23662
rect 6524 22370 6580 22428
rect 6524 22318 6526 22370
rect 6578 22318 6580 22370
rect 6524 22306 6580 22318
rect 6636 21700 6692 21710
rect 6636 21606 6692 21644
rect 6076 20750 6078 20802
rect 6130 20750 6132 20802
rect 6076 20738 6132 20750
rect 4396 20066 4452 20076
rect 5628 20132 5684 20142
rect 5964 20132 6132 20188
rect 5628 20038 5684 20076
rect 4956 20020 5012 20030
rect 4284 19842 4340 19852
rect 4844 19964 4956 20020
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 3276 19236 3332 19246
rect 3276 19142 3332 19180
rect 4620 19234 4676 19246
rect 4620 19182 4622 19234
rect 4674 19182 4676 19234
rect 1596 18676 1652 18686
rect 2044 18676 2100 19068
rect 3164 19124 3220 19134
rect 3164 19030 3220 19068
rect 4620 19124 4676 19182
rect 4620 19058 4676 19068
rect 4844 19236 4900 19964
rect 4956 19954 5012 19964
rect 1596 18674 2100 18676
rect 1596 18622 1598 18674
rect 1650 18622 2100 18674
rect 1596 18620 2100 18622
rect 2380 18676 2436 18686
rect 1596 18610 1652 18620
rect 2380 18582 2436 18620
rect 4732 18452 4788 18462
rect 4844 18452 4900 19180
rect 4956 19348 5012 19358
rect 4956 19234 5012 19292
rect 6076 19348 6132 20132
rect 6076 19282 6132 19292
rect 6524 19348 6580 19358
rect 4956 19182 4958 19234
rect 5010 19182 5012 19234
rect 4956 19170 5012 19182
rect 5068 19236 5124 19246
rect 5068 19142 5124 19180
rect 5964 19236 6020 19246
rect 5964 19142 6020 19180
rect 5628 19010 5684 19022
rect 5628 18958 5630 19010
rect 5682 18958 5684 19010
rect 5628 18676 5684 18958
rect 5628 18610 5684 18620
rect 4732 18450 4900 18452
rect 4732 18398 4734 18450
rect 4786 18398 4900 18450
rect 4732 18396 4900 18398
rect 5180 18450 5236 18462
rect 5180 18398 5182 18450
rect 5234 18398 5236 18450
rect 4732 18386 4788 18396
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 5180 17780 5236 18398
rect 6412 18340 6468 18350
rect 6524 18340 6580 19292
rect 6860 19236 6916 24108
rect 7196 24098 7252 24108
rect 7196 23940 7252 23950
rect 7308 23940 7364 25454
rect 7756 25506 7924 25508
rect 7756 25454 7870 25506
rect 7922 25454 7924 25506
rect 7756 25452 7924 25454
rect 7756 25284 7812 25452
rect 7868 25442 7924 25452
rect 7756 24946 7812 25228
rect 7756 24894 7758 24946
rect 7810 24894 7812 24946
rect 7756 24882 7812 24894
rect 8092 24724 8148 24734
rect 7196 23938 7364 23940
rect 7196 23886 7198 23938
rect 7250 23886 7364 23938
rect 7196 23884 7364 23886
rect 7756 24722 8148 24724
rect 7756 24670 8094 24722
rect 8146 24670 8148 24722
rect 7756 24668 8148 24670
rect 7756 23938 7812 24668
rect 8092 24658 8148 24668
rect 8652 24612 8708 24622
rect 8764 24612 8820 27020
rect 8988 26290 9044 27132
rect 9212 27186 9268 27244
rect 9212 27134 9214 27186
rect 9266 27134 9268 27186
rect 9212 27122 9268 27134
rect 10108 27188 10164 27198
rect 9660 27076 9716 27086
rect 9660 26982 9716 27020
rect 10108 27074 10164 27132
rect 10108 27022 10110 27074
rect 10162 27022 10164 27074
rect 10108 27010 10164 27022
rect 10220 26964 10276 26974
rect 10108 26292 10164 26302
rect 8988 26238 8990 26290
rect 9042 26238 9044 26290
rect 8988 26226 9044 26238
rect 9660 26290 10164 26292
rect 9660 26238 10110 26290
rect 10162 26238 10164 26290
rect 9660 26236 10164 26238
rect 9660 26180 9716 26236
rect 10108 26226 10164 26236
rect 9548 26178 9716 26180
rect 9548 26126 9662 26178
rect 9714 26126 9716 26178
rect 9548 26124 9716 26126
rect 9548 25618 9604 26124
rect 9660 26114 9716 26124
rect 9772 26068 9828 26078
rect 9772 25974 9828 26012
rect 9548 25566 9550 25618
rect 9602 25566 9604 25618
rect 9548 25554 9604 25566
rect 10108 25396 10164 25406
rect 10220 25396 10276 26908
rect 10556 26962 10612 26974
rect 10556 26910 10558 26962
rect 10610 26910 10612 26962
rect 10556 26404 10612 26910
rect 10556 26338 10612 26348
rect 10668 26292 10724 26302
rect 10780 26292 10836 27580
rect 11004 27076 11060 27086
rect 11116 27076 11172 27694
rect 11060 27020 11172 27076
rect 11228 27188 11284 27916
rect 12236 27906 12292 27916
rect 13804 27972 13860 27982
rect 13804 27878 13860 27916
rect 16044 27858 16100 28476
rect 17388 27972 17444 27982
rect 17388 27878 17444 27916
rect 17500 27970 17556 29484
rect 17500 27918 17502 27970
rect 17554 27918 17556 27970
rect 17500 27906 17556 27918
rect 16044 27806 16046 27858
rect 16098 27806 16100 27858
rect 16044 27794 16100 27806
rect 16604 27860 16660 27870
rect 16604 27858 16772 27860
rect 16604 27806 16606 27858
rect 16658 27806 16772 27858
rect 16604 27804 16772 27806
rect 16604 27794 16660 27804
rect 11564 27748 11620 27758
rect 11564 27654 11620 27692
rect 12012 27746 12068 27758
rect 12012 27694 12014 27746
rect 12066 27694 12068 27746
rect 11900 27636 11956 27646
rect 11900 27542 11956 27580
rect 12012 27188 12068 27694
rect 12460 27748 12516 27758
rect 12012 27132 12404 27188
rect 11228 27074 11284 27132
rect 11228 27022 11230 27074
rect 11282 27022 11284 27074
rect 11004 26982 11060 27020
rect 11228 27010 11284 27022
rect 11900 26964 11956 26974
rect 12236 26964 12292 26974
rect 11900 26962 12180 26964
rect 11900 26910 11902 26962
rect 11954 26910 12180 26962
rect 11900 26908 12180 26910
rect 11900 26898 11956 26908
rect 10668 26290 10836 26292
rect 10668 26238 10670 26290
rect 10722 26238 10836 26290
rect 10668 26236 10836 26238
rect 12124 26292 12180 26908
rect 12236 26870 12292 26908
rect 12348 26628 12404 27132
rect 12460 27074 12516 27692
rect 15820 27300 15876 27310
rect 15820 27298 16660 27300
rect 15820 27246 15822 27298
rect 15874 27246 16660 27298
rect 15820 27244 16660 27246
rect 15820 27234 15876 27244
rect 12460 27022 12462 27074
rect 12514 27022 12516 27074
rect 12460 27010 12516 27022
rect 16268 27074 16324 27086
rect 16268 27022 16270 27074
rect 16322 27022 16324 27074
rect 15372 26964 15428 26974
rect 15708 26964 15764 26974
rect 15372 26962 15708 26964
rect 15372 26910 15374 26962
rect 15426 26910 15708 26962
rect 15372 26908 15708 26910
rect 15372 26898 15428 26908
rect 15708 26870 15764 26908
rect 12348 26562 12404 26572
rect 13468 26628 13524 26638
rect 13132 26516 13188 26526
rect 13132 26422 13188 26460
rect 12124 26236 12516 26292
rect 10668 26226 10724 26236
rect 10108 25394 10276 25396
rect 10108 25342 10110 25394
rect 10162 25342 10276 25394
rect 10108 25340 10276 25342
rect 12348 26068 12404 26078
rect 12348 25506 12404 26012
rect 12348 25454 12350 25506
rect 12402 25454 12404 25506
rect 10108 25330 10164 25340
rect 10332 25284 10388 25294
rect 8652 24610 8820 24612
rect 8652 24558 8654 24610
rect 8706 24558 8820 24610
rect 8652 24556 8820 24558
rect 8652 24546 8708 24556
rect 8764 24050 8820 24556
rect 8764 23998 8766 24050
rect 8818 23998 8820 24050
rect 8764 23986 8820 23998
rect 9884 24948 9940 24958
rect 7756 23886 7758 23938
rect 7810 23886 7812 23938
rect 7196 23154 7252 23884
rect 7196 23102 7198 23154
rect 7250 23102 7252 23154
rect 7196 23044 7252 23102
rect 7756 23156 7812 23886
rect 8540 23940 8596 23950
rect 8540 23846 8596 23884
rect 7868 23828 7924 23838
rect 7868 23734 7924 23772
rect 9212 23826 9268 23838
rect 9212 23774 9214 23826
rect 9266 23774 9268 23826
rect 8652 23266 8708 23278
rect 8652 23214 8654 23266
rect 8706 23214 8708 23266
rect 7756 23062 7812 23100
rect 7868 23156 7924 23166
rect 8316 23156 8372 23166
rect 7868 23154 8372 23156
rect 7868 23102 7870 23154
rect 7922 23102 8318 23154
rect 8370 23102 8372 23154
rect 7868 23100 8372 23102
rect 7868 23090 7924 23100
rect 8316 23090 8372 23100
rect 7196 22978 7252 22988
rect 6972 22372 7028 22382
rect 7420 22372 7476 22382
rect 6972 22370 7252 22372
rect 6972 22318 6974 22370
rect 7026 22318 7252 22370
rect 6972 22316 7252 22318
rect 6972 22306 7028 22316
rect 7196 21700 7252 22316
rect 7420 22278 7476 22316
rect 8652 22260 8708 23214
rect 9212 23044 9268 23774
rect 9548 23828 9604 23838
rect 9548 23734 9604 23772
rect 9884 23826 9940 24892
rect 10332 24946 10388 25228
rect 11676 25284 11732 25294
rect 10332 24894 10334 24946
rect 10386 24894 10388 24946
rect 10332 24882 10388 24894
rect 10892 24948 10948 24958
rect 10892 24854 10948 24892
rect 9884 23774 9886 23826
rect 9938 23774 9940 23826
rect 9884 23762 9940 23774
rect 9212 22978 9268 22988
rect 10780 23154 10836 23166
rect 11228 23156 11284 23166
rect 10780 23102 10782 23154
rect 10834 23102 10836 23154
rect 10444 22596 10500 22606
rect 10500 22540 10612 22596
rect 10444 22502 10500 22540
rect 10444 22372 10500 22382
rect 9660 22260 9716 22270
rect 8652 22258 9716 22260
rect 8652 22206 9662 22258
rect 9714 22206 9716 22258
rect 8652 22204 9716 22206
rect 9660 22194 9716 22204
rect 9212 21924 9268 21934
rect 7644 21700 7700 21710
rect 7196 21698 7700 21700
rect 7196 21646 7646 21698
rect 7698 21646 7700 21698
rect 7196 21644 7700 21646
rect 7196 21474 7252 21644
rect 7644 21634 7700 21644
rect 7756 21588 7812 21598
rect 7756 21494 7812 21532
rect 7196 21422 7198 21474
rect 7250 21422 7252 21474
rect 7196 21410 7252 21422
rect 9212 20690 9268 21868
rect 9212 20638 9214 20690
rect 9266 20638 9268 20690
rect 9212 20626 9268 20638
rect 10444 21362 10500 22316
rect 10556 21698 10612 22540
rect 10668 22146 10724 22158
rect 10668 22094 10670 22146
rect 10722 22094 10724 22146
rect 10668 21924 10724 22094
rect 10780 22148 10836 23102
rect 11116 23154 11284 23156
rect 11116 23102 11230 23154
rect 11282 23102 11284 23154
rect 11116 23100 11284 23102
rect 10892 23044 10948 23054
rect 10892 22370 10948 22988
rect 10892 22318 10894 22370
rect 10946 22318 10948 22370
rect 10892 22306 10948 22318
rect 10892 22148 10948 22158
rect 10780 22092 10892 22148
rect 10892 22082 10948 22092
rect 10668 21858 10724 21868
rect 10556 21646 10558 21698
rect 10610 21646 10612 21698
rect 10556 21634 10612 21646
rect 11004 21812 11060 21822
rect 11116 21812 11172 23100
rect 11228 23090 11284 23100
rect 11004 21810 11172 21812
rect 11004 21758 11006 21810
rect 11058 21758 11172 21810
rect 11004 21756 11172 21758
rect 11340 22372 11396 22382
rect 10444 21310 10446 21362
rect 10498 21310 10500 21362
rect 8428 20578 8484 20590
rect 8428 20526 8430 20578
rect 8482 20526 8484 20578
rect 8428 20132 8484 20526
rect 10444 20580 10500 21310
rect 10892 21474 10948 21486
rect 10892 21422 10894 21474
rect 10946 21422 10948 21474
rect 10892 21364 10948 21422
rect 10892 21298 10948 21308
rect 10444 20514 10500 20524
rect 8428 20066 8484 20076
rect 6636 19234 6916 19236
rect 6636 19182 6862 19234
rect 6914 19182 6916 19234
rect 6636 19180 6916 19182
rect 6636 19124 6692 19180
rect 6860 19170 6916 19180
rect 11004 19236 11060 21756
rect 11340 21586 11396 22316
rect 11676 22258 11732 25228
rect 11900 22708 11956 22718
rect 11788 22652 11900 22708
rect 11788 22594 11844 22652
rect 11900 22642 11956 22652
rect 11788 22542 11790 22594
rect 11842 22542 11844 22594
rect 11788 22530 11844 22542
rect 12348 22372 12404 25454
rect 12460 23938 12516 26236
rect 13468 26178 13524 26572
rect 13916 26516 13972 26526
rect 13916 26422 13972 26460
rect 14140 26404 14196 26414
rect 14140 26290 14196 26348
rect 14140 26238 14142 26290
rect 14194 26238 14196 26290
rect 14140 26226 14196 26238
rect 13468 26126 13470 26178
rect 13522 26126 13524 26178
rect 12796 25506 12852 25518
rect 12796 25454 12798 25506
rect 12850 25454 12852 25506
rect 12796 25284 12852 25454
rect 12796 25218 12852 25228
rect 13356 24724 13412 24734
rect 12460 23886 12462 23938
rect 12514 23886 12516 23938
rect 12460 23874 12516 23886
rect 12684 24722 13412 24724
rect 12684 24670 13358 24722
rect 13410 24670 13412 24722
rect 12684 24668 13412 24670
rect 12684 22708 12740 24668
rect 13356 24658 13412 24668
rect 13468 24500 13524 26126
rect 16268 25732 16324 27022
rect 16604 27074 16660 27244
rect 16604 27022 16606 27074
rect 16658 27022 16660 27074
rect 16604 27010 16660 27022
rect 16716 26964 16772 27804
rect 16772 26908 16884 26964
rect 16716 26870 16772 26908
rect 16828 26292 16884 26908
rect 16828 26198 16884 26236
rect 17500 26178 17556 26190
rect 17500 26126 17502 26178
rect 17554 26126 17556 26178
rect 16268 25666 16324 25676
rect 16716 26068 16772 26078
rect 16156 25508 16212 25518
rect 15708 25506 16212 25508
rect 15708 25454 16158 25506
rect 16210 25454 16212 25506
rect 15708 25452 16212 25454
rect 15708 25394 15764 25452
rect 16156 25442 16212 25452
rect 16716 25506 16772 26012
rect 17388 26068 17444 26078
rect 17388 25974 17444 26012
rect 17500 25732 17556 26126
rect 17500 25666 17556 25676
rect 16716 25454 16718 25506
rect 16770 25454 16772 25506
rect 16716 25442 16772 25454
rect 15708 25342 15710 25394
rect 15762 25342 15764 25394
rect 13804 24724 13860 24734
rect 13244 24444 13524 24500
rect 13692 24722 13860 24724
rect 13692 24670 13806 24722
rect 13858 24670 13860 24722
rect 13692 24668 13860 24670
rect 12796 23714 12852 23726
rect 12796 23662 12798 23714
rect 12850 23662 12852 23714
rect 12796 23380 12852 23662
rect 12796 23314 12852 23324
rect 12348 22278 12404 22316
rect 12572 22372 12628 22382
rect 11676 22206 11678 22258
rect 11730 22206 11732 22258
rect 11340 21534 11342 21586
rect 11394 21534 11396 21586
rect 11340 21522 11396 21534
rect 11564 21812 11620 21822
rect 11564 21586 11620 21756
rect 11676 21700 11732 22206
rect 12460 22260 12516 22270
rect 12572 22260 12628 22316
rect 12684 22370 12740 22652
rect 12796 22484 12852 22494
rect 12796 22482 12964 22484
rect 12796 22430 12798 22482
rect 12850 22430 12964 22482
rect 12796 22428 12964 22430
rect 12796 22418 12852 22428
rect 12684 22318 12686 22370
rect 12738 22318 12740 22370
rect 12684 22306 12740 22318
rect 12460 22258 12628 22260
rect 12460 22206 12462 22258
rect 12514 22206 12628 22258
rect 12460 22204 12628 22206
rect 12796 22260 12852 22270
rect 12460 21812 12516 22204
rect 12796 22166 12852 22204
rect 12460 21746 12516 21756
rect 12908 21810 12964 22428
rect 12908 21758 12910 21810
rect 12962 21758 12964 21810
rect 12908 21746 12964 21758
rect 13244 22148 13300 24444
rect 13580 23380 13636 23390
rect 13580 23286 13636 23324
rect 13692 22596 13748 24668
rect 13804 24658 13860 24668
rect 15484 24052 15540 24062
rect 15708 24052 15764 25342
rect 15820 25282 15876 25294
rect 15820 25230 15822 25282
rect 15874 25230 15876 25282
rect 15820 24500 15876 25230
rect 15820 24434 15876 24444
rect 16044 25284 16100 25294
rect 15484 24050 15764 24052
rect 15484 23998 15486 24050
rect 15538 23998 15764 24050
rect 15484 23996 15764 23998
rect 15484 23986 15540 23996
rect 16044 23826 16100 25228
rect 16044 23774 16046 23826
rect 16098 23774 16100 23826
rect 16044 23762 16100 23774
rect 13580 22372 13636 22382
rect 13692 22372 13748 22540
rect 13580 22370 13748 22372
rect 13580 22318 13582 22370
rect 13634 22318 13748 22370
rect 13580 22316 13748 22318
rect 14140 23042 14196 23054
rect 14140 22990 14142 23042
rect 14194 22990 14196 23042
rect 13580 22306 13636 22316
rect 11676 21634 11732 21644
rect 11564 21534 11566 21586
rect 11618 21534 11620 21586
rect 11564 21522 11620 21534
rect 11788 21588 11844 21598
rect 11788 21494 11844 21532
rect 12012 21588 12068 21598
rect 12012 21586 12180 21588
rect 12012 21534 12014 21586
rect 12066 21534 12180 21586
rect 12012 21532 12180 21534
rect 12012 21522 12068 21532
rect 11900 21474 11956 21486
rect 11900 21422 11902 21474
rect 11954 21422 11956 21474
rect 11900 21028 11956 21422
rect 11788 20972 11956 21028
rect 12012 21364 12068 21374
rect 11564 20916 11620 20926
rect 11564 20804 11620 20860
rect 11452 20802 11620 20804
rect 11452 20750 11566 20802
rect 11618 20750 11620 20802
rect 11452 20748 11620 20750
rect 11452 20242 11508 20748
rect 11564 20738 11620 20748
rect 11452 20190 11454 20242
rect 11506 20190 11508 20242
rect 11452 20178 11508 20190
rect 11788 20188 11844 20972
rect 12012 20802 12068 21308
rect 12012 20750 12014 20802
rect 12066 20750 12068 20802
rect 12012 20738 12068 20750
rect 12124 20804 12180 21532
rect 13132 21586 13188 21598
rect 13132 21534 13134 21586
rect 13186 21534 13188 21586
rect 12348 21476 12404 21486
rect 12236 20804 12292 20814
rect 12124 20748 12236 20804
rect 12236 20738 12292 20748
rect 11340 20132 11396 20142
rect 11004 19170 11060 19180
rect 11116 19908 11172 19918
rect 6636 18450 6692 19068
rect 7420 19124 7476 19134
rect 7420 19122 7924 19124
rect 7420 19070 7422 19122
rect 7474 19070 7924 19122
rect 7420 19068 7924 19070
rect 7420 19058 7476 19068
rect 7644 18562 7700 18574
rect 7644 18510 7646 18562
rect 7698 18510 7700 18562
rect 6636 18398 6638 18450
rect 6690 18398 6692 18450
rect 6636 18386 6692 18398
rect 7196 18452 7252 18462
rect 7196 18358 7252 18396
rect 6412 18338 6580 18340
rect 6412 18286 6414 18338
rect 6466 18286 6580 18338
rect 6412 18284 6580 18286
rect 6412 18274 6468 18284
rect 5180 17714 5236 17724
rect 5964 17780 6020 17790
rect 5964 17686 6020 17724
rect 6524 17556 6580 17566
rect 6524 17462 6580 17500
rect 7644 17556 7700 18510
rect 7868 18450 7924 19068
rect 11116 19012 11172 19852
rect 11340 19124 11396 20076
rect 11676 20132 11844 20188
rect 11340 19068 11620 19124
rect 7868 18398 7870 18450
rect 7922 18398 7924 18450
rect 7868 18386 7924 18398
rect 8316 18562 8372 18574
rect 8316 18510 8318 18562
rect 8370 18510 8372 18562
rect 8316 17780 8372 18510
rect 8876 18564 8932 18574
rect 8540 18452 8596 18462
rect 8540 18358 8596 18396
rect 7644 17490 7700 17500
rect 8204 17724 8372 17780
rect 6076 17108 6132 17118
rect 6076 17014 6132 17052
rect 8204 17108 8260 17724
rect 8876 17666 8932 18508
rect 9772 18564 9828 18574
rect 10444 18564 10500 18574
rect 9772 17890 9828 18508
rect 9772 17838 9774 17890
rect 9826 17838 9828 17890
rect 9772 17826 9828 17838
rect 10220 18562 10500 18564
rect 10220 18510 10446 18562
rect 10498 18510 10500 18562
rect 10220 18508 10500 18510
rect 9660 17780 9716 17790
rect 8876 17614 8878 17666
rect 8930 17614 8932 17666
rect 8876 17602 8932 17614
rect 9324 17666 9380 17678
rect 9324 17614 9326 17666
rect 9378 17614 9380 17666
rect 8204 17042 8260 17052
rect 8988 17108 9044 17118
rect 7196 16996 7252 17006
rect 5292 16884 5348 16894
rect 5292 16790 5348 16828
rect 7084 16884 7140 16894
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 7084 16210 7140 16828
rect 7196 16322 7252 16940
rect 8316 16996 8372 17006
rect 8316 16882 8372 16940
rect 8316 16830 8318 16882
rect 8370 16830 8372 16882
rect 8316 16818 8372 16830
rect 8988 16884 9044 17052
rect 9324 16884 9380 17614
rect 8988 16882 9156 16884
rect 8988 16830 8990 16882
rect 9042 16830 9156 16882
rect 8988 16828 9156 16830
rect 8988 16818 9044 16828
rect 7196 16270 7198 16322
rect 7250 16270 7252 16322
rect 7196 16258 7252 16270
rect 9100 16212 9156 16828
rect 9324 16818 9380 16828
rect 9660 16324 9716 17724
rect 10108 17442 10164 17454
rect 10108 17390 10110 17442
rect 10162 17390 10164 17442
rect 9996 16884 10052 16894
rect 10108 16884 10164 17390
rect 9996 16882 10164 16884
rect 9996 16830 9998 16882
rect 10050 16830 10164 16882
rect 9996 16828 10164 16830
rect 9884 16324 9940 16334
rect 9660 16322 9940 16324
rect 9660 16270 9886 16322
rect 9938 16270 9940 16322
rect 9660 16268 9940 16270
rect 9884 16258 9940 16268
rect 7084 16158 7086 16210
rect 7138 16158 7140 16210
rect 7084 16146 7140 16158
rect 8652 16210 9156 16212
rect 8652 16158 9102 16210
rect 9154 16158 9156 16210
rect 8652 16156 9156 16158
rect 8428 15316 8484 15326
rect 8428 15222 8484 15260
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 8652 8428 8708 16156
rect 9100 16146 9156 16156
rect 9548 15988 9604 15998
rect 9548 15894 9604 15932
rect 8764 15876 8820 15886
rect 8764 15538 8820 15820
rect 9436 15876 9492 15886
rect 9436 15782 9492 15820
rect 8764 15486 8766 15538
rect 8818 15486 8820 15538
rect 8764 15474 8820 15486
rect 8988 15428 9044 15438
rect 8988 15334 9044 15372
rect 8876 15314 8932 15326
rect 8876 15262 8878 15314
rect 8930 15262 8932 15314
rect 8876 14868 8932 15262
rect 9660 15316 9716 15326
rect 9996 15316 10052 16828
rect 10108 16098 10164 16110
rect 10108 16046 10110 16098
rect 10162 16046 10164 16098
rect 10108 15876 10164 16046
rect 10220 15988 10276 18508
rect 10444 18498 10500 18508
rect 10668 18564 10724 18574
rect 10668 18470 10724 18508
rect 10892 18452 10948 18462
rect 10892 18358 10948 18396
rect 11116 18450 11172 18956
rect 11116 18398 11118 18450
rect 11170 18398 11172 18450
rect 11116 18386 11172 18398
rect 10556 18340 10612 18350
rect 11452 18340 11508 18350
rect 10556 18246 10612 18284
rect 11340 18338 11508 18340
rect 11340 18286 11454 18338
rect 11506 18286 11508 18338
rect 11340 18284 11508 18286
rect 10332 17666 10388 17678
rect 10332 17614 10334 17666
rect 10386 17614 10388 17666
rect 10332 16996 10388 17614
rect 10332 16940 10612 16996
rect 10332 16772 10388 16782
rect 10332 16098 10388 16716
rect 10444 16660 10500 16670
rect 10444 16210 10500 16604
rect 10444 16158 10446 16210
rect 10498 16158 10500 16210
rect 10444 16146 10500 16158
rect 10332 16046 10334 16098
rect 10386 16046 10388 16098
rect 10332 16034 10388 16046
rect 10556 16100 10612 16940
rect 10668 16882 10724 16894
rect 10668 16830 10670 16882
rect 10722 16830 10724 16882
rect 10668 16772 10724 16830
rect 10668 16706 10724 16716
rect 11340 16660 11396 18284
rect 11452 18274 11508 18284
rect 11452 17892 11508 17902
rect 11564 17892 11620 19068
rect 11676 18450 11732 20132
rect 12348 20130 12404 21420
rect 12460 21362 12516 21374
rect 12460 21310 12462 21362
rect 12514 21310 12516 21362
rect 12460 20916 12516 21310
rect 12572 21364 12628 21374
rect 12572 21362 12852 21364
rect 12572 21310 12574 21362
rect 12626 21310 12852 21362
rect 12572 21308 12852 21310
rect 12572 21298 12628 21308
rect 12460 20850 12516 20860
rect 12572 21140 12628 21150
rect 12348 20078 12350 20130
rect 12402 20078 12404 20130
rect 12348 20066 12404 20078
rect 12572 20130 12628 21084
rect 12572 20078 12574 20130
rect 12626 20078 12628 20130
rect 12572 20066 12628 20078
rect 12684 20132 12740 20142
rect 12684 20038 12740 20076
rect 12012 20020 12068 20030
rect 12012 19926 12068 19964
rect 12124 20018 12180 20030
rect 12124 19966 12126 20018
rect 12178 19966 12180 20018
rect 12124 19348 12180 19966
rect 12236 19348 12292 19358
rect 12124 19346 12292 19348
rect 12124 19294 12238 19346
rect 12290 19294 12292 19346
rect 12124 19292 12292 19294
rect 12236 19282 12292 19292
rect 11900 19236 11956 19246
rect 11900 19142 11956 19180
rect 12124 19124 12180 19134
rect 12124 19030 12180 19068
rect 12348 19012 12404 19022
rect 12348 18918 12404 18956
rect 12460 19010 12516 19022
rect 12460 18958 12462 19010
rect 12514 18958 12516 19010
rect 11676 18398 11678 18450
rect 11730 18398 11732 18450
rect 11676 18386 11732 18398
rect 12460 18452 12516 18958
rect 11900 18340 11956 18350
rect 11900 18246 11956 18284
rect 11452 17890 11620 17892
rect 11452 17838 11454 17890
rect 11506 17838 11620 17890
rect 11452 17836 11620 17838
rect 12124 18226 12180 18238
rect 12124 18174 12126 18226
rect 12178 18174 12180 18226
rect 11452 17826 11508 17836
rect 11676 17780 11732 17790
rect 11676 17686 11732 17724
rect 12012 17780 12068 17790
rect 12124 17780 12180 18174
rect 12012 17778 12180 17780
rect 12012 17726 12014 17778
rect 12066 17726 12180 17778
rect 12012 17724 12180 17726
rect 12012 17714 12068 17724
rect 11900 17442 11956 17454
rect 11900 17390 11902 17442
rect 11954 17390 11956 17442
rect 11900 16996 11956 17390
rect 11900 16930 11956 16940
rect 12124 17442 12180 17454
rect 12124 17390 12126 17442
rect 12178 17390 12180 17442
rect 11340 16594 11396 16604
rect 11788 16884 11844 16894
rect 11228 16212 11284 16222
rect 11228 16118 11284 16156
rect 10556 16034 10612 16044
rect 10220 15922 10276 15932
rect 11788 15986 11844 16828
rect 12124 16212 12180 17390
rect 12460 16884 12516 18396
rect 12572 18676 12628 18686
rect 12572 18450 12628 18620
rect 12796 18564 12852 21308
rect 12908 20692 12964 20702
rect 12908 20130 12964 20636
rect 12908 20078 12910 20130
rect 12962 20078 12964 20130
rect 12908 20066 12964 20078
rect 13132 19572 13188 21534
rect 13244 20188 13300 22092
rect 13692 22146 13748 22158
rect 13692 22094 13694 22146
rect 13746 22094 13748 22146
rect 13692 21812 13748 22094
rect 13692 21746 13748 21756
rect 13804 22146 13860 22158
rect 13804 22094 13806 22146
rect 13858 22094 13860 22146
rect 13356 21586 13412 21598
rect 13356 21534 13358 21586
rect 13410 21534 13412 21586
rect 13356 21252 13412 21534
rect 13468 21476 13524 21486
rect 13468 21474 13748 21476
rect 13468 21422 13470 21474
rect 13522 21422 13748 21474
rect 13468 21420 13748 21422
rect 13468 21410 13524 21420
rect 13356 21196 13636 21252
rect 13468 20692 13524 20702
rect 13468 20598 13524 20636
rect 13244 20132 13412 20188
rect 13356 20018 13412 20132
rect 13356 19966 13358 20018
rect 13410 19966 13412 20018
rect 13356 19954 13412 19966
rect 13580 19908 13636 21196
rect 13692 21026 13748 21420
rect 13804 21140 13860 22094
rect 13916 22146 13972 22158
rect 13916 22094 13918 22146
rect 13970 22094 13972 22146
rect 13916 21588 13972 22094
rect 13916 21522 13972 21532
rect 14028 22146 14084 22158
rect 14028 22094 14030 22146
rect 14082 22094 14084 22146
rect 13804 21074 13860 21084
rect 13692 20974 13694 21026
rect 13746 20974 13748 21026
rect 13692 20962 13748 20974
rect 13916 20802 13972 20814
rect 13916 20750 13918 20802
rect 13970 20750 13972 20802
rect 13916 20132 13972 20750
rect 14028 20804 14084 22094
rect 14140 21586 14196 22990
rect 14588 23044 14644 23054
rect 14476 21700 14532 21710
rect 14476 21606 14532 21644
rect 14140 21534 14142 21586
rect 14194 21534 14196 21586
rect 14140 21364 14196 21534
rect 14140 21298 14196 21308
rect 14252 21586 14308 21598
rect 14252 21534 14254 21586
rect 14306 21534 14308 21586
rect 14028 20738 14084 20748
rect 14140 20802 14196 20814
rect 14140 20750 14142 20802
rect 14194 20750 14196 20802
rect 14140 20188 14196 20750
rect 14252 20804 14308 21534
rect 14364 21476 14420 21486
rect 14364 21382 14420 21420
rect 14252 20748 14532 20804
rect 13916 20066 13972 20076
rect 14028 20132 14196 20188
rect 14252 20580 14308 20590
rect 13580 19842 13636 19852
rect 13804 19906 13860 19918
rect 13804 19854 13806 19906
rect 13858 19854 13860 19906
rect 13804 19796 13860 19854
rect 13804 19730 13860 19740
rect 13132 19506 13188 19516
rect 14028 18676 14084 20132
rect 14252 20130 14308 20524
rect 14476 20468 14532 20748
rect 14588 20690 14644 22988
rect 15260 22482 15316 22494
rect 15260 22430 15262 22482
rect 15314 22430 15316 22482
rect 15260 22260 15316 22430
rect 15260 22194 15316 22204
rect 15820 22260 15876 22270
rect 15484 21812 15540 21822
rect 15484 21718 15540 21756
rect 14700 21700 14756 21710
rect 14700 21586 14756 21644
rect 15820 21698 15876 22204
rect 17388 22258 17444 22270
rect 17388 22206 17390 22258
rect 17442 22206 17444 22258
rect 16492 21812 16548 21822
rect 17388 21812 17444 22206
rect 17500 21812 17556 21822
rect 17388 21810 17556 21812
rect 17388 21758 17502 21810
rect 17554 21758 17556 21810
rect 17388 21756 17556 21758
rect 15820 21646 15822 21698
rect 15874 21646 15876 21698
rect 15820 21634 15876 21646
rect 15932 21700 15988 21710
rect 15932 21606 15988 21644
rect 16492 21698 16548 21756
rect 17500 21746 17556 21756
rect 16492 21646 16494 21698
rect 16546 21646 16548 21698
rect 16492 21634 16548 21646
rect 14700 21534 14702 21586
rect 14754 21534 14756 21586
rect 14700 21522 14756 21534
rect 16380 21588 16436 21598
rect 16380 21494 16436 21532
rect 16940 21588 16996 21598
rect 17276 21588 17332 21598
rect 16940 21586 17332 21588
rect 16940 21534 16942 21586
rect 16994 21534 17278 21586
rect 17330 21534 17332 21586
rect 16940 21532 17332 21534
rect 16940 21522 16996 21532
rect 14588 20638 14590 20690
rect 14642 20638 14644 20690
rect 14588 20626 14644 20638
rect 15372 21474 15428 21486
rect 15372 21422 15374 21474
rect 15426 21422 15428 21474
rect 15372 20914 15428 21422
rect 16716 21476 16772 21486
rect 16716 21382 16772 21420
rect 17276 21364 17332 21532
rect 17276 21298 17332 21308
rect 17500 21476 17556 21486
rect 15372 20862 15374 20914
rect 15426 20862 15428 20914
rect 14476 20412 15092 20468
rect 14476 20244 14532 20282
rect 14476 20178 14532 20188
rect 14252 20078 14254 20130
rect 14306 20078 14308 20130
rect 14252 20066 14308 20078
rect 14588 20020 14644 20030
rect 14588 19926 14644 19964
rect 14700 20018 14756 20030
rect 14700 19966 14702 20018
rect 14754 19966 14756 20018
rect 14140 19908 14196 19918
rect 14140 19346 14196 19852
rect 14700 19684 14756 19966
rect 14700 19618 14756 19628
rect 14812 20018 14868 20030
rect 14812 19966 14814 20018
rect 14866 19966 14868 20018
rect 14140 19294 14142 19346
rect 14194 19294 14196 19346
rect 14140 19124 14196 19294
rect 14140 19058 14196 19068
rect 14812 19572 14868 19966
rect 15036 19684 15092 20412
rect 15372 20244 15428 20862
rect 17500 20914 17556 21420
rect 17500 20862 17502 20914
rect 17554 20862 17556 20914
rect 17500 20850 17556 20862
rect 15372 20178 15428 20188
rect 17388 20692 17444 20702
rect 17612 20692 17668 30156
rect 17836 30118 17892 30156
rect 18284 29540 18340 29550
rect 18172 29484 18284 29540
rect 17836 29428 17892 29438
rect 17836 29334 17892 29372
rect 18172 27970 18228 29484
rect 18284 29446 18340 29484
rect 18396 29428 18452 30940
rect 19292 31892 19572 31948
rect 20188 32564 20244 32574
rect 20300 32564 20356 35644
rect 20412 34804 20468 34814
rect 20412 34710 20468 34748
rect 20524 34802 20580 34814
rect 20524 34750 20526 34802
rect 20578 34750 20580 34802
rect 20524 33348 20580 34750
rect 20860 34132 20916 35644
rect 23772 35634 23828 35644
rect 24108 35698 24164 35710
rect 24108 35646 24110 35698
rect 24162 35646 24164 35698
rect 20972 35586 21028 35598
rect 20972 35534 20974 35586
rect 21026 35534 21028 35586
rect 20972 34692 21028 35534
rect 23100 35586 23156 35598
rect 23100 35534 23102 35586
rect 23154 35534 23156 35586
rect 20972 34626 21028 34636
rect 21084 35476 21140 35486
rect 20972 34356 21028 34366
rect 21084 34356 21140 35420
rect 23100 35476 23156 35534
rect 23436 35476 23492 35486
rect 23100 35410 23156 35420
rect 23212 35474 23492 35476
rect 23212 35422 23438 35474
rect 23490 35422 23492 35474
rect 23212 35420 23492 35422
rect 21980 34916 22036 34926
rect 22540 34916 22596 34926
rect 23212 34916 23268 35420
rect 23436 35410 23492 35420
rect 21980 34914 22260 34916
rect 21980 34862 21982 34914
rect 22034 34862 22260 34914
rect 21980 34860 22260 34862
rect 21980 34850 22036 34860
rect 20972 34354 21084 34356
rect 20972 34302 20974 34354
rect 21026 34302 21084 34354
rect 20972 34300 21084 34302
rect 20972 34290 21028 34300
rect 21084 34262 21140 34300
rect 22092 34356 22148 34366
rect 21196 34132 21252 34142
rect 20860 34130 21252 34132
rect 20860 34078 21198 34130
rect 21250 34078 21252 34130
rect 20860 34076 21252 34078
rect 21196 34066 21252 34076
rect 21980 34132 22036 34142
rect 21980 34038 22036 34076
rect 22092 33458 22148 34300
rect 22092 33406 22094 33458
rect 22146 33406 22148 33458
rect 22092 33394 22148 33406
rect 20524 33282 20580 33292
rect 21308 33346 21364 33358
rect 21308 33294 21310 33346
rect 21362 33294 21364 33346
rect 20188 32562 20356 32564
rect 20188 32510 20190 32562
rect 20242 32510 20356 32562
rect 20188 32508 20356 32510
rect 18620 30772 18676 30782
rect 18620 30210 18676 30716
rect 18620 30158 18622 30210
rect 18674 30158 18676 30210
rect 18620 30146 18676 30158
rect 18396 29362 18452 29372
rect 19180 29316 19236 29326
rect 18396 29202 18452 29214
rect 18396 29150 18398 29202
rect 18450 29150 18452 29202
rect 18396 28532 18452 29150
rect 19180 28756 19236 29260
rect 18732 28754 19236 28756
rect 18732 28702 19182 28754
rect 19234 28702 19236 28754
rect 18732 28700 19236 28702
rect 18620 28532 18676 28542
rect 18396 28530 18676 28532
rect 18396 28478 18622 28530
rect 18674 28478 18676 28530
rect 18396 28476 18676 28478
rect 18620 28466 18676 28476
rect 18172 27918 18174 27970
rect 18226 27918 18228 27970
rect 18172 27906 18228 27918
rect 18732 27858 18788 28700
rect 19180 28690 19236 28700
rect 18732 27806 18734 27858
rect 18786 27806 18788 27858
rect 18732 27794 18788 27806
rect 19180 27860 19236 27870
rect 19180 27766 19236 27804
rect 18284 27634 18340 27646
rect 18284 27582 18286 27634
rect 18338 27582 18340 27634
rect 18284 26964 18340 27582
rect 18284 26898 18340 26908
rect 18956 26964 19012 26974
rect 19292 26908 19348 31892
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20076 31220 20132 31230
rect 20188 31220 20244 32508
rect 20860 32452 20916 32462
rect 20860 32358 20916 32396
rect 21308 31948 21364 33294
rect 20076 31218 20244 31220
rect 20076 31166 20078 31218
rect 20130 31166 20244 31218
rect 20076 31164 20244 31166
rect 20076 31154 20132 31164
rect 20188 31108 20244 31164
rect 20748 31892 21364 31948
rect 22204 33236 22260 34860
rect 22540 34914 23268 34916
rect 22540 34862 22542 34914
rect 22594 34862 23268 34914
rect 22540 34860 23268 34862
rect 22540 34850 22596 34860
rect 24108 34244 24164 35646
rect 24220 35698 24276 35980
rect 24668 35924 24724 35934
rect 24220 35646 24222 35698
rect 24274 35646 24276 35698
rect 24220 35140 24276 35646
rect 24444 35700 24500 35710
rect 24444 35606 24500 35644
rect 24668 35698 24724 35868
rect 24668 35646 24670 35698
rect 24722 35646 24724 35698
rect 24332 35588 24388 35598
rect 24332 35494 24388 35532
rect 24444 35252 24500 35262
rect 24220 35084 24388 35140
rect 24108 34018 24164 34188
rect 24108 33966 24110 34018
rect 24162 33966 24164 34018
rect 24108 33954 24164 33966
rect 24220 33458 24276 33470
rect 24220 33406 24222 33458
rect 24274 33406 24276 33458
rect 24220 33348 24276 33406
rect 24220 33282 24276 33292
rect 20524 31108 20580 31118
rect 20188 31106 20580 31108
rect 20188 31054 20526 31106
rect 20578 31054 20580 31106
rect 20188 31052 20580 31054
rect 20524 31042 20580 31052
rect 19852 30996 19908 31006
rect 19852 30902 19908 30940
rect 20748 30996 20804 31892
rect 20412 30772 20468 30782
rect 20412 30678 20468 30716
rect 20748 30322 20804 30940
rect 20748 30270 20750 30322
rect 20802 30270 20804 30322
rect 20748 30258 20804 30270
rect 20972 30882 21028 30894
rect 20972 30830 20974 30882
rect 21026 30830 21028 30882
rect 20972 30212 21028 30830
rect 21420 30884 21476 30894
rect 21420 30790 21476 30828
rect 22204 30884 22260 33180
rect 24332 32676 24388 35084
rect 24444 34242 24500 35196
rect 24556 34804 24612 34814
rect 24556 34354 24612 34748
rect 24556 34302 24558 34354
rect 24610 34302 24612 34354
rect 24556 34290 24612 34302
rect 24444 34190 24446 34242
rect 24498 34190 24500 34242
rect 24444 34178 24500 34190
rect 24668 33122 24724 35646
rect 25228 35700 25284 37102
rect 25340 37044 25396 37054
rect 25340 37042 25844 37044
rect 25340 36990 25342 37042
rect 25394 36990 25844 37042
rect 25340 36988 25844 36990
rect 25340 36978 25396 36988
rect 25788 36484 25844 36988
rect 25900 36484 25956 36494
rect 25788 36482 25956 36484
rect 25788 36430 25902 36482
rect 25954 36430 25956 36482
rect 25788 36428 25956 36430
rect 25900 36418 25956 36428
rect 26012 36260 26068 36270
rect 25452 35700 25508 35710
rect 25228 35644 25452 35700
rect 25452 35606 25508 35644
rect 26012 35698 26068 36204
rect 26124 36036 26180 37214
rect 26124 35970 26180 35980
rect 26236 36372 26292 37326
rect 27804 37378 27860 37390
rect 27804 37326 27806 37378
rect 27858 37326 27860 37378
rect 26908 37266 26964 37278
rect 26908 37214 26910 37266
rect 26962 37214 26964 37266
rect 26012 35646 26014 35698
rect 26066 35646 26068 35698
rect 26012 35634 26068 35646
rect 25228 35476 25284 35486
rect 24892 35252 24948 35262
rect 24892 35026 24948 35196
rect 24892 34974 24894 35026
rect 24946 34974 24948 35026
rect 24892 34962 24948 34974
rect 25228 34914 25284 35420
rect 26236 35476 26292 36316
rect 26460 36484 26516 36494
rect 26460 35812 26516 36428
rect 26908 36370 26964 37214
rect 27244 37268 27300 37278
rect 27804 37268 27860 37326
rect 29820 37378 29876 38668
rect 29932 38612 30100 38668
rect 29932 37490 29988 38612
rect 30156 38500 30212 39228
rect 30268 39228 30436 39284
rect 30268 38836 30324 39228
rect 30380 39060 30436 39070
rect 30380 38966 30436 39004
rect 30828 39058 30884 40348
rect 30828 39006 30830 39058
rect 30882 39006 30884 39058
rect 30492 38948 30548 38958
rect 30492 38854 30548 38892
rect 30604 38836 30660 38846
rect 30268 38780 30436 38836
rect 30044 38444 30212 38500
rect 30268 38612 30324 38622
rect 30044 38050 30100 38444
rect 30156 38164 30212 38174
rect 30268 38164 30324 38556
rect 30156 38162 30324 38164
rect 30156 38110 30158 38162
rect 30210 38110 30324 38162
rect 30156 38108 30324 38110
rect 30156 38098 30212 38108
rect 30044 37998 30046 38050
rect 30098 37998 30100 38050
rect 30044 37986 30100 37998
rect 30268 37940 30324 37950
rect 30380 37940 30436 38780
rect 30604 38742 30660 38780
rect 30828 38164 30884 39006
rect 31276 39284 31332 40348
rect 31612 40516 31668 41916
rect 33068 41970 33124 41982
rect 33068 41918 33070 41970
rect 33122 41918 33124 41970
rect 32508 41860 32564 41870
rect 33068 41860 33124 41918
rect 32508 41858 33124 41860
rect 32508 41806 32510 41858
rect 32562 41806 33124 41858
rect 32508 41804 33124 41806
rect 33852 41970 33908 41982
rect 33852 41918 33854 41970
rect 33906 41918 33908 41970
rect 32508 41794 32564 41804
rect 32508 41300 32564 41310
rect 32396 41244 32508 41300
rect 31612 40402 31668 40460
rect 31612 40350 31614 40402
rect 31666 40350 31668 40402
rect 31612 40338 31668 40350
rect 31836 41186 31892 41198
rect 31836 41134 31838 41186
rect 31890 41134 31892 41186
rect 31836 40514 31892 41134
rect 31836 40462 31838 40514
rect 31890 40462 31892 40514
rect 31836 39620 31892 40462
rect 32172 40404 32228 40414
rect 31836 39554 31892 39564
rect 31948 40402 32228 40404
rect 31948 40350 32174 40402
rect 32226 40350 32228 40402
rect 31948 40348 32228 40350
rect 31276 38946 31332 39228
rect 31948 39058 32004 40348
rect 32172 40338 32228 40348
rect 32060 39732 32116 39742
rect 32060 39638 32116 39676
rect 31948 39006 31950 39058
rect 32002 39006 32004 39058
rect 31948 38994 32004 39006
rect 31276 38894 31278 38946
rect 31330 38894 31332 38946
rect 31276 38882 31332 38894
rect 31500 38946 31556 38958
rect 31500 38894 31502 38946
rect 31554 38894 31556 38946
rect 30716 38052 30772 38062
rect 30828 38052 30884 38108
rect 30716 38050 30884 38052
rect 30716 37998 30718 38050
rect 30770 37998 30884 38050
rect 30716 37996 30884 37998
rect 30716 37986 30772 37996
rect 30268 37938 30436 37940
rect 30268 37886 30270 37938
rect 30322 37886 30436 37938
rect 30268 37884 30436 37886
rect 30268 37874 30324 37884
rect 31500 37828 31556 38894
rect 32396 38836 32452 41244
rect 32508 41234 32564 41244
rect 32508 41074 32564 41086
rect 32508 41022 32510 41074
rect 32562 41022 32564 41074
rect 32508 40626 32564 41022
rect 32508 40574 32510 40626
rect 32562 40574 32564 40626
rect 32508 40562 32564 40574
rect 32508 39620 32564 39630
rect 32564 39564 32676 39620
rect 32508 39526 32564 39564
rect 32508 38836 32564 38846
rect 32396 38834 32564 38836
rect 32396 38782 32510 38834
rect 32562 38782 32564 38834
rect 32396 38780 32564 38782
rect 32508 38770 32564 38780
rect 32620 38836 32676 39564
rect 32620 38770 32676 38780
rect 31612 38724 31668 38762
rect 31612 38658 31668 38668
rect 32284 38724 32340 38762
rect 32284 38658 32340 38668
rect 31836 37828 31892 37838
rect 31500 37826 31892 37828
rect 31500 37774 31838 37826
rect 31890 37774 31892 37826
rect 31500 37772 31892 37774
rect 29932 37438 29934 37490
rect 29986 37438 29988 37490
rect 29932 37426 29988 37438
rect 29820 37326 29822 37378
rect 29874 37326 29876 37378
rect 29820 37314 29876 37326
rect 28028 37268 28084 37278
rect 27244 37266 27860 37268
rect 27244 37214 27246 37266
rect 27298 37214 27860 37266
rect 27244 37212 27860 37214
rect 27916 37266 28084 37268
rect 27916 37214 28030 37266
rect 28082 37214 28084 37266
rect 27916 37212 28084 37214
rect 27132 37044 27188 37054
rect 26908 36318 26910 36370
rect 26962 36318 26964 36370
rect 26908 35924 26964 36318
rect 26908 35858 26964 35868
rect 27020 37042 27188 37044
rect 27020 36990 27134 37042
rect 27186 36990 27188 37042
rect 27020 36988 27188 36990
rect 26460 35746 26516 35756
rect 26236 35410 26292 35420
rect 26348 35700 26404 35710
rect 26124 35028 26180 35038
rect 26124 34934 26180 34972
rect 25228 34862 25230 34914
rect 25282 34862 25284 34914
rect 25228 34850 25284 34862
rect 25340 34860 26068 34916
rect 25340 34802 25396 34860
rect 25340 34750 25342 34802
rect 25394 34750 25396 34802
rect 25340 34738 25396 34750
rect 25564 34690 25620 34702
rect 25564 34638 25566 34690
rect 25618 34638 25620 34690
rect 24780 34132 24836 34142
rect 24780 34038 24836 34076
rect 25452 34018 25508 34030
rect 25452 33966 25454 34018
rect 25506 33966 25508 34018
rect 25340 33572 25396 33582
rect 24668 33070 24670 33122
rect 24722 33070 24724 33122
rect 24668 33012 24724 33070
rect 25004 33124 25060 33134
rect 25004 33030 25060 33068
rect 24668 32946 24724 32956
rect 24668 32788 24724 32798
rect 24668 32694 24724 32732
rect 24332 32582 24388 32620
rect 22988 32564 23044 32574
rect 22988 32450 23044 32508
rect 25340 32564 25396 33516
rect 25452 32788 25508 33966
rect 25564 34020 25620 34638
rect 25900 34690 25956 34702
rect 25900 34638 25902 34690
rect 25954 34638 25956 34690
rect 25788 34244 25844 34254
rect 25788 34150 25844 34188
rect 25564 33954 25620 33964
rect 25676 34130 25732 34142
rect 25676 34078 25678 34130
rect 25730 34078 25732 34130
rect 25676 33124 25732 34078
rect 25788 33572 25844 33582
rect 25900 33572 25956 34638
rect 26012 34690 26068 34860
rect 26012 34638 26014 34690
rect 26066 34638 26068 34690
rect 26012 34356 26068 34638
rect 26236 34692 26292 34702
rect 26236 34598 26292 34636
rect 26012 34300 26180 34356
rect 25844 33516 25956 33572
rect 25788 33506 25844 33516
rect 25676 33058 25732 33068
rect 25788 33348 25844 33358
rect 25564 32788 25620 32798
rect 25452 32732 25564 32788
rect 25564 32722 25620 32732
rect 25788 32786 25844 33292
rect 25900 33236 25956 33246
rect 25900 33142 25956 33180
rect 26124 33012 26180 34300
rect 26236 34132 26292 34142
rect 26348 34132 26404 35644
rect 27020 34914 27076 36988
rect 27132 36978 27188 36988
rect 27132 36484 27188 36494
rect 27244 36484 27300 37212
rect 27916 36484 27972 37212
rect 28028 37202 28084 37212
rect 30156 37268 30212 37278
rect 30156 37266 30548 37268
rect 30156 37214 30158 37266
rect 30210 37214 30548 37266
rect 30156 37212 30548 37214
rect 30156 37202 30212 37212
rect 27188 36428 27300 36484
rect 27804 36428 27972 36484
rect 27132 36390 27188 36428
rect 27468 36372 27524 36382
rect 27468 36278 27524 36316
rect 27244 36258 27300 36270
rect 27244 36206 27246 36258
rect 27298 36206 27300 36258
rect 27244 35028 27300 36206
rect 27356 36258 27412 36270
rect 27356 36206 27358 36258
rect 27410 36206 27412 36258
rect 27356 36036 27412 36206
rect 27356 35970 27412 35980
rect 27804 35252 27860 36428
rect 28028 36370 28084 36382
rect 28028 36318 28030 36370
rect 28082 36318 28084 36370
rect 27916 36260 27972 36270
rect 27916 36166 27972 36204
rect 28028 35588 28084 36318
rect 30380 35812 30436 35822
rect 29036 35700 29092 35710
rect 29036 35698 29204 35700
rect 29036 35646 29038 35698
rect 29090 35646 29204 35698
rect 29036 35644 29204 35646
rect 29036 35634 29092 35644
rect 28364 35588 28420 35598
rect 28028 35586 28420 35588
rect 28028 35534 28366 35586
rect 28418 35534 28420 35586
rect 28028 35532 28420 35534
rect 27804 35186 27860 35196
rect 27356 35028 27412 35038
rect 27244 35026 27412 35028
rect 27244 34974 27358 35026
rect 27410 34974 27412 35026
rect 27244 34972 27412 34974
rect 27356 34962 27412 34972
rect 27020 34862 27022 34914
rect 27074 34862 27076 34914
rect 27020 34850 27076 34862
rect 27468 34914 27524 34926
rect 27468 34862 27470 34914
rect 27522 34862 27524 34914
rect 26460 34804 26516 34814
rect 26516 34748 26628 34804
rect 26460 34710 26516 34748
rect 26460 34356 26516 34366
rect 26460 34262 26516 34300
rect 26236 34130 26404 34132
rect 26236 34078 26238 34130
rect 26290 34078 26404 34130
rect 26236 34076 26404 34078
rect 26236 34066 26292 34076
rect 25788 32734 25790 32786
rect 25842 32734 25844 32786
rect 25788 32722 25844 32734
rect 25900 32956 26180 33012
rect 26236 33236 26292 33246
rect 25340 32498 25396 32508
rect 25900 32562 25956 32956
rect 26124 32788 26180 32798
rect 26236 32788 26292 33180
rect 26124 32786 26292 32788
rect 26124 32734 26126 32786
rect 26178 32734 26292 32786
rect 26124 32732 26292 32734
rect 26124 32722 26180 32732
rect 25900 32510 25902 32562
rect 25954 32510 25956 32562
rect 22988 32398 22990 32450
rect 23042 32398 23044 32450
rect 22988 32386 23044 32398
rect 23436 31778 23492 31790
rect 23436 31726 23438 31778
rect 23490 31726 23492 31778
rect 22204 30818 22260 30828
rect 22764 30884 22820 30894
rect 21308 30772 21364 30782
rect 20972 30146 21028 30156
rect 21084 30770 21364 30772
rect 21084 30718 21310 30770
rect 21362 30718 21364 30770
rect 21084 30716 21364 30718
rect 21084 29988 21140 30716
rect 21308 30706 21364 30716
rect 21644 30100 21700 30110
rect 21644 30006 21700 30044
rect 20636 29932 21140 29988
rect 21308 29986 21364 29998
rect 21308 29934 21310 29986
rect 21362 29934 21364 29986
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20636 29538 20692 29932
rect 20636 29486 20638 29538
rect 20690 29486 20692 29538
rect 20636 29474 20692 29486
rect 19852 29428 19908 29438
rect 18956 26870 19012 26908
rect 19068 26852 19348 26908
rect 19516 29426 19908 29428
rect 19516 29374 19854 29426
rect 19906 29374 19908 29426
rect 19516 29372 19908 29374
rect 19068 26514 19124 26852
rect 19068 26462 19070 26514
rect 19122 26462 19124 26514
rect 18732 26292 18788 26302
rect 18620 25396 18676 25406
rect 17948 24836 18004 24846
rect 17948 24742 18004 24780
rect 18060 24724 18116 24734
rect 18060 24630 18116 24668
rect 18508 24722 18564 24734
rect 18508 24670 18510 24722
rect 18562 24670 18564 24722
rect 18284 24500 18340 24510
rect 18284 23938 18340 24444
rect 18508 24164 18564 24670
rect 18284 23886 18286 23938
rect 18338 23886 18340 23938
rect 18284 23874 18340 23886
rect 18396 24108 18508 24164
rect 17836 23154 17892 23166
rect 17836 23102 17838 23154
rect 17890 23102 17892 23154
rect 17836 23044 17892 23102
rect 18396 23154 18452 24108
rect 18508 24098 18564 24108
rect 18396 23102 18398 23154
rect 18450 23102 18452 23154
rect 18396 23090 18452 23102
rect 17836 22978 17892 22988
rect 18508 22930 18564 22942
rect 18508 22878 18510 22930
rect 18562 22878 18564 22930
rect 18508 22484 18564 22878
rect 18508 22418 18564 22428
rect 18172 22370 18228 22382
rect 18172 22318 18174 22370
rect 18226 22318 18228 22370
rect 17724 21700 17780 21710
rect 17724 21606 17780 21644
rect 17948 21586 18004 21598
rect 17948 21534 17950 21586
rect 18002 21534 18004 21586
rect 17948 21028 18004 21534
rect 17948 20962 18004 20972
rect 18172 21476 18228 22318
rect 18620 22260 18676 25340
rect 18732 23716 18788 26236
rect 19068 24836 19124 26462
rect 19292 26290 19348 26302
rect 19292 26238 19294 26290
rect 19346 26238 19348 26290
rect 19292 25396 19348 26238
rect 19292 25330 19348 25340
rect 18844 24724 18900 24734
rect 18844 24630 18900 24668
rect 18844 23940 18900 23950
rect 19068 23940 19124 24780
rect 19180 25282 19236 25294
rect 19180 25230 19182 25282
rect 19234 25230 19236 25282
rect 19180 24500 19236 25230
rect 19180 24434 19236 24444
rect 19404 24164 19460 24174
rect 19516 24164 19572 29372
rect 19852 29362 19908 29372
rect 21308 29428 21364 29934
rect 20636 28644 20692 28654
rect 20636 28550 20692 28588
rect 21308 28644 21364 29372
rect 22764 29314 22820 30828
rect 23436 30212 23492 31726
rect 23884 31780 23940 31790
rect 23884 31778 24276 31780
rect 23884 31726 23886 31778
rect 23938 31726 24276 31778
rect 23884 31724 24276 31726
rect 23884 31714 23940 31724
rect 24220 31218 24276 31724
rect 25900 31668 25956 32510
rect 26348 32676 26404 32686
rect 26572 32676 26628 34748
rect 27244 34692 27300 34702
rect 26796 34020 26852 34030
rect 26796 33926 26852 33964
rect 27020 33348 27076 33358
rect 27020 33346 27188 33348
rect 27020 33294 27022 33346
rect 27074 33294 27188 33346
rect 27020 33292 27188 33294
rect 27020 33282 27076 33292
rect 26908 33236 26964 33246
rect 26796 33234 26964 33236
rect 26796 33182 26910 33234
rect 26962 33182 26964 33234
rect 26796 33180 26964 33182
rect 26796 32788 26852 33180
rect 26908 33170 26964 33180
rect 27132 33124 27188 33292
rect 26348 32674 26628 32676
rect 26348 32622 26350 32674
rect 26402 32622 26628 32674
rect 26348 32620 26628 32622
rect 26684 32676 26740 32686
rect 26012 32452 26068 32462
rect 26012 32358 26068 32396
rect 26348 31948 26404 32620
rect 26684 32562 26740 32620
rect 26684 32510 26686 32562
rect 26738 32510 26740 32562
rect 26684 32498 26740 32510
rect 25900 31602 25956 31612
rect 26236 31892 26404 31948
rect 24220 31166 24222 31218
rect 24274 31166 24276 31218
rect 24220 31154 24276 31166
rect 26236 31556 26292 31892
rect 26796 31780 26852 32732
rect 26908 33012 26964 33022
rect 26908 32674 26964 32956
rect 26908 32622 26910 32674
rect 26962 32622 26964 32674
rect 26908 32610 26964 32622
rect 27020 32564 27076 32574
rect 27020 32470 27076 32508
rect 27132 32340 27188 33068
rect 27244 32562 27300 34636
rect 27356 34244 27412 34254
rect 27468 34244 27524 34862
rect 27356 34242 27468 34244
rect 27356 34190 27358 34242
rect 27410 34190 27468 34242
rect 27356 34188 27468 34190
rect 27356 33458 27412 34188
rect 27468 34150 27524 34188
rect 27692 34916 27748 34926
rect 27356 33406 27358 33458
rect 27410 33406 27412 33458
rect 27356 33394 27412 33406
rect 27692 32786 27748 34860
rect 28140 34804 28196 34814
rect 28140 34710 28196 34748
rect 28364 34692 28420 35532
rect 28700 35588 28756 35598
rect 28700 35494 28756 35532
rect 28812 35586 28868 35598
rect 28812 35534 28814 35586
rect 28866 35534 28868 35586
rect 28364 34626 28420 34636
rect 28700 34804 28756 34814
rect 28588 34356 28644 34366
rect 28476 34300 28588 34356
rect 28252 34132 28308 34142
rect 28252 34038 28308 34076
rect 27692 32734 27694 32786
rect 27746 32734 27748 32786
rect 27692 32722 27748 32734
rect 28028 33684 28084 33694
rect 28028 32786 28084 33628
rect 28028 32734 28030 32786
rect 28082 32734 28084 32786
rect 28028 32722 28084 32734
rect 28476 32674 28532 34300
rect 28588 34290 28644 34300
rect 28476 32622 28478 32674
rect 28530 32622 28532 32674
rect 28476 32610 28532 32622
rect 28700 32676 28756 34748
rect 28700 32610 28756 32620
rect 27244 32510 27246 32562
rect 27298 32510 27300 32562
rect 27244 32498 27300 32510
rect 28812 32564 28868 35534
rect 29148 34914 29204 35644
rect 29148 34862 29150 34914
rect 29202 34862 29204 34914
rect 29148 34356 29204 34862
rect 29372 35698 29428 35710
rect 29372 35646 29374 35698
rect 29426 35646 29428 35698
rect 29372 35138 29428 35646
rect 29596 35700 29652 35710
rect 29596 35698 30100 35700
rect 29596 35646 29598 35698
rect 29650 35646 30100 35698
rect 29596 35644 30100 35646
rect 29596 35634 29652 35644
rect 29372 35086 29374 35138
rect 29426 35086 29428 35138
rect 29372 34916 29428 35086
rect 29708 35474 29764 35486
rect 29708 35422 29710 35474
rect 29762 35422 29764 35474
rect 29708 35028 29764 35422
rect 29372 34850 29428 34860
rect 29596 34914 29652 34926
rect 29596 34862 29598 34914
rect 29650 34862 29652 34914
rect 29484 34692 29540 34702
rect 29148 34290 29204 34300
rect 29372 34690 29540 34692
rect 29372 34638 29486 34690
rect 29538 34638 29540 34690
rect 29372 34636 29540 34638
rect 28924 34132 28980 34142
rect 28924 34038 28980 34076
rect 29260 33346 29316 33358
rect 29260 33294 29262 33346
rect 29314 33294 29316 33346
rect 29260 32900 29316 33294
rect 28924 32844 29316 32900
rect 28924 32786 28980 32844
rect 28924 32734 28926 32786
rect 28978 32734 28980 32786
rect 28924 32722 28980 32734
rect 29036 32676 29092 32686
rect 29036 32582 29092 32620
rect 29372 32674 29428 34636
rect 29484 34626 29540 34636
rect 29596 34356 29652 34862
rect 29372 32622 29374 32674
rect 29426 32622 29428 32674
rect 29372 32610 29428 32622
rect 29484 34300 29652 34356
rect 29484 34130 29540 34300
rect 29484 34078 29486 34130
rect 29538 34078 29540 34130
rect 28812 32562 28980 32564
rect 28812 32510 28814 32562
rect 28866 32510 28980 32562
rect 28812 32508 28980 32510
rect 28812 32498 28868 32508
rect 27916 32452 27972 32462
rect 28924 32452 28980 32508
rect 29484 32452 29540 34078
rect 29708 34020 29764 34972
rect 29596 33964 29764 34020
rect 29932 34804 29988 34814
rect 29932 34018 29988 34748
rect 29932 33966 29934 34018
rect 29986 33966 29988 34018
rect 29596 32786 29652 33964
rect 29932 33954 29988 33966
rect 29708 33348 29764 33358
rect 30044 33348 30100 35644
rect 30380 34242 30436 35756
rect 30380 34190 30382 34242
rect 30434 34190 30436 34242
rect 30380 34178 30436 34190
rect 29708 33346 30100 33348
rect 29708 33294 29710 33346
rect 29762 33294 30100 33346
rect 29708 33292 30100 33294
rect 29708 33282 29764 33292
rect 30156 33236 30212 33246
rect 30156 33142 30212 33180
rect 29596 32734 29598 32786
rect 29650 32734 29652 32786
rect 29596 32722 29652 32734
rect 28924 32396 29540 32452
rect 27916 32358 27972 32396
rect 26908 32284 27188 32340
rect 26908 32002 26964 32284
rect 26908 31950 26910 32002
rect 26962 31950 26964 32002
rect 26908 31938 26964 31950
rect 27132 31948 27188 32284
rect 29708 32338 29764 32350
rect 29708 32286 29710 32338
rect 29762 32286 29764 32338
rect 27132 31892 27412 31948
rect 26796 31724 26964 31780
rect 25676 31106 25732 31118
rect 25676 31054 25678 31106
rect 25730 31054 25732 31106
rect 24556 30994 24612 31006
rect 24556 30942 24558 30994
rect 24610 30942 24612 30994
rect 23548 30212 23604 30222
rect 23436 30210 23604 30212
rect 23436 30158 23550 30210
rect 23602 30158 23604 30210
rect 23436 30156 23604 30158
rect 23548 29540 23604 30156
rect 23996 30212 24052 30222
rect 23996 30210 24388 30212
rect 23996 30158 23998 30210
rect 24050 30158 24388 30210
rect 23996 30156 24388 30158
rect 23996 30146 24052 30156
rect 24332 29650 24388 30156
rect 24332 29598 24334 29650
rect 24386 29598 24388 29650
rect 24332 29586 24388 29598
rect 24556 29652 24612 30942
rect 24556 29586 24612 29596
rect 24780 29764 24836 29774
rect 23660 29540 23716 29550
rect 23548 29538 23716 29540
rect 23548 29486 23662 29538
rect 23714 29486 23716 29538
rect 23548 29484 23716 29486
rect 22764 29262 22766 29314
rect 22818 29262 22820 29314
rect 22764 29250 22820 29262
rect 21308 28578 21364 28588
rect 20300 28420 20356 28430
rect 20300 28418 20468 28420
rect 20300 28366 20302 28418
rect 20354 28366 20468 28418
rect 20300 28364 20468 28366
rect 20300 28354 20356 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20188 27860 20244 27870
rect 20188 27298 20244 27804
rect 20188 27246 20190 27298
rect 20242 27246 20244 27298
rect 20188 27234 20244 27246
rect 20300 27748 20356 27758
rect 19628 27186 19684 27198
rect 19628 27134 19630 27186
rect 19682 27134 19684 27186
rect 19628 26292 19684 27134
rect 20300 27186 20356 27692
rect 20300 27134 20302 27186
rect 20354 27134 20356 27186
rect 20300 27122 20356 27134
rect 20412 26852 20468 28364
rect 21420 27970 21476 27982
rect 21420 27918 21422 27970
rect 21474 27918 21476 27970
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26226 19684 26236
rect 19852 26180 19908 26190
rect 20300 26180 20356 26190
rect 19852 26086 19908 26124
rect 20188 26178 20356 26180
rect 20188 26126 20302 26178
rect 20354 26126 20356 26178
rect 20188 26124 20356 26126
rect 19740 26068 19796 26078
rect 19628 26066 19796 26068
rect 19628 26014 19742 26066
rect 19794 26014 19796 26066
rect 19628 26012 19796 26014
rect 19628 25284 19684 26012
rect 19740 26002 19796 26012
rect 19740 25732 19796 25742
rect 19740 25638 19796 25676
rect 19964 25396 20020 25406
rect 20188 25396 20244 26124
rect 20300 26114 20356 26124
rect 20412 26180 20468 26796
rect 20860 27748 20916 27758
rect 20860 26290 20916 27692
rect 21420 27298 21476 27918
rect 21980 27748 22036 27758
rect 21980 27654 22036 27692
rect 21420 27246 21422 27298
rect 21474 27246 21476 27298
rect 21420 27234 21476 27246
rect 21308 26962 21364 26974
rect 21308 26910 21310 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 21308 26852 21476 26908
rect 21308 26786 21364 26796
rect 20860 26238 20862 26290
rect 20914 26238 20916 26290
rect 20860 26226 20916 26238
rect 21308 26292 21364 26302
rect 21308 26198 21364 26236
rect 20412 26114 20468 26124
rect 21420 25620 21476 26852
rect 22540 26404 22596 26414
rect 22540 25730 22596 26348
rect 23548 26404 23604 26414
rect 23548 26310 23604 26348
rect 22540 25678 22542 25730
rect 22594 25678 22596 25730
rect 22540 25666 22596 25678
rect 21420 25526 21476 25564
rect 22428 25620 22484 25630
rect 22428 25526 22484 25564
rect 20020 25340 20244 25396
rect 19964 25302 20020 25340
rect 19628 25218 19684 25228
rect 20300 25282 20356 25294
rect 20300 25230 20302 25282
rect 20354 25230 20356 25282
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20300 24948 20356 25230
rect 20300 24882 20356 24892
rect 21308 25282 21364 25294
rect 21308 25230 21310 25282
rect 21362 25230 21364 25282
rect 21308 24946 21364 25230
rect 21308 24894 21310 24946
rect 21362 24894 21364 24946
rect 21308 24882 21364 24894
rect 21980 24948 22036 24958
rect 21980 24854 22036 24892
rect 22540 24836 22596 24846
rect 22540 24742 22596 24780
rect 23660 24836 23716 29484
rect 23996 29426 24052 29438
rect 23996 29374 23998 29426
rect 24050 29374 24052 29426
rect 23996 28420 24052 29374
rect 24668 29428 24724 29438
rect 24668 29334 24724 29372
rect 24780 28642 24836 29708
rect 25228 29764 25284 29774
rect 25228 29204 25284 29708
rect 25676 29764 25732 31054
rect 26012 31108 26068 31118
rect 26012 31014 26068 31052
rect 26236 30884 26292 31500
rect 25676 29698 25732 29708
rect 26012 30828 26292 30884
rect 26348 31554 26404 31566
rect 26348 31502 26350 31554
rect 26402 31502 26404 31554
rect 25340 29652 25396 29662
rect 25340 29558 25396 29596
rect 25676 29428 25732 29438
rect 26012 29428 26068 30828
rect 26236 29764 26292 29774
rect 26236 29538 26292 29708
rect 26348 29652 26404 31502
rect 26684 31106 26740 31118
rect 26684 31054 26686 31106
rect 26738 31054 26740 31106
rect 26460 29988 26516 29998
rect 26460 29894 26516 29932
rect 26348 29586 26404 29596
rect 26236 29486 26238 29538
rect 26290 29486 26292 29538
rect 26236 29474 26292 29486
rect 26684 29540 26740 31054
rect 26908 30772 26964 31724
rect 27356 31778 27412 31892
rect 29708 31892 29764 32286
rect 29708 31826 29764 31836
rect 27356 31726 27358 31778
rect 27410 31726 27412 31778
rect 27356 31714 27412 31726
rect 28028 31778 28084 31790
rect 28028 31726 28030 31778
rect 28082 31726 28084 31778
rect 27244 31668 27300 31678
rect 27132 31556 27188 31566
rect 27132 31462 27188 31500
rect 27020 31444 27076 31454
rect 27020 31218 27076 31388
rect 27020 31166 27022 31218
rect 27074 31166 27076 31218
rect 27020 31154 27076 31166
rect 27244 30996 27300 31612
rect 27804 31668 27860 31678
rect 27804 31574 27860 31612
rect 27916 31444 27972 31454
rect 27916 31218 27972 31388
rect 27916 31166 27918 31218
rect 27970 31166 27972 31218
rect 27916 31154 27972 31166
rect 27244 30940 27412 30996
rect 27244 30772 27300 30782
rect 26908 30770 27300 30772
rect 26908 30718 27246 30770
rect 27298 30718 27300 30770
rect 26908 30716 27300 30718
rect 26908 30436 26964 30716
rect 27244 30706 27300 30716
rect 27020 30436 27076 30446
rect 26908 30434 27076 30436
rect 26908 30382 27022 30434
rect 27074 30382 27076 30434
rect 26908 30380 27076 30382
rect 27020 30370 27076 30380
rect 27244 29986 27300 29998
rect 27244 29934 27246 29986
rect 27298 29934 27300 29986
rect 26684 29474 26740 29484
rect 27132 29764 27188 29774
rect 25676 29426 26068 29428
rect 25676 29374 25678 29426
rect 25730 29374 26068 29426
rect 25676 29372 26068 29374
rect 26460 29426 26516 29438
rect 26460 29374 26462 29426
rect 26514 29374 26516 29426
rect 25676 29362 25732 29372
rect 25228 29148 25396 29204
rect 24780 28590 24782 28642
rect 24834 28590 24836 28642
rect 24780 28578 24836 28590
rect 25004 28642 25060 28654
rect 25004 28590 25006 28642
rect 25058 28590 25060 28642
rect 24444 28420 24500 28430
rect 25004 28420 25060 28590
rect 23996 28418 25060 28420
rect 23996 28366 24446 28418
rect 24498 28366 25060 28418
rect 23996 28364 25060 28366
rect 25116 28644 25172 28654
rect 23996 27748 24052 27758
rect 23996 27654 24052 27692
rect 24332 27074 24388 28364
rect 24444 28354 24500 28364
rect 24668 28084 24724 28094
rect 25116 28084 25172 28588
rect 24668 28082 25172 28084
rect 24668 28030 24670 28082
rect 24722 28030 25172 28082
rect 24668 28028 25172 28030
rect 24668 28018 24724 28028
rect 25228 27972 25284 27982
rect 24780 27970 25284 27972
rect 24780 27918 25230 27970
rect 25282 27918 25284 27970
rect 24780 27916 25284 27918
rect 24444 27860 24500 27870
rect 24444 27766 24500 27804
rect 24332 27022 24334 27074
rect 24386 27022 24388 27074
rect 24332 27010 24388 27022
rect 24780 27074 24836 27916
rect 25228 27906 25284 27916
rect 24780 27022 24782 27074
rect 24834 27022 24836 27074
rect 24780 27010 24836 27022
rect 23996 26292 24052 26302
rect 23996 25732 24052 26236
rect 23996 25638 24052 25676
rect 24108 26178 24164 26190
rect 24108 26126 24110 26178
rect 24162 26126 24164 26178
rect 24108 25618 24164 26126
rect 24108 25566 24110 25618
rect 24162 25566 24164 25618
rect 24108 25554 24164 25566
rect 25116 25732 25172 25742
rect 25116 25394 25172 25676
rect 25116 25342 25118 25394
rect 25170 25342 25172 25394
rect 25116 25330 25172 25342
rect 23660 24770 23716 24780
rect 24108 24836 24164 24846
rect 25228 24836 25284 24846
rect 19404 24162 19572 24164
rect 19404 24110 19406 24162
rect 19458 24110 19572 24162
rect 19404 24108 19572 24110
rect 19628 24500 19684 24510
rect 19404 24098 19460 24108
rect 18844 23938 19124 23940
rect 18844 23886 18846 23938
rect 18898 23886 19124 23938
rect 18844 23884 19124 23886
rect 18844 23874 18900 23884
rect 19292 23826 19348 23838
rect 19292 23774 19294 23826
rect 19346 23774 19348 23826
rect 19068 23716 19124 23726
rect 18732 23660 19012 23716
rect 15260 19908 15316 19918
rect 15260 19814 15316 19852
rect 15372 19794 15428 19806
rect 15372 19742 15374 19794
rect 15426 19742 15428 19794
rect 15372 19684 15428 19742
rect 15036 19628 15428 19684
rect 14812 18676 14868 19516
rect 14028 18610 14084 18620
rect 14588 18620 14868 18676
rect 15372 18676 15428 19628
rect 17052 19236 17108 19246
rect 17052 19142 17108 19180
rect 17388 19234 17444 20636
rect 17500 20636 17668 20692
rect 18172 20802 18228 21420
rect 18508 22204 18676 22260
rect 18844 22594 18900 22606
rect 18844 22542 18846 22594
rect 18898 22542 18900 22594
rect 18508 21140 18564 22204
rect 18844 21810 18900 22542
rect 18844 21758 18846 21810
rect 18898 21758 18900 21810
rect 18844 21746 18900 21758
rect 18732 21588 18788 21598
rect 18732 21494 18788 21532
rect 18620 21364 18676 21374
rect 18620 21270 18676 21308
rect 18956 21252 19012 23660
rect 19068 21924 19124 23660
rect 19180 23154 19236 23166
rect 19180 23102 19182 23154
rect 19234 23102 19236 23154
rect 19180 22148 19236 23102
rect 19292 23044 19348 23774
rect 19516 23156 19572 23166
rect 19628 23156 19684 24444
rect 22428 24500 22484 24510
rect 22428 24406 22484 24444
rect 23772 24500 23828 24510
rect 19740 24164 19796 24174
rect 19740 24070 19796 24108
rect 19852 23826 19908 23838
rect 19852 23774 19854 23826
rect 19906 23774 19908 23826
rect 19852 23716 19908 23774
rect 19852 23650 19908 23660
rect 20300 23716 20356 23726
rect 20300 23622 20356 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20748 23436 21588 23492
rect 19516 23154 19684 23156
rect 19516 23102 19518 23154
rect 19570 23102 19684 23154
rect 19516 23100 19684 23102
rect 20188 23266 20244 23278
rect 20188 23214 20190 23266
rect 20242 23214 20244 23266
rect 19516 23090 19572 23100
rect 19292 22978 19348 22988
rect 19180 22082 19236 22092
rect 19292 22594 19348 22606
rect 19292 22542 19294 22594
rect 19346 22542 19348 22594
rect 19292 22482 19348 22542
rect 19292 22430 19294 22482
rect 19346 22430 19348 22482
rect 19292 21924 19348 22430
rect 20188 22372 20244 23214
rect 20524 23156 20580 23166
rect 20748 23156 20804 23436
rect 21532 23378 21588 23436
rect 21532 23326 21534 23378
rect 21586 23326 21588 23378
rect 21532 23314 21588 23326
rect 20524 23154 20804 23156
rect 20524 23102 20526 23154
rect 20578 23102 20804 23154
rect 20524 23100 20804 23102
rect 20860 23266 20916 23278
rect 20860 23214 20862 23266
rect 20914 23214 20916 23266
rect 20412 22372 20468 22382
rect 20188 22370 20468 22372
rect 20188 22318 20414 22370
rect 20466 22318 20468 22370
rect 20188 22316 20468 22318
rect 19740 22148 19796 22158
rect 19628 22146 19796 22148
rect 19628 22094 19742 22146
rect 19794 22094 19796 22146
rect 19628 22092 19796 22094
rect 19628 21924 19684 22092
rect 19740 22082 19796 22092
rect 20188 22146 20244 22158
rect 20188 22094 20190 22146
rect 20242 22094 20244 22146
rect 19292 21868 19572 21924
rect 19068 21858 19124 21868
rect 18956 21186 19012 21196
rect 19068 21700 19124 21710
rect 18508 21084 18788 21140
rect 18172 20750 18174 20802
rect 18226 20750 18228 20802
rect 18172 20692 18228 20750
rect 17500 19684 17556 20636
rect 18172 20626 18228 20636
rect 17836 20132 17892 20142
rect 17836 20130 18228 20132
rect 17836 20078 17838 20130
rect 17890 20078 18228 20130
rect 17836 20076 18228 20078
rect 17836 20066 17892 20076
rect 17612 20020 17668 20030
rect 17612 19926 17668 19964
rect 17500 19628 18004 19684
rect 17388 19182 17390 19234
rect 17442 19182 17444 19234
rect 17388 19170 17444 19182
rect 16268 19124 16324 19134
rect 12796 18498 12852 18508
rect 13692 18564 13748 18574
rect 13692 18452 13748 18508
rect 12572 18398 12574 18450
rect 12626 18398 12628 18450
rect 12572 18386 12628 18398
rect 13468 18450 13748 18452
rect 13468 18398 13694 18450
rect 13746 18398 13748 18450
rect 13468 18396 13748 18398
rect 13468 17778 13524 18396
rect 13692 18386 13748 18396
rect 14476 18450 14532 18462
rect 14476 18398 14478 18450
rect 14530 18398 14532 18450
rect 13468 17726 13470 17778
rect 13522 17726 13524 17778
rect 13468 17714 13524 17726
rect 13804 18228 13860 18238
rect 13804 17780 13860 18172
rect 14476 17892 14532 18398
rect 14476 17826 14532 17836
rect 13804 17714 13860 17724
rect 14028 17668 14084 17678
rect 12460 16772 12516 16828
rect 13132 16994 13188 17006
rect 13132 16942 13134 16994
rect 13186 16942 13188 16994
rect 12796 16772 12852 16782
rect 12460 16770 12852 16772
rect 12460 16718 12798 16770
rect 12850 16718 12852 16770
rect 12460 16716 12852 16718
rect 12796 16706 12852 16716
rect 13132 16772 13188 16942
rect 13356 16884 13412 16894
rect 13132 16706 13188 16716
rect 13244 16882 13412 16884
rect 13244 16830 13358 16882
rect 13410 16830 13412 16882
rect 13244 16828 13412 16830
rect 13244 16436 13300 16828
rect 13356 16818 13412 16828
rect 14028 16884 14084 17612
rect 14028 16882 14532 16884
rect 14028 16830 14030 16882
rect 14082 16830 14532 16882
rect 14028 16828 14532 16830
rect 14028 16818 14084 16828
rect 12796 16380 13300 16436
rect 14252 16660 14308 16670
rect 12796 16322 12852 16380
rect 12796 16270 12798 16322
rect 12850 16270 12852 16322
rect 12796 16258 12852 16270
rect 12460 16212 12516 16222
rect 12180 16156 12404 16212
rect 12124 16146 12180 16156
rect 11788 15934 11790 15986
rect 11842 15934 11844 15986
rect 11788 15922 11844 15934
rect 11900 15988 11956 15998
rect 10108 15810 10164 15820
rect 10556 15876 10612 15886
rect 11116 15876 11172 15886
rect 10556 15874 11172 15876
rect 10556 15822 10558 15874
rect 10610 15822 11118 15874
rect 11170 15822 11172 15874
rect 10556 15820 11172 15822
rect 10556 15810 10612 15820
rect 11116 15540 11172 15820
rect 11116 15474 11172 15484
rect 9660 15314 10052 15316
rect 9660 15262 9662 15314
rect 9714 15262 10052 15314
rect 9660 15260 10052 15262
rect 9660 15250 9716 15260
rect 8876 14812 9828 14868
rect 9772 14642 9828 14812
rect 9772 14590 9774 14642
rect 9826 14590 9828 14642
rect 9772 14578 9828 14590
rect 9100 14530 9156 14542
rect 9100 14478 9102 14530
rect 9154 14478 9156 14530
rect 9100 13748 9156 14478
rect 9100 13682 9156 13692
rect 9884 13748 9940 15260
rect 10332 15204 10388 15214
rect 10332 15110 10388 15148
rect 11900 14642 11956 15932
rect 12236 15986 12292 15998
rect 12236 15934 12238 15986
rect 12290 15934 12292 15986
rect 12236 15876 12292 15934
rect 12236 15810 12292 15820
rect 11900 14590 11902 14642
rect 11954 14590 11956 14642
rect 11900 14578 11956 14590
rect 12236 15428 12292 15438
rect 12236 14530 12292 15372
rect 12348 15204 12404 16156
rect 12460 16118 12516 16156
rect 14252 16212 14308 16604
rect 13692 16044 13972 16100
rect 13468 15876 13524 15886
rect 13356 15874 13524 15876
rect 13356 15822 13470 15874
rect 13522 15822 13524 15874
rect 13356 15820 13524 15822
rect 13132 15540 13188 15550
rect 13132 15446 13188 15484
rect 13356 15428 13412 15820
rect 13468 15810 13524 15820
rect 12684 15316 12740 15326
rect 12572 15314 12740 15316
rect 12572 15262 12686 15314
rect 12738 15262 12740 15314
rect 12572 15260 12740 15262
rect 12460 15204 12516 15214
rect 12348 15202 12516 15204
rect 12348 15150 12462 15202
rect 12514 15150 12516 15202
rect 12348 15148 12516 15150
rect 12460 15138 12516 15148
rect 12236 14478 12238 14530
rect 12290 14478 12292 14530
rect 12236 14466 12292 14478
rect 12572 14530 12628 15260
rect 12684 15250 12740 15260
rect 13244 15204 13300 15214
rect 13244 15110 13300 15148
rect 13356 14644 13412 15372
rect 13468 15316 13524 15326
rect 13524 15260 13636 15316
rect 13468 15250 13524 15260
rect 13580 14754 13636 15260
rect 13580 14702 13582 14754
rect 13634 14702 13636 14754
rect 13580 14690 13636 14702
rect 13692 14756 13748 16044
rect 13916 15988 13972 16044
rect 14140 15988 14196 15998
rect 13916 15932 14140 15988
rect 14140 15894 14196 15932
rect 13804 15876 13860 15886
rect 13804 15540 13860 15820
rect 14140 15540 14196 15550
rect 13804 15484 14140 15540
rect 14140 15446 14196 15484
rect 13692 14700 13860 14756
rect 13356 14588 13524 14644
rect 12572 14478 12574 14530
rect 12626 14478 12628 14530
rect 12572 14466 12628 14478
rect 13468 14532 13524 14588
rect 13692 14532 13748 14542
rect 13468 14530 13748 14532
rect 13468 14478 13694 14530
rect 13746 14478 13748 14530
rect 13468 14476 13748 14478
rect 13692 14466 13748 14476
rect 12348 14306 12404 14318
rect 12348 14254 12350 14306
rect 12402 14254 12404 14306
rect 9884 13682 9940 13692
rect 10892 13748 10948 13758
rect 10892 13654 10948 13692
rect 11676 13634 11732 13646
rect 11676 13582 11678 13634
rect 11730 13582 11732 13634
rect 11676 12852 11732 13582
rect 12348 13524 12404 14254
rect 12348 13458 12404 13468
rect 12796 14308 12852 14318
rect 12796 12962 12852 14252
rect 13020 14308 13076 14318
rect 13580 14308 13636 14318
rect 13020 14306 13636 14308
rect 13020 14254 13022 14306
rect 13074 14254 13582 14306
rect 13634 14254 13636 14306
rect 13020 14252 13636 14254
rect 13020 14242 13076 14252
rect 13356 13748 13412 14252
rect 13580 14242 13636 14252
rect 13804 13860 13860 14700
rect 14252 14642 14308 16156
rect 14476 15988 14532 16828
rect 14588 16772 14644 18620
rect 15372 18610 15428 18620
rect 15708 19122 16324 19124
rect 15708 19070 16270 19122
rect 16322 19070 16324 19122
rect 15708 19068 16324 19070
rect 15708 18674 15764 19068
rect 16268 19058 16324 19068
rect 15708 18622 15710 18674
rect 15762 18622 15764 18674
rect 15708 18610 15764 18622
rect 15820 18676 15876 18686
rect 15820 18582 15876 18620
rect 15036 18564 15092 18574
rect 15036 18470 15092 18508
rect 15596 18564 15652 18574
rect 15596 18470 15652 18508
rect 16940 18564 16996 18574
rect 14812 18450 14868 18462
rect 14812 18398 14814 18450
rect 14866 18398 14868 18450
rect 14812 18228 14868 18398
rect 16268 18452 16324 18462
rect 16268 18358 16324 18396
rect 14812 18162 14868 18172
rect 14924 18338 14980 18350
rect 14924 18286 14926 18338
rect 14978 18286 14980 18338
rect 14924 17780 14980 18286
rect 14924 17714 14980 17724
rect 15596 17780 15652 17790
rect 15596 17686 15652 17724
rect 16268 17668 16324 17678
rect 16268 17574 16324 17612
rect 16604 17668 16660 17678
rect 16604 17574 16660 17612
rect 16940 17666 16996 18508
rect 17500 18562 17556 18574
rect 17500 18510 17502 18562
rect 17554 18510 17556 18562
rect 17276 18452 17332 18462
rect 17276 18358 17332 18396
rect 16940 17614 16942 17666
rect 16994 17614 16996 17666
rect 16940 17602 16996 17614
rect 17500 17668 17556 18510
rect 17612 18564 17668 18574
rect 17612 18470 17668 18508
rect 17500 17612 17668 17668
rect 16828 17444 16884 17454
rect 17500 17444 17556 17454
rect 16828 17442 17556 17444
rect 16828 17390 16830 17442
rect 16882 17390 17502 17442
rect 17554 17390 17556 17442
rect 16828 17388 17556 17390
rect 17612 17444 17668 17612
rect 17836 17444 17892 17454
rect 17612 17442 17892 17444
rect 17612 17390 17838 17442
rect 17890 17390 17892 17442
rect 17612 17388 17892 17390
rect 16828 17378 16884 17388
rect 14588 16706 14644 16716
rect 14700 16772 14756 16782
rect 16828 16772 16884 16782
rect 14700 16770 15092 16772
rect 14700 16718 14702 16770
rect 14754 16718 15092 16770
rect 14700 16716 15092 16718
rect 14700 16706 14756 16716
rect 14812 15988 14868 15998
rect 14476 15986 14756 15988
rect 14476 15934 14478 15986
rect 14530 15934 14756 15986
rect 14476 15932 14756 15934
rect 14476 15922 14532 15932
rect 14588 15540 14644 15550
rect 14588 15446 14644 15484
rect 14252 14590 14254 14642
rect 14306 14590 14308 14642
rect 14252 14578 14308 14590
rect 13356 13682 13412 13692
rect 13468 13804 13860 13860
rect 12796 12910 12798 12962
rect 12850 12910 12852 12962
rect 12796 12898 12852 12910
rect 13356 13524 13412 13534
rect 11676 12786 11732 12796
rect 12460 12852 12516 12862
rect 12460 12758 12516 12796
rect 12348 11282 12404 11294
rect 12348 11230 12350 11282
rect 12402 11230 12404 11282
rect 12012 11172 12068 11182
rect 11676 11170 12068 11172
rect 11676 11118 12014 11170
rect 12066 11118 12068 11170
rect 11676 11116 12068 11118
rect 11004 10724 11060 10734
rect 11004 10630 11060 10668
rect 11228 10610 11284 10622
rect 11228 10558 11230 10610
rect 11282 10558 11284 10610
rect 11116 10498 11172 10510
rect 11116 10446 11118 10498
rect 11170 10446 11172 10498
rect 11116 10164 11172 10446
rect 10108 10108 11172 10164
rect 10108 9938 10164 10108
rect 10108 9886 10110 9938
rect 10162 9886 10164 9938
rect 10108 9874 10164 9886
rect 9436 9828 9492 9838
rect 9436 9734 9492 9772
rect 11228 9268 11284 10558
rect 11676 10610 11732 11116
rect 12012 11106 12068 11116
rect 12236 11172 12292 11182
rect 12236 11078 12292 11116
rect 11900 10724 11956 10734
rect 11900 10630 11956 10668
rect 12348 10724 12404 11230
rect 12796 11172 12852 11182
rect 12796 11078 12852 11116
rect 13356 11172 13412 13468
rect 13356 11106 13412 11116
rect 13132 10948 13188 10958
rect 13132 10836 13188 10892
rect 12908 10834 13188 10836
rect 12908 10782 13134 10834
rect 13186 10782 13188 10834
rect 12908 10780 13188 10782
rect 12348 10658 12404 10668
rect 12796 10724 12852 10734
rect 12796 10630 12852 10668
rect 11676 10558 11678 10610
rect 11730 10558 11732 10610
rect 11676 10546 11732 10558
rect 12124 10610 12180 10622
rect 12124 10558 12126 10610
rect 12178 10558 12180 10610
rect 12012 10498 12068 10510
rect 12012 10446 12014 10498
rect 12066 10446 12068 10498
rect 12012 10276 12068 10446
rect 11228 9202 11284 9212
rect 11676 10220 12068 10276
rect 11676 9154 11732 10220
rect 12124 9492 12180 10558
rect 12572 10610 12628 10622
rect 12572 10558 12574 10610
rect 12626 10558 12628 10610
rect 11676 9102 11678 9154
rect 11730 9102 11732 9154
rect 11676 9090 11732 9102
rect 12012 9436 12180 9492
rect 12236 9938 12292 9950
rect 12236 9886 12238 9938
rect 12290 9886 12292 9938
rect 9548 8930 9604 8942
rect 9548 8878 9550 8930
rect 9602 8878 9604 8930
rect 8652 8372 8932 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 8876 6690 8932 8372
rect 9548 8372 9604 8878
rect 9548 8306 9604 8316
rect 11228 8372 11284 8382
rect 11228 8278 11284 8316
rect 11900 8372 11956 8382
rect 11340 8260 11396 8270
rect 11340 8166 11396 8204
rect 11900 8258 11956 8316
rect 11900 8206 11902 8258
rect 11954 8206 11956 8258
rect 11900 8194 11956 8206
rect 12012 8260 12068 9436
rect 12124 8708 12180 8718
rect 12124 8370 12180 8652
rect 12124 8318 12126 8370
rect 12178 8318 12180 8370
rect 12124 8306 12180 8318
rect 12012 8194 12068 8204
rect 12236 8260 12292 9886
rect 12460 9828 12516 9838
rect 12460 9042 12516 9772
rect 12572 9826 12628 10558
rect 12572 9774 12574 9826
rect 12626 9774 12628 9826
rect 12572 9762 12628 9774
rect 12908 9826 12964 10780
rect 13132 10770 13188 10780
rect 12908 9774 12910 9826
rect 12962 9774 12964 9826
rect 12908 9762 12964 9774
rect 13468 9828 13524 13804
rect 13468 9734 13524 9772
rect 13580 13636 13636 13646
rect 13804 13636 13860 13646
rect 13580 11506 13636 13580
rect 13580 11454 13582 11506
rect 13634 11454 13636 11506
rect 12796 9716 12852 9726
rect 12796 9622 12852 9660
rect 13580 9716 13636 11454
rect 13580 9650 13636 9660
rect 13692 13580 13804 13636
rect 12460 8990 12462 9042
rect 12514 8990 12516 9042
rect 12460 8978 12516 8990
rect 12796 9268 12852 9278
rect 12796 9042 12852 9212
rect 12796 8990 12798 9042
rect 12850 8990 12852 9042
rect 12796 8482 12852 8990
rect 12796 8430 12798 8482
rect 12850 8430 12852 8482
rect 12796 8418 12852 8430
rect 13020 9042 13076 9054
rect 13020 8990 13022 9042
rect 13074 8990 13076 9042
rect 12684 8260 12740 8270
rect 12236 8258 12740 8260
rect 12236 8206 12238 8258
rect 12290 8206 12686 8258
rect 12738 8206 12740 8258
rect 12236 8204 12740 8206
rect 12236 8194 12292 8204
rect 12684 8194 12740 8204
rect 10892 8148 10948 8158
rect 8876 6638 8878 6690
rect 8930 6638 8932 6690
rect 8876 6132 8932 6638
rect 9324 8036 9380 8046
rect 9324 6690 9380 7980
rect 10780 8036 10836 8046
rect 10780 7942 10836 7980
rect 10780 7476 10836 7486
rect 10892 7476 10948 8092
rect 11676 8146 11732 8158
rect 11676 8094 11678 8146
rect 11730 8094 11732 8146
rect 10780 7474 10948 7476
rect 10780 7422 10782 7474
rect 10834 7422 10948 7474
rect 10780 7420 10948 7422
rect 11228 7476 11284 7486
rect 11676 7476 11732 8094
rect 13020 8148 13076 8990
rect 13132 9044 13188 9054
rect 13132 8950 13188 8988
rect 13244 9042 13300 9054
rect 13244 8990 13246 9042
rect 13298 8990 13300 9042
rect 13244 8932 13300 8990
rect 13244 8866 13300 8876
rect 13468 9042 13524 9054
rect 13468 8990 13470 9042
rect 13522 8990 13524 9042
rect 13020 8082 13076 8092
rect 13468 8148 13524 8990
rect 13692 8932 13748 13580
rect 13804 13542 13860 13580
rect 14252 13634 14308 13646
rect 14252 13582 14254 13634
rect 14306 13582 14308 13634
rect 14140 13524 14196 13534
rect 14252 13524 14308 13582
rect 14196 13468 14308 13524
rect 14364 13524 14420 13534
rect 14140 13458 14196 13468
rect 14364 12962 14420 13468
rect 14700 12964 14756 15932
rect 14812 15894 14868 15932
rect 15036 15540 15092 16716
rect 16716 16716 16828 16772
rect 16604 16436 16660 16446
rect 15932 16324 15988 16334
rect 15932 16230 15988 16268
rect 15148 16100 15204 16110
rect 15148 16006 15204 16044
rect 16604 16098 16660 16380
rect 16604 16046 16606 16098
rect 16658 16046 16660 16098
rect 15596 15876 15652 15886
rect 15484 15874 15652 15876
rect 15484 15822 15598 15874
rect 15650 15822 15652 15874
rect 15484 15820 15652 15822
rect 15148 15540 15204 15550
rect 15036 15538 15204 15540
rect 15036 15486 15150 15538
rect 15202 15486 15204 15538
rect 15036 15484 15204 15486
rect 15148 15474 15204 15484
rect 15484 15426 15540 15820
rect 15596 15810 15652 15820
rect 16604 15540 16660 16046
rect 16716 15986 16772 16716
rect 16828 16678 16884 16716
rect 17276 16436 17332 16446
rect 17276 16210 17332 16380
rect 17276 16158 17278 16210
rect 17330 16158 17332 16210
rect 17276 16146 17332 16158
rect 17500 16324 17556 17388
rect 17836 17108 17892 17388
rect 17836 17042 17892 17052
rect 16716 15934 16718 15986
rect 16770 15934 16772 15986
rect 16716 15922 16772 15934
rect 17500 15876 17556 16268
rect 17724 15876 17780 15886
rect 17500 15874 17780 15876
rect 17500 15822 17726 15874
rect 17778 15822 17780 15874
rect 17500 15820 17780 15822
rect 16604 15474 16660 15484
rect 17724 15540 17780 15820
rect 17724 15474 17780 15484
rect 15484 15374 15486 15426
rect 15538 15374 15540 15426
rect 15484 15362 15540 15374
rect 15148 14530 15204 14542
rect 15148 14478 15150 14530
rect 15202 14478 15204 14530
rect 14812 14308 14868 14318
rect 14812 14214 14868 14252
rect 15148 13636 15204 14478
rect 15484 14418 15540 14430
rect 15484 14366 15486 14418
rect 15538 14366 15540 14418
rect 15148 13570 15204 13580
rect 15372 13860 15428 13870
rect 14924 12964 14980 12974
rect 14364 12910 14366 12962
rect 14418 12910 14420 12962
rect 14364 12898 14420 12910
rect 14476 12962 14980 12964
rect 14476 12910 14926 12962
rect 14978 12910 14980 12962
rect 14476 12908 14980 12910
rect 14476 12740 14532 12908
rect 14924 12898 14980 12908
rect 14028 12684 14532 12740
rect 14588 12740 14644 12750
rect 14588 12738 14756 12740
rect 14588 12686 14590 12738
rect 14642 12686 14756 12738
rect 14588 12684 14756 12686
rect 14028 12178 14084 12684
rect 14588 12674 14644 12684
rect 14700 12290 14756 12684
rect 14700 12238 14702 12290
rect 14754 12238 14756 12290
rect 14700 12226 14756 12238
rect 14028 12126 14030 12178
rect 14082 12126 14084 12178
rect 14028 12114 14084 12126
rect 15372 10948 15428 13804
rect 15484 13636 15540 14366
rect 15708 14418 15764 14430
rect 15708 14366 15710 14418
rect 15762 14366 15764 14418
rect 15708 14308 15764 14366
rect 16716 14418 16772 14430
rect 16716 14366 16718 14418
rect 16770 14366 16772 14418
rect 16380 14308 16436 14318
rect 15708 14242 15764 14252
rect 15820 14306 16436 14308
rect 15820 14254 16382 14306
rect 16434 14254 16436 14306
rect 15820 14252 16436 14254
rect 15484 13570 15540 13580
rect 15596 13524 15652 13534
rect 15596 13430 15652 13468
rect 15708 13076 15764 13086
rect 15820 13076 15876 14252
rect 16380 14242 16436 14252
rect 15932 14084 15988 14094
rect 15932 13746 15988 14028
rect 15932 13694 15934 13746
rect 15986 13694 15988 13746
rect 15932 13682 15988 13694
rect 16492 13860 16548 13870
rect 16492 13746 16548 13804
rect 16492 13694 16494 13746
rect 16546 13694 16548 13746
rect 16492 13682 16548 13694
rect 16604 13858 16660 13870
rect 16604 13806 16606 13858
rect 16658 13806 16660 13858
rect 15708 13074 15876 13076
rect 15708 13022 15710 13074
rect 15762 13022 15876 13074
rect 15708 13020 15876 13022
rect 15708 13010 15764 13020
rect 16604 12068 16660 13806
rect 16716 12404 16772 14366
rect 17164 14308 17220 14318
rect 17948 14308 18004 19628
rect 18172 19346 18228 20076
rect 18284 20020 18340 20030
rect 18284 19926 18340 19964
rect 18620 19796 18676 19806
rect 18172 19294 18174 19346
rect 18226 19294 18228 19346
rect 18172 19282 18228 19294
rect 18508 19794 18676 19796
rect 18508 19742 18622 19794
rect 18674 19742 18676 19794
rect 18508 19740 18676 19742
rect 18508 19012 18564 19740
rect 18620 19730 18676 19740
rect 18284 18564 18340 18574
rect 18284 18470 18340 18508
rect 18396 17892 18452 17902
rect 18508 17892 18564 18956
rect 18620 18452 18676 18462
rect 18620 18358 18676 18396
rect 18508 17836 18676 17892
rect 18284 17108 18340 17118
rect 18396 17108 18452 17836
rect 18508 17108 18564 17118
rect 18284 17106 18564 17108
rect 18284 17054 18286 17106
rect 18338 17054 18510 17106
rect 18562 17054 18564 17106
rect 18284 17052 18564 17054
rect 18284 17042 18340 17052
rect 18508 15428 18564 17052
rect 18508 15362 18564 15372
rect 18620 15148 18676 17836
rect 18732 17220 18788 21084
rect 19068 20916 19124 21644
rect 19404 21588 19460 21598
rect 19404 21494 19460 21532
rect 19292 21364 19348 21374
rect 18956 20860 19124 20916
rect 19180 21028 19236 21038
rect 19180 20914 19236 20972
rect 19292 21026 19348 21308
rect 19292 20974 19294 21026
rect 19346 20974 19348 21026
rect 19292 20962 19348 20974
rect 19516 20916 19572 21868
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21858 19684 21868
rect 19180 20862 19182 20914
rect 19234 20862 19236 20914
rect 18956 20804 19012 20860
rect 19180 20850 19236 20862
rect 19404 20860 19572 20916
rect 19628 21698 19684 21710
rect 19628 21646 19630 21698
rect 19682 21646 19684 21698
rect 18844 20802 19012 20804
rect 18844 20750 18958 20802
rect 19010 20750 19012 20802
rect 18844 20748 19012 20750
rect 18844 17780 18900 20748
rect 18956 20738 19012 20748
rect 19404 20188 19460 20860
rect 19180 20130 19236 20142
rect 19180 20078 19182 20130
rect 19234 20078 19236 20130
rect 19180 19796 19236 20078
rect 19180 19730 19236 19740
rect 19292 20132 19460 20188
rect 19628 20132 19684 21646
rect 19964 21588 20020 21598
rect 20188 21588 20244 22094
rect 19964 21586 20244 21588
rect 19964 21534 19966 21586
rect 20018 21534 20244 21586
rect 19964 21532 20244 21534
rect 20300 22148 20356 22158
rect 19964 21476 20020 21532
rect 19964 21410 20020 21420
rect 19740 21364 19796 21374
rect 19740 20690 19796 21308
rect 20188 21364 20244 21374
rect 19740 20638 19742 20690
rect 19794 20638 19796 20690
rect 19740 20626 19796 20638
rect 20076 20692 20132 20702
rect 20076 20598 20132 20636
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19292 18228 19348 20132
rect 19628 20066 19684 20076
rect 19964 20244 20020 20254
rect 19404 20018 19460 20030
rect 19404 19966 19406 20018
rect 19458 19966 19460 20018
rect 19404 18452 19460 19966
rect 19964 20018 20020 20188
rect 19964 19966 19966 20018
rect 20018 19966 20020 20018
rect 19964 19954 20020 19966
rect 20188 19236 20244 21308
rect 20300 20020 20356 22092
rect 20412 20244 20468 22316
rect 20524 21364 20580 23100
rect 20860 23044 20916 23214
rect 21196 23268 21252 23278
rect 21196 23174 21252 23212
rect 21756 23156 21812 23166
rect 21644 23154 21812 23156
rect 21644 23102 21758 23154
rect 21810 23102 21812 23154
rect 21644 23100 21812 23102
rect 21644 23044 21700 23100
rect 21756 23090 21812 23100
rect 20860 22988 21700 23044
rect 21420 22148 21476 22158
rect 21084 22146 21476 22148
rect 21084 22094 21422 22146
rect 21474 22094 21476 22146
rect 21084 22092 21476 22094
rect 21084 21700 21140 22092
rect 21420 22082 21476 22092
rect 20524 21298 20580 21308
rect 20636 21644 21140 21700
rect 20636 20916 20692 21644
rect 21532 21588 21588 21598
rect 20524 20860 20692 20916
rect 20748 21474 20804 21486
rect 20748 21422 20750 21474
rect 20802 21422 20804 21474
rect 20524 20802 20580 20860
rect 20524 20750 20526 20802
rect 20578 20750 20580 20802
rect 20524 20738 20580 20750
rect 20748 20690 20804 21422
rect 21532 21026 21588 21532
rect 21532 20974 21534 21026
rect 21586 20974 21588 21026
rect 21532 20962 21588 20974
rect 20748 20638 20750 20690
rect 20802 20638 20804 20690
rect 20748 20626 20804 20638
rect 20412 20178 20468 20188
rect 20636 20132 20692 20142
rect 20636 20038 20692 20076
rect 20300 19964 20468 20020
rect 20300 19796 20356 19806
rect 20300 19346 20356 19740
rect 20300 19294 20302 19346
rect 20354 19294 20356 19346
rect 20300 19282 20356 19294
rect 20188 19170 20244 19180
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19404 18386 19460 18396
rect 19292 18162 19348 18172
rect 18844 17714 18900 17724
rect 19852 18004 19908 18014
rect 19180 17666 19236 17678
rect 19180 17614 19182 17666
rect 19234 17614 19236 17666
rect 18844 17556 18900 17566
rect 19180 17556 19236 17614
rect 19852 17666 19908 17948
rect 19852 17614 19854 17666
rect 19906 17614 19908 17666
rect 19852 17602 19908 17614
rect 20300 17666 20356 17678
rect 20300 17614 20302 17666
rect 20354 17614 20356 17666
rect 19516 17556 19572 17566
rect 18844 17554 19124 17556
rect 18844 17502 18846 17554
rect 18898 17502 19124 17554
rect 18844 17500 19124 17502
rect 19180 17554 19572 17556
rect 19180 17502 19518 17554
rect 19570 17502 19572 17554
rect 19180 17500 19572 17502
rect 18844 17490 18900 17500
rect 19068 17444 19124 17500
rect 19068 17388 19236 17444
rect 18732 17154 18788 17164
rect 18956 17220 19012 17230
rect 18956 16884 19012 17164
rect 18844 16828 19012 16884
rect 19068 17108 19124 17118
rect 19068 16882 19124 17052
rect 19068 16830 19070 16882
rect 19122 16830 19124 16882
rect 18844 16210 18900 16828
rect 19068 16818 19124 16830
rect 19180 16436 19236 17388
rect 19404 16882 19460 16894
rect 19404 16830 19406 16882
rect 19458 16830 19460 16882
rect 19404 16436 19460 16830
rect 18844 16158 18846 16210
rect 18898 16158 18900 16210
rect 18844 16146 18900 16158
rect 18956 16380 19460 16436
rect 18956 15204 19012 16380
rect 19068 16100 19124 16110
rect 19516 16100 19572 17500
rect 19836 17276 20100 17286
rect 19124 16044 19572 16100
rect 19628 17220 19684 17230
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16100 19684 17164
rect 20188 16770 20244 16782
rect 20188 16718 20190 16770
rect 20242 16718 20244 16770
rect 20188 16548 20244 16718
rect 20188 16482 20244 16492
rect 20300 16436 20356 17614
rect 20412 17444 20468 19964
rect 20972 19124 21028 19134
rect 20748 19012 20804 19022
rect 20748 18918 20804 18956
rect 20636 18452 20692 18462
rect 20636 18358 20692 18396
rect 20972 18226 21028 19068
rect 21196 18452 21252 18462
rect 21196 18358 21252 18396
rect 20972 18174 20974 18226
rect 21026 18174 21028 18226
rect 20972 17892 21028 18174
rect 21532 18004 21588 18014
rect 21644 18004 21700 22988
rect 21756 22372 21812 22382
rect 21756 22278 21812 22316
rect 22876 22372 22932 22382
rect 22092 22258 22148 22270
rect 22092 22206 22094 22258
rect 22146 22206 22148 22258
rect 21868 20804 21924 20814
rect 21868 20710 21924 20748
rect 22092 20692 22148 22206
rect 22092 19346 22148 20636
rect 22092 19294 22094 19346
rect 22146 19294 22148 19346
rect 22092 19282 22148 19294
rect 22540 22258 22596 22270
rect 22540 22206 22542 22258
rect 22594 22206 22596 22258
rect 22540 22148 22596 22206
rect 22316 19236 22372 19246
rect 22316 19142 22372 19180
rect 21980 19124 22036 19134
rect 21980 19030 22036 19068
rect 21588 17948 21700 18004
rect 21756 18338 21812 18350
rect 21756 18286 21758 18338
rect 21810 18286 21812 18338
rect 21532 17938 21588 17948
rect 20860 17836 21028 17892
rect 20524 17668 20580 17678
rect 20524 17574 20580 17612
rect 20860 17668 20916 17836
rect 21196 17724 21588 17780
rect 21196 17668 21252 17724
rect 20860 17666 21028 17668
rect 20860 17614 20862 17666
rect 20914 17614 21028 17666
rect 20860 17612 21028 17614
rect 20860 17602 20916 17612
rect 20524 17444 20580 17454
rect 20412 17442 20580 17444
rect 20412 17390 20526 17442
rect 20578 17390 20580 17442
rect 20412 17388 20580 17390
rect 20524 17378 20580 17388
rect 20300 16370 20356 16380
rect 20636 16324 20692 16334
rect 19964 16212 20020 16222
rect 19964 16118 20020 16156
rect 19740 16100 19796 16110
rect 19628 16098 19796 16100
rect 19628 16046 19742 16098
rect 19794 16046 19796 16098
rect 19628 16044 19796 16046
rect 19068 16006 19124 16044
rect 19404 15874 19460 15886
rect 19404 15822 19406 15874
rect 19458 15822 19460 15874
rect 18508 15092 18676 15148
rect 18844 15148 19012 15204
rect 19068 15764 19124 15774
rect 19068 15538 19124 15708
rect 19404 15652 19460 15822
rect 19740 15876 19796 16044
rect 20076 16100 20132 16110
rect 20636 16100 20692 16268
rect 20748 16100 20804 16110
rect 20636 16098 20804 16100
rect 20636 16046 20750 16098
rect 20802 16046 20804 16098
rect 20636 16044 20804 16046
rect 20076 16006 20132 16044
rect 20748 16034 20804 16044
rect 20524 15876 20580 15886
rect 19740 15820 20244 15876
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19068 15486 19070 15538
rect 19122 15486 19124 15538
rect 18172 14308 18228 14318
rect 17948 14252 18172 14308
rect 17164 13972 17220 14252
rect 18172 14214 18228 14252
rect 17500 13972 17556 13982
rect 17164 13916 17500 13972
rect 17500 13878 17556 13916
rect 18060 13636 18116 13646
rect 18060 13188 18116 13580
rect 17836 13074 17892 13086
rect 17836 13022 17838 13074
rect 17890 13022 17892 13074
rect 16716 12338 16772 12348
rect 17500 12404 17556 12414
rect 17500 12310 17556 12348
rect 16828 12068 16884 12078
rect 16604 12012 16828 12068
rect 16828 11974 16884 12012
rect 17612 12068 17668 12078
rect 16156 11506 16212 11518
rect 16156 11454 16158 11506
rect 16210 11454 16212 11506
rect 15260 10836 15316 10846
rect 15260 10742 15316 10780
rect 13804 10724 13860 10734
rect 13804 10630 13860 10668
rect 15372 10722 15428 10892
rect 15820 11396 15876 11406
rect 15820 10836 15876 11340
rect 15820 10742 15876 10780
rect 15372 10670 15374 10722
rect 15426 10670 15428 10722
rect 15372 10658 15428 10670
rect 14028 10612 14084 10622
rect 14476 10612 14532 10622
rect 15036 10612 15092 10622
rect 14028 10610 14420 10612
rect 14028 10558 14030 10610
rect 14082 10558 14420 10610
rect 14028 10556 14420 10558
rect 14028 10546 14084 10556
rect 13916 10498 13972 10510
rect 13916 10446 13918 10498
rect 13970 10446 13972 10498
rect 13916 10052 13972 10446
rect 13916 9996 14308 10052
rect 14252 9938 14308 9996
rect 14252 9886 14254 9938
rect 14306 9886 14308 9938
rect 14252 9874 14308 9886
rect 14364 9268 14420 10556
rect 14476 10610 15092 10612
rect 14476 10558 14478 10610
rect 14530 10558 15038 10610
rect 15090 10558 15092 10610
rect 14476 10556 15092 10558
rect 14476 10546 14532 10556
rect 15036 10546 15092 10556
rect 16156 9940 16212 11454
rect 16156 9874 16212 9884
rect 16380 9938 16436 9950
rect 16380 9886 16382 9938
rect 16434 9886 16436 9938
rect 14028 9154 14084 9166
rect 14028 9102 14030 9154
rect 14082 9102 14084 9154
rect 13804 8932 13860 8942
rect 13692 8876 13804 8932
rect 13804 8866 13860 8876
rect 14028 8370 14084 9102
rect 14140 9042 14196 9054
rect 14140 8990 14142 9042
rect 14194 8990 14196 9042
rect 14140 8708 14196 8990
rect 14140 8642 14196 8652
rect 14364 8428 14420 9212
rect 15820 9268 15876 9278
rect 15820 9174 15876 9212
rect 16380 9156 16436 9886
rect 15932 9100 16436 9156
rect 17500 9716 17556 9726
rect 14924 9042 14980 9054
rect 14924 8990 14926 9042
rect 14978 8990 14980 9042
rect 14924 8708 14980 8990
rect 15260 9044 15316 9054
rect 15260 8950 15316 8988
rect 15932 8930 15988 9100
rect 15932 8878 15934 8930
rect 15986 8878 15988 8930
rect 15596 8820 15652 8830
rect 15596 8726 15652 8764
rect 14924 8642 14980 8652
rect 14028 8318 14030 8370
rect 14082 8318 14084 8370
rect 14028 8306 14084 8318
rect 14140 8372 14420 8428
rect 13692 8260 13748 8270
rect 13692 8166 13748 8204
rect 14140 8258 14196 8372
rect 14140 8206 14142 8258
rect 14194 8206 14196 8258
rect 14140 8194 14196 8206
rect 12124 8036 12180 8046
rect 12124 7942 12180 7980
rect 12348 8036 12404 8046
rect 11228 7474 11732 7476
rect 11228 7422 11230 7474
rect 11282 7422 11732 7474
rect 11228 7420 11732 7422
rect 10780 7410 10836 7420
rect 9324 6638 9326 6690
rect 9378 6638 9380 6690
rect 9324 6626 9380 6638
rect 11228 6692 11284 7420
rect 11228 6626 11284 6636
rect 12124 6916 12180 6926
rect 11788 6468 11844 6478
rect 11788 6374 11844 6412
rect 8876 6066 8932 6076
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 12124 4338 12180 6860
rect 12348 6690 12404 7980
rect 13468 7028 13524 8092
rect 14364 8146 14420 8158
rect 14364 8094 14366 8146
rect 14418 8094 14420 8146
rect 13916 8036 13972 8046
rect 13916 8034 14084 8036
rect 13916 7982 13918 8034
rect 13970 7982 14084 8034
rect 13916 7980 14084 7982
rect 13916 7970 13972 7980
rect 13692 7700 13748 7710
rect 13692 7698 13860 7700
rect 13692 7646 13694 7698
rect 13746 7646 13860 7698
rect 13692 7644 13860 7646
rect 13692 7634 13748 7644
rect 13356 6972 13524 7028
rect 13356 6916 13412 6972
rect 13244 6860 13412 6916
rect 12684 6804 12740 6814
rect 12348 6638 12350 6690
rect 12402 6638 12404 6690
rect 12348 6626 12404 6638
rect 12572 6692 12628 6702
rect 12572 6598 12628 6636
rect 12684 6690 12740 6748
rect 12684 6638 12686 6690
rect 12738 6638 12740 6690
rect 12684 6626 12740 6638
rect 12236 6468 12292 6478
rect 12236 6130 12292 6412
rect 12236 6078 12238 6130
rect 12290 6078 12292 6130
rect 12236 6066 12292 6078
rect 13132 6132 13188 6142
rect 13132 6038 13188 6076
rect 12460 5908 12516 5918
rect 12348 5906 12516 5908
rect 12348 5854 12462 5906
rect 12514 5854 12516 5906
rect 12348 5852 12516 5854
rect 12348 5346 12404 5852
rect 12460 5842 12516 5852
rect 12348 5294 12350 5346
rect 12402 5294 12404 5346
rect 12348 5282 12404 5294
rect 12460 5684 12516 5694
rect 13244 5684 13300 6860
rect 13468 6804 13524 6814
rect 13356 6748 13468 6804
rect 13356 5906 13412 6748
rect 13468 6738 13524 6748
rect 13804 6578 13860 7644
rect 14028 7362 14084 7980
rect 14028 7310 14030 7362
rect 14082 7310 14084 7362
rect 14028 6804 14084 7310
rect 14028 6738 14084 6748
rect 13804 6526 13806 6578
rect 13858 6526 13860 6578
rect 13804 6514 13860 6526
rect 14140 6578 14196 6590
rect 14140 6526 14142 6578
rect 14194 6526 14196 6578
rect 13356 5854 13358 5906
rect 13410 5854 13412 5906
rect 13356 5842 13412 5854
rect 13916 6468 13972 6478
rect 13916 5906 13972 6412
rect 13916 5854 13918 5906
rect 13970 5854 13972 5906
rect 13916 5842 13972 5854
rect 13356 5684 13412 5694
rect 13244 5628 13356 5684
rect 12124 4286 12126 4338
rect 12178 4286 12180 4338
rect 12124 4274 12180 4286
rect 12460 4338 12516 5628
rect 13356 5618 13412 5628
rect 14140 5346 14196 6526
rect 14364 6020 14420 8094
rect 15820 8148 15876 8158
rect 15820 8054 15876 8092
rect 15932 7812 15988 8878
rect 16044 8932 16100 8942
rect 16044 8258 16100 8876
rect 16044 8206 16046 8258
rect 16098 8206 16100 8258
rect 16044 8194 16100 8206
rect 17052 8258 17108 8270
rect 17052 8206 17054 8258
rect 17106 8206 17108 8258
rect 17052 8148 17108 8206
rect 17052 8082 17108 8092
rect 17388 8258 17444 8270
rect 17388 8206 17390 8258
rect 17442 8206 17444 8258
rect 15932 7746 15988 7756
rect 17388 8036 17444 8206
rect 16828 7476 16884 7486
rect 16828 7382 16884 7420
rect 16716 7364 16772 7374
rect 16716 6916 16772 7308
rect 16828 6916 16884 6926
rect 16772 6914 16884 6916
rect 16772 6862 16830 6914
rect 16882 6862 16884 6914
rect 16772 6860 16884 6862
rect 16716 6822 16772 6860
rect 16828 6850 16884 6860
rect 14364 5954 14420 5964
rect 14476 6578 14532 6590
rect 14476 6526 14478 6578
rect 14530 6526 14532 6578
rect 14140 5294 14142 5346
rect 14194 5294 14196 5346
rect 14140 5282 14196 5294
rect 12572 5236 12628 5246
rect 12572 5142 12628 5180
rect 14252 5236 14308 5246
rect 12460 4286 12462 4338
rect 12514 4286 12516 4338
rect 12460 4274 12516 4286
rect 12684 5122 12740 5134
rect 12684 5070 12686 5122
rect 12738 5070 12740 5122
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 12684 3556 12740 5070
rect 14252 3666 14308 5180
rect 14476 3778 14532 6526
rect 15260 6580 15316 6590
rect 15260 6578 15428 6580
rect 15260 6526 15262 6578
rect 15314 6526 15428 6578
rect 15260 6524 15428 6526
rect 15260 6514 15316 6524
rect 14812 6466 14868 6478
rect 14812 6414 14814 6466
rect 14866 6414 14868 6466
rect 14812 4562 14868 6414
rect 15148 6466 15204 6478
rect 15148 6414 15150 6466
rect 15202 6414 15204 6466
rect 15148 5684 15204 6414
rect 15148 5618 15204 5628
rect 14924 5236 14980 5246
rect 14924 5122 14980 5180
rect 14924 5070 14926 5122
rect 14978 5070 14980 5122
rect 14924 5058 14980 5070
rect 14812 4510 14814 4562
rect 14866 4510 14868 4562
rect 14812 4498 14868 4510
rect 15372 4226 15428 6524
rect 16604 6578 16660 6590
rect 16604 6526 16606 6578
rect 16658 6526 16660 6578
rect 16492 6468 16548 6478
rect 16492 6374 16548 6412
rect 16380 6132 16436 6142
rect 16380 6130 16548 6132
rect 16380 6078 16382 6130
rect 16434 6078 16548 6130
rect 16380 6076 16548 6078
rect 16380 6066 16436 6076
rect 15708 5236 15764 5246
rect 15708 5122 15764 5180
rect 15708 5070 15710 5122
rect 15762 5070 15764 5122
rect 15708 5058 15764 5070
rect 16380 5124 16436 5134
rect 16380 4788 16436 5068
rect 16380 4722 16436 4732
rect 16492 4562 16548 6076
rect 16604 5796 16660 6526
rect 17388 6468 17444 7980
rect 17500 7586 17556 9660
rect 17612 8258 17668 12012
rect 17836 11954 17892 13022
rect 18060 12962 18116 13132
rect 18060 12910 18062 12962
rect 18114 12910 18116 12962
rect 18060 12290 18116 12910
rect 18396 12962 18452 12974
rect 18396 12910 18398 12962
rect 18450 12910 18452 12962
rect 18284 12738 18340 12750
rect 18284 12686 18286 12738
rect 18338 12686 18340 12738
rect 18284 12404 18340 12686
rect 18396 12516 18452 12910
rect 18508 12740 18564 15092
rect 18844 14756 18900 15148
rect 19068 14868 19124 15486
rect 18844 14690 18900 14700
rect 18956 14812 19124 14868
rect 19180 15596 19684 15652
rect 19836 15642 20100 15652
rect 18732 14532 18788 14542
rect 18956 14532 19012 14812
rect 18732 14530 19012 14532
rect 18732 14478 18734 14530
rect 18786 14478 19012 14530
rect 18732 14476 19012 14478
rect 19068 14644 19124 14654
rect 18732 14466 18788 14476
rect 18508 12674 18564 12684
rect 18620 14308 18676 14318
rect 18396 12460 18564 12516
rect 18060 12238 18062 12290
rect 18114 12238 18116 12290
rect 18060 12226 18116 12238
rect 18172 12348 18340 12404
rect 17836 11902 17838 11954
rect 17890 11902 17892 11954
rect 17836 9940 17892 11902
rect 18172 11508 18228 12348
rect 18396 12292 18452 12302
rect 18396 12198 18452 12236
rect 18284 11508 18340 11518
rect 18172 11506 18340 11508
rect 18172 11454 18286 11506
rect 18338 11454 18340 11506
rect 18172 11452 18340 11454
rect 18284 11442 18340 11452
rect 18396 10498 18452 10510
rect 18396 10446 18398 10498
rect 18450 10446 18452 10498
rect 17948 9940 18004 9950
rect 17836 9938 18004 9940
rect 17836 9886 17950 9938
rect 18002 9886 18004 9938
rect 17836 9884 18004 9886
rect 18396 9940 18452 10446
rect 18508 10052 18564 12460
rect 18620 12404 18676 14252
rect 18844 14308 18900 14318
rect 18844 14214 18900 14252
rect 18956 14306 19012 14318
rect 18956 14254 18958 14306
rect 19010 14254 19012 14306
rect 18956 14084 19012 14254
rect 18732 14028 19012 14084
rect 18732 13970 18788 14028
rect 18732 13918 18734 13970
rect 18786 13918 18788 13970
rect 18732 13906 18788 13918
rect 18956 13858 19012 13870
rect 18956 13806 18958 13858
rect 19010 13806 19012 13858
rect 18956 13748 19012 13806
rect 19068 13858 19124 14588
rect 19180 14530 19236 15596
rect 19628 15540 19684 15596
rect 19628 15484 20020 15540
rect 19404 15428 19460 15438
rect 19180 14478 19182 14530
rect 19234 14478 19236 14530
rect 19180 14466 19236 14478
rect 19292 15314 19348 15326
rect 19292 15262 19294 15314
rect 19346 15262 19348 15314
rect 19068 13806 19070 13858
rect 19122 13806 19124 13858
rect 19068 13794 19124 13806
rect 18956 13682 19012 13692
rect 19292 13748 19348 15262
rect 19292 13682 19348 13692
rect 19404 13970 19460 15372
rect 19516 15426 19572 15438
rect 19516 15374 19518 15426
rect 19570 15374 19572 15426
rect 19516 15316 19572 15374
rect 19516 15250 19572 15260
rect 19628 15314 19684 15326
rect 19628 15262 19630 15314
rect 19682 15262 19684 15314
rect 19628 15204 19684 15262
rect 19964 15314 20020 15484
rect 19964 15262 19966 15314
rect 20018 15262 20020 15314
rect 19964 15250 20020 15262
rect 19628 15138 19684 15148
rect 19516 14756 19572 14766
rect 19572 14700 19684 14756
rect 19516 14690 19572 14700
rect 19404 13918 19406 13970
rect 19458 13918 19460 13970
rect 19404 13524 19460 13918
rect 19180 13468 19460 13524
rect 19516 14530 19572 14542
rect 19516 14478 19518 14530
rect 19570 14478 19572 14530
rect 19068 13074 19124 13086
rect 19068 13022 19070 13074
rect 19122 13022 19124 13074
rect 18732 12964 18788 12974
rect 19068 12964 19124 13022
rect 18732 12962 19124 12964
rect 18732 12910 18734 12962
rect 18786 12910 19124 12962
rect 18732 12908 19124 12910
rect 19180 13076 19236 13468
rect 19404 13188 19460 13198
rect 19516 13188 19572 14478
rect 19460 13132 19572 13188
rect 19404 13094 19460 13132
rect 18732 12898 18788 12908
rect 19180 12850 19236 13020
rect 19180 12798 19182 12850
rect 19234 12798 19236 12850
rect 19180 12786 19236 12798
rect 19404 12404 19460 12414
rect 18620 12402 19460 12404
rect 18620 12350 19406 12402
rect 19458 12350 19460 12402
rect 18620 12348 19460 12350
rect 19404 12338 19460 12348
rect 19180 12178 19236 12190
rect 19180 12126 19182 12178
rect 19234 12126 19236 12178
rect 19068 11620 19124 11630
rect 19068 11394 19124 11564
rect 19068 11342 19070 11394
rect 19122 11342 19124 11394
rect 18732 10164 18788 10174
rect 18732 10052 18788 10108
rect 18508 10050 18788 10052
rect 18508 9998 18734 10050
rect 18786 9998 18788 10050
rect 18508 9996 18788 9998
rect 18732 9986 18788 9996
rect 18844 9940 18900 9950
rect 18396 9884 18676 9940
rect 17948 9874 18004 9884
rect 17724 9826 17780 9838
rect 17724 9774 17726 9826
rect 17778 9774 17780 9826
rect 17724 8708 17780 9774
rect 18396 9716 18452 9726
rect 18396 9622 18452 9660
rect 18620 9716 18676 9884
rect 18844 9846 18900 9884
rect 18620 9380 18676 9660
rect 18620 9324 18900 9380
rect 18172 9042 18228 9054
rect 18172 8990 18174 9042
rect 18226 8990 18228 9042
rect 18172 8932 18228 8990
rect 18284 8988 18564 9044
rect 18284 8932 18340 8988
rect 18172 8876 18340 8932
rect 18396 8818 18452 8830
rect 18396 8766 18398 8818
rect 18450 8766 18452 8818
rect 17724 8652 18116 8708
rect 17612 8206 17614 8258
rect 17666 8206 17668 8258
rect 17612 7924 17668 8206
rect 17612 7858 17668 7868
rect 17948 8482 18004 8494
rect 17948 8430 17950 8482
rect 18002 8430 18004 8482
rect 17500 7534 17502 7586
rect 17554 7534 17556 7586
rect 17500 7522 17556 7534
rect 17948 7474 18004 8430
rect 17948 7422 17950 7474
rect 18002 7422 18004 7474
rect 17948 7410 18004 7422
rect 18060 6692 18116 8652
rect 18396 7476 18452 8766
rect 18508 8370 18564 8988
rect 18508 8318 18510 8370
rect 18562 8318 18564 8370
rect 18508 8306 18564 8318
rect 18732 9042 18788 9054
rect 18732 8990 18734 9042
rect 18786 8990 18788 9042
rect 18732 8372 18788 8990
rect 18732 8306 18788 8316
rect 18844 8258 18900 9324
rect 19068 8932 19124 11342
rect 19068 8866 19124 8876
rect 18844 8206 18846 8258
rect 18898 8206 18900 8258
rect 18844 8194 18900 8206
rect 18956 8820 19012 8830
rect 18508 8034 18564 8046
rect 18508 7982 18510 8034
rect 18562 7982 18564 8034
rect 18508 7924 18564 7982
rect 18620 8036 18676 8046
rect 18620 7942 18676 7980
rect 18508 7858 18564 7868
rect 18844 7698 18900 7710
rect 18844 7646 18846 7698
rect 18898 7646 18900 7698
rect 18508 7476 18564 7486
rect 18396 7474 18564 7476
rect 18396 7422 18510 7474
rect 18562 7422 18564 7474
rect 18396 7420 18564 7422
rect 18508 7410 18564 7420
rect 18844 7364 18900 7646
rect 18956 7586 19012 8764
rect 18956 7534 18958 7586
rect 19010 7534 19012 7586
rect 18956 7522 19012 7534
rect 19068 8146 19124 8158
rect 19068 8094 19070 8146
rect 19122 8094 19124 8146
rect 19068 7588 19124 8094
rect 19068 7522 19124 7532
rect 19180 7364 19236 12126
rect 19628 11620 19684 14700
rect 20076 14644 20132 14654
rect 20076 14530 20132 14588
rect 20076 14478 20078 14530
rect 20130 14478 20132 14530
rect 20076 14466 20132 14478
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13972 20244 15820
rect 20524 15782 20580 15820
rect 20636 15874 20692 15886
rect 20636 15822 20638 15874
rect 20690 15822 20692 15874
rect 20636 15204 20692 15822
rect 20860 15428 20916 15438
rect 20748 15372 20860 15428
rect 20748 15314 20804 15372
rect 20860 15362 20916 15372
rect 20748 15262 20750 15314
rect 20802 15262 20804 15314
rect 20748 15250 20804 15262
rect 20972 15148 21028 17612
rect 20524 14532 20580 14542
rect 20636 14532 20692 15148
rect 20524 14530 20692 14532
rect 20524 14478 20526 14530
rect 20578 14478 20692 14530
rect 20524 14476 20692 14478
rect 20748 15092 21028 15148
rect 20524 14466 20580 14476
rect 20748 14420 20804 15092
rect 21196 14756 21252 17612
rect 21532 17666 21588 17724
rect 21532 17614 21534 17666
rect 21586 17614 21588 17666
rect 21532 17602 21588 17614
rect 21308 17556 21364 17566
rect 21308 17462 21364 17500
rect 21420 17442 21476 17454
rect 21420 17390 21422 17442
rect 21474 17390 21476 17442
rect 21308 16212 21364 16222
rect 21308 16098 21364 16156
rect 21308 16046 21310 16098
rect 21362 16046 21364 16098
rect 21308 16034 21364 16046
rect 21420 15428 21476 17390
rect 21644 16996 21700 17006
rect 21644 16098 21700 16940
rect 21756 16884 21812 18286
rect 22428 18228 22484 18238
rect 22316 17780 22372 17790
rect 21868 17778 22372 17780
rect 21868 17726 22318 17778
rect 22370 17726 22372 17778
rect 21868 17724 22372 17726
rect 21868 17666 21924 17724
rect 22316 17714 22372 17724
rect 21868 17614 21870 17666
rect 21922 17614 21924 17666
rect 21868 17602 21924 17614
rect 22204 17556 22260 17566
rect 21756 16828 21924 16884
rect 21756 16548 21812 16558
rect 21868 16548 21924 16828
rect 21980 16548 22036 16558
rect 21868 16492 21980 16548
rect 21756 16210 21812 16492
rect 21980 16482 22036 16492
rect 21756 16158 21758 16210
rect 21810 16158 21812 16210
rect 21756 16146 21812 16158
rect 21644 16046 21646 16098
rect 21698 16046 21700 16098
rect 21644 16034 21700 16046
rect 21868 16100 21924 16110
rect 22204 16100 22260 17500
rect 22428 17554 22484 18172
rect 22428 17502 22430 17554
rect 22482 17502 22484 17554
rect 22428 17490 22484 17502
rect 21924 16044 22260 16100
rect 21868 16006 21924 16044
rect 21420 15362 21476 15372
rect 21532 15988 21588 15998
rect 21532 15316 21588 15932
rect 22204 15986 22260 16044
rect 22204 15934 22206 15986
rect 22258 15934 22260 15986
rect 22204 15922 22260 15934
rect 22316 16772 22372 16782
rect 22316 15876 22372 16716
rect 22428 16660 22484 16670
rect 22540 16660 22596 22092
rect 22876 21474 22932 22316
rect 23772 22370 23828 24444
rect 24108 23938 24164 24780
rect 24780 24834 25284 24836
rect 24780 24782 25230 24834
rect 25282 24782 25284 24834
rect 24780 24780 25284 24782
rect 24780 24050 24836 24780
rect 25228 24770 25284 24780
rect 24780 23998 24782 24050
rect 24834 23998 24836 24050
rect 24780 23986 24836 23998
rect 24108 23886 24110 23938
rect 24162 23886 24164 23938
rect 24108 23874 24164 23886
rect 23996 23156 24052 23166
rect 23996 22482 24052 23100
rect 23996 22430 23998 22482
rect 24050 22430 24052 22482
rect 23996 22418 24052 22430
rect 25340 23154 25396 29148
rect 25564 28644 25620 28654
rect 25564 28550 25620 28588
rect 26012 28084 26068 28094
rect 26012 27990 26068 28028
rect 25900 27972 25956 27982
rect 25900 27878 25956 27916
rect 25564 27860 25620 27870
rect 25564 27858 25844 27860
rect 25564 27806 25566 27858
rect 25618 27806 25844 27858
rect 25564 27804 25844 27806
rect 25564 27794 25620 27804
rect 25788 26516 25844 27804
rect 26012 27634 26068 27646
rect 26012 27582 26014 27634
rect 26066 27582 26068 27634
rect 26012 26964 26068 27582
rect 26012 26898 26068 26908
rect 26236 27300 26292 27310
rect 25900 26516 25956 26526
rect 25788 26514 25956 26516
rect 25788 26462 25902 26514
rect 25954 26462 25956 26514
rect 25788 26460 25956 26462
rect 25900 26450 25956 26460
rect 26236 26290 26292 27244
rect 26460 27076 26516 29374
rect 27020 29428 27076 29438
rect 27020 29334 27076 29372
rect 26908 28644 26964 28654
rect 26572 27860 26628 27870
rect 26572 27766 26628 27804
rect 26908 27858 26964 28588
rect 26908 27806 26910 27858
rect 26962 27806 26964 27858
rect 26908 27794 26964 27806
rect 26572 27076 26628 27086
rect 26460 27020 26572 27076
rect 26236 26238 26238 26290
rect 26290 26238 26292 26290
rect 26236 26226 26292 26238
rect 26572 26402 26628 27020
rect 27020 26964 27076 26974
rect 27020 26870 27076 26908
rect 27132 26628 27188 29708
rect 27244 27972 27300 29934
rect 27356 29426 27412 30940
rect 27580 30882 27636 30894
rect 27580 30830 27582 30882
rect 27634 30830 27636 30882
rect 27468 30210 27524 30222
rect 27468 30158 27470 30210
rect 27522 30158 27524 30210
rect 27468 30100 27524 30158
rect 27468 30034 27524 30044
rect 27580 29764 27636 30830
rect 28028 30770 28084 31726
rect 30268 31106 30324 31118
rect 30268 31054 30270 31106
rect 30322 31054 30324 31106
rect 28028 30718 28030 30770
rect 28082 30718 28084 30770
rect 28028 30706 28084 30718
rect 29932 30996 29988 31006
rect 29596 30212 29652 30222
rect 28140 30098 28196 30110
rect 28140 30046 28142 30098
rect 28194 30046 28196 30098
rect 27804 29988 27860 29998
rect 27804 29894 27860 29932
rect 28028 29986 28084 29998
rect 28028 29934 28030 29986
rect 28082 29934 28084 29986
rect 27580 29698 27636 29708
rect 27356 29374 27358 29426
rect 27410 29374 27412 29426
rect 27356 29362 27412 29374
rect 27580 29538 27636 29550
rect 27580 29486 27582 29538
rect 27634 29486 27636 29538
rect 27580 28196 27636 29486
rect 27916 29538 27972 29550
rect 27916 29486 27918 29538
rect 27970 29486 27972 29538
rect 27916 29428 27972 29486
rect 27244 27906 27300 27916
rect 27356 28140 27636 28196
rect 27804 28532 27860 28542
rect 27356 27858 27412 28140
rect 27356 27806 27358 27858
rect 27410 27806 27412 27858
rect 27356 27076 27412 27806
rect 27468 27970 27524 27982
rect 27468 27918 27470 27970
rect 27522 27918 27524 27970
rect 27468 27748 27524 27918
rect 27524 27692 27748 27748
rect 27468 27682 27524 27692
rect 27356 27010 27412 27020
rect 26572 26350 26574 26402
rect 26626 26350 26628 26402
rect 25676 25508 25732 25546
rect 25676 25442 25732 25452
rect 26348 25508 26404 25518
rect 26348 25414 26404 25452
rect 25452 25282 25508 25294
rect 25452 25230 25454 25282
rect 25506 25230 25508 25282
rect 25452 23716 25508 25230
rect 25564 24724 25620 24734
rect 26124 24724 26180 24734
rect 25564 24722 26180 24724
rect 25564 24670 25566 24722
rect 25618 24670 26126 24722
rect 26178 24670 26180 24722
rect 25564 24668 26180 24670
rect 25564 24658 25620 24668
rect 26124 24658 26180 24668
rect 26460 24612 26516 24622
rect 26460 24518 26516 24556
rect 25452 23650 25508 23660
rect 25340 23102 25342 23154
rect 25394 23102 25396 23154
rect 23772 22318 23774 22370
rect 23826 22318 23828 22370
rect 23772 22306 23828 22318
rect 24108 22258 24164 22270
rect 24108 22206 24110 22258
rect 24162 22206 24164 22258
rect 23100 22148 23156 22158
rect 23100 22054 23156 22092
rect 22876 21422 22878 21474
rect 22930 21422 22932 21474
rect 22876 21410 22932 21422
rect 22764 20804 22820 20814
rect 22652 20692 22708 20702
rect 22652 20598 22708 20636
rect 22764 19906 22820 20748
rect 23212 20692 23268 20702
rect 23212 20598 23268 20636
rect 22764 19854 22766 19906
rect 22818 19854 22820 19906
rect 22764 19842 22820 19854
rect 24108 19236 24164 22206
rect 25340 21586 25396 23102
rect 26012 23044 26068 23054
rect 25788 23042 26068 23044
rect 25788 22990 26014 23042
rect 26066 22990 26068 23042
rect 25788 22988 26068 22990
rect 25564 22370 25620 22382
rect 25564 22318 25566 22370
rect 25618 22318 25620 22370
rect 25564 22036 25620 22318
rect 25788 22258 25844 22988
rect 26012 22978 26068 22988
rect 25788 22206 25790 22258
rect 25842 22206 25844 22258
rect 25788 22194 25844 22206
rect 26348 22146 26404 22158
rect 26348 22094 26350 22146
rect 26402 22094 26404 22146
rect 26348 22036 26404 22094
rect 25564 21980 26404 22036
rect 25340 21534 25342 21586
rect 25394 21534 25396 21586
rect 25340 21522 25396 21534
rect 26348 21812 26404 21822
rect 26012 21476 26068 21486
rect 26012 21474 26180 21476
rect 26012 21422 26014 21474
rect 26066 21422 26180 21474
rect 26012 21420 26180 21422
rect 26012 21410 26068 21420
rect 25340 20804 25396 20814
rect 26012 20804 26068 20814
rect 25340 20802 26068 20804
rect 25340 20750 25342 20802
rect 25394 20750 26014 20802
rect 26066 20750 26068 20802
rect 25340 20748 26068 20750
rect 25340 20738 25396 20748
rect 26012 20738 26068 20748
rect 25564 20580 25620 20590
rect 26124 20580 26180 21420
rect 26348 21026 26404 21756
rect 26348 20974 26350 21026
rect 26402 20974 26404 21026
rect 26348 20962 26404 20974
rect 25564 20578 26180 20580
rect 25564 20526 25566 20578
rect 25618 20526 26180 20578
rect 25564 20524 26180 20526
rect 25564 20514 25620 20524
rect 25900 20244 25956 20254
rect 25900 20130 25956 20188
rect 26572 20242 26628 26350
rect 26908 26572 27188 26628
rect 26908 24276 26964 26572
rect 27020 26402 27076 26414
rect 27020 26350 27022 26402
rect 27074 26350 27076 26402
rect 27020 26292 27076 26350
rect 27020 26236 27524 26292
rect 27468 26180 27524 26236
rect 27580 26180 27636 26190
rect 27468 26178 27636 26180
rect 27468 26126 27582 26178
rect 27634 26126 27636 26178
rect 27468 26124 27636 26126
rect 27244 24836 27300 24874
rect 27244 24770 27300 24780
rect 27132 24722 27188 24734
rect 27132 24670 27134 24722
rect 27186 24670 27188 24722
rect 26908 24210 26964 24220
rect 27020 24612 27076 24622
rect 26908 24052 26964 24062
rect 27020 24052 27076 24556
rect 26908 24050 27076 24052
rect 26908 23998 26910 24050
rect 26962 23998 27076 24050
rect 26908 23996 27076 23998
rect 26908 23986 26964 23996
rect 27132 22484 27188 24670
rect 26684 22370 26740 22382
rect 26684 22318 26686 22370
rect 26738 22318 26740 22370
rect 26684 22148 26740 22318
rect 27132 22370 27188 22428
rect 27132 22318 27134 22370
rect 27186 22318 27188 22370
rect 27132 22306 27188 22318
rect 27244 24276 27300 24286
rect 26908 22260 26964 22270
rect 27244 22260 27300 24220
rect 27468 22260 27524 22270
rect 26964 22204 27076 22260
rect 27244 22258 27524 22260
rect 27244 22206 27470 22258
rect 27522 22206 27524 22258
rect 27244 22204 27524 22206
rect 26908 22194 26964 22204
rect 26684 22082 26740 22092
rect 26572 20190 26574 20242
rect 26626 20190 26628 20242
rect 26572 20178 26628 20190
rect 26796 21700 26852 21710
rect 26796 20244 26852 21644
rect 26908 20692 26964 20702
rect 26908 20598 26964 20636
rect 27020 20468 27076 22204
rect 27468 22036 27524 22204
rect 27468 21970 27524 21980
rect 25900 20078 25902 20130
rect 25954 20078 25956 20130
rect 25788 20018 25844 20030
rect 25788 19966 25790 20018
rect 25842 19966 25844 20018
rect 24220 19236 24276 19246
rect 24108 19180 24220 19236
rect 24108 18562 24164 18574
rect 24108 18510 24110 18562
rect 24162 18510 24164 18562
rect 23884 18340 23940 18350
rect 22484 16604 22596 16660
rect 22652 18228 22708 18238
rect 22428 16594 22484 16604
rect 22652 16436 22708 18172
rect 23436 18228 23492 18238
rect 23436 17778 23492 18172
rect 23436 17726 23438 17778
rect 23490 17726 23492 17778
rect 23436 17714 23492 17726
rect 22988 17554 23044 17566
rect 22988 17502 22990 17554
rect 23042 17502 23044 17554
rect 22876 17442 22932 17454
rect 22876 17390 22878 17442
rect 22930 17390 22932 17442
rect 22876 16996 22932 17390
rect 22876 16882 22932 16940
rect 22876 16830 22878 16882
rect 22930 16830 22932 16882
rect 22876 16818 22932 16830
rect 22988 16772 23044 17502
rect 23884 17108 23940 18284
rect 23996 17668 24052 17678
rect 24108 17668 24164 18510
rect 23996 17666 24164 17668
rect 23996 17614 23998 17666
rect 24050 17614 24164 17666
rect 23996 17612 24164 17614
rect 23996 17602 24052 17612
rect 23436 17106 23940 17108
rect 23436 17054 23886 17106
rect 23938 17054 23940 17106
rect 23436 17052 23940 17054
rect 23436 16994 23492 17052
rect 23884 17042 23940 17052
rect 23436 16942 23438 16994
rect 23490 16942 23492 16994
rect 23436 16930 23492 16942
rect 23996 16884 24052 16894
rect 23996 16790 24052 16828
rect 22988 16706 23044 16716
rect 23100 16770 23156 16782
rect 23100 16718 23102 16770
rect 23154 16718 23156 16770
rect 22316 15428 22372 15820
rect 22316 15362 22372 15372
rect 22428 16380 22708 16436
rect 21532 15148 21588 15260
rect 21420 15092 21588 15148
rect 21308 14756 21364 14766
rect 21196 14754 21364 14756
rect 21196 14702 21310 14754
rect 21362 14702 21364 14754
rect 21196 14700 21364 14702
rect 21308 14690 21364 14700
rect 21420 14642 21476 15092
rect 21420 14590 21422 14642
rect 21474 14590 21476 14642
rect 21420 14578 21476 14590
rect 21868 14642 21924 14654
rect 21868 14590 21870 14642
rect 21922 14590 21924 14642
rect 21644 14530 21700 14542
rect 21644 14478 21646 14530
rect 21698 14478 21700 14530
rect 21644 14420 21700 14478
rect 20748 14418 21700 14420
rect 20748 14366 20750 14418
rect 20802 14366 21700 14418
rect 20748 14364 21700 14366
rect 20748 14354 20804 14364
rect 20076 13916 20244 13972
rect 19852 13636 19908 13646
rect 19852 13542 19908 13580
rect 20076 13188 20132 13916
rect 20300 13860 20356 13870
rect 20300 13766 20356 13804
rect 20412 13748 20468 13786
rect 20412 13682 20468 13692
rect 20860 13748 20916 13758
rect 20860 13654 20916 13692
rect 21868 13412 21924 14590
rect 21980 14306 22036 14318
rect 21980 14254 21982 14306
rect 22034 14254 22036 14306
rect 21980 13972 22036 14254
rect 21980 13906 22036 13916
rect 22204 14308 22260 14318
rect 22204 13748 22260 14252
rect 22204 13682 22260 13692
rect 20076 13122 20132 13132
rect 21756 13356 21924 13412
rect 20188 13076 20244 13086
rect 20188 12982 20244 13020
rect 20636 13076 20692 13086
rect 20636 12982 20692 13020
rect 21644 12850 21700 12862
rect 21644 12798 21646 12850
rect 21698 12798 21700 12850
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19852 12292 19908 12302
rect 19852 12198 19908 12236
rect 21420 12290 21476 12302
rect 21420 12238 21422 12290
rect 21474 12238 21476 12290
rect 19628 11554 19684 11564
rect 21196 11620 21252 11630
rect 20748 11508 20804 11518
rect 20748 11414 20804 11452
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 21196 10610 21252 11564
rect 21196 10558 21198 10610
rect 21250 10558 21252 10610
rect 21196 10546 21252 10558
rect 21420 10724 21476 12238
rect 21644 11620 21700 12798
rect 21756 12404 21812 13356
rect 22428 13300 22484 16380
rect 23100 16324 23156 16718
rect 23884 16660 23940 16670
rect 24108 16660 24164 17612
rect 24220 16772 24276 19180
rect 25228 18562 25284 18574
rect 25228 18510 25230 18562
rect 25282 18510 25284 18562
rect 24444 18452 24500 18462
rect 24444 18450 24612 18452
rect 24444 18398 24446 18450
rect 24498 18398 24612 18450
rect 24444 18396 24612 18398
rect 24444 18386 24500 18396
rect 24220 16706 24276 16716
rect 24556 17556 24612 18396
rect 25228 18116 25284 18510
rect 25788 18564 25844 19966
rect 25788 18498 25844 18508
rect 25452 18452 25508 18462
rect 24668 18060 25284 18116
rect 25340 18450 25508 18452
rect 25340 18398 25454 18450
rect 25506 18398 25508 18450
rect 25340 18396 25508 18398
rect 24668 17778 24724 18060
rect 24668 17726 24670 17778
rect 24722 17726 24724 17778
rect 24668 17714 24724 17726
rect 23100 16258 23156 16268
rect 23772 16658 23940 16660
rect 23772 16606 23886 16658
rect 23938 16606 23940 16658
rect 23772 16604 23940 16606
rect 23436 16210 23492 16222
rect 23436 16158 23438 16210
rect 23490 16158 23492 16210
rect 23100 16100 23156 16110
rect 23100 16006 23156 16044
rect 22540 15874 22596 15886
rect 22540 15822 22542 15874
rect 22594 15822 22596 15874
rect 22540 15652 22596 15822
rect 22540 15586 22596 15596
rect 22876 15204 22932 15242
rect 22876 15138 22932 15148
rect 23324 15092 23380 15102
rect 22988 15090 23380 15092
rect 22988 15038 23326 15090
rect 23378 15038 23380 15090
rect 22988 15036 23380 15038
rect 22652 14532 22708 14542
rect 22652 14438 22708 14476
rect 22876 13748 22932 13758
rect 22988 13748 23044 15036
rect 23324 15026 23380 15036
rect 23324 14420 23380 14430
rect 23100 14418 23380 14420
rect 23100 14366 23326 14418
rect 23378 14366 23380 14418
rect 23100 14364 23380 14366
rect 23100 13970 23156 14364
rect 23324 14354 23380 14364
rect 23100 13918 23102 13970
rect 23154 13918 23156 13970
rect 23100 13906 23156 13918
rect 23436 13972 23492 16158
rect 23660 15202 23716 15214
rect 23660 15150 23662 15202
rect 23714 15150 23716 15202
rect 23660 14308 23716 15150
rect 23772 14644 23828 16604
rect 23884 16594 23940 16604
rect 23996 16604 24164 16660
rect 23884 16100 23940 16110
rect 23884 16006 23940 16044
rect 23772 14578 23828 14588
rect 23660 14242 23716 14252
rect 23436 13906 23492 13916
rect 22876 13746 23044 13748
rect 22876 13694 22878 13746
rect 22930 13694 23044 13746
rect 22876 13692 23044 13694
rect 22876 13682 22932 13692
rect 21868 13244 22484 13300
rect 21868 12850 21924 13244
rect 21868 12798 21870 12850
rect 21922 12798 21924 12850
rect 21868 12786 21924 12798
rect 21980 13074 22036 13086
rect 21980 13022 21982 13074
rect 22034 13022 22036 13074
rect 21756 12310 21812 12348
rect 21756 11620 21812 11630
rect 21644 11564 21756 11620
rect 21756 11526 21812 11564
rect 21532 11508 21588 11518
rect 21532 11282 21588 11452
rect 21532 11230 21534 11282
rect 21586 11230 21588 11282
rect 21532 11218 21588 11230
rect 20524 10500 20580 10510
rect 20524 10498 21140 10500
rect 20524 10446 20526 10498
rect 20578 10446 21140 10498
rect 20524 10444 21140 10446
rect 20524 10434 20580 10444
rect 20972 10276 21028 10286
rect 19516 10164 19572 10174
rect 20636 10164 20692 10174
rect 19572 10108 19684 10164
rect 19516 10098 19572 10108
rect 19628 9268 19684 10108
rect 20524 10108 20636 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19628 9212 20020 9268
rect 19404 9154 19460 9166
rect 19404 9102 19406 9154
rect 19458 9102 19460 9154
rect 18844 7308 19236 7364
rect 19292 8036 19348 8046
rect 19404 8036 19460 9102
rect 19516 9042 19572 9054
rect 19516 8990 19518 9042
rect 19570 8990 19572 9042
rect 19516 8260 19572 8990
rect 19852 9042 19908 9054
rect 19852 8990 19854 9042
rect 19906 8990 19908 9042
rect 19740 8932 19796 8942
rect 19852 8932 19908 8990
rect 19796 8876 19908 8932
rect 19740 8866 19796 8876
rect 19516 8194 19572 8204
rect 19964 8258 20020 9212
rect 20524 9156 20580 10108
rect 20636 10098 20692 10108
rect 20636 9716 20692 9726
rect 20972 9716 21028 10220
rect 21084 10052 21140 10444
rect 21420 10276 21476 10668
rect 21644 11170 21700 11182
rect 21644 11118 21646 11170
rect 21698 11118 21700 11170
rect 21644 10722 21700 11118
rect 21644 10670 21646 10722
rect 21698 10670 21700 10722
rect 21644 10658 21700 10670
rect 21420 10210 21476 10220
rect 21868 10610 21924 10622
rect 21868 10558 21870 10610
rect 21922 10558 21924 10610
rect 21868 10052 21924 10558
rect 21084 9996 21476 10052
rect 21420 9938 21476 9996
rect 21868 9986 21924 9996
rect 21420 9886 21422 9938
rect 21474 9886 21476 9938
rect 21420 9874 21476 9886
rect 21532 9826 21588 9838
rect 21532 9774 21534 9826
rect 21586 9774 21588 9826
rect 21308 9716 21364 9726
rect 20972 9714 21364 9716
rect 20972 9662 21310 9714
rect 21362 9662 21364 9714
rect 20972 9660 21364 9662
rect 20636 9622 20692 9660
rect 21308 9650 21364 9660
rect 20748 9604 20804 9614
rect 20748 9602 21252 9604
rect 20748 9550 20750 9602
rect 20802 9550 21252 9602
rect 20748 9548 21252 9550
rect 20748 9538 20804 9548
rect 21196 9492 21252 9548
rect 21532 9492 21588 9774
rect 21868 9828 21924 9838
rect 21980 9828 22036 13022
rect 22428 13074 22484 13244
rect 22428 13022 22430 13074
rect 22482 13022 22484 13074
rect 22428 13010 22484 13022
rect 22988 13188 23044 13198
rect 22876 12740 22932 12750
rect 22540 12684 22876 12740
rect 22092 12404 22148 12414
rect 22092 12290 22148 12348
rect 22092 12238 22094 12290
rect 22146 12238 22148 12290
rect 22092 12226 22148 12238
rect 22428 12290 22484 12302
rect 22428 12238 22430 12290
rect 22482 12238 22484 12290
rect 22428 11732 22484 12238
rect 22092 11620 22148 11630
rect 22428 11620 22484 11676
rect 22148 11564 22484 11620
rect 22092 11526 22148 11564
rect 22428 11396 22484 11406
rect 22540 11396 22596 12684
rect 22876 12646 22932 12684
rect 22988 12404 23044 13132
rect 22988 12310 23044 12348
rect 23660 12404 23716 12414
rect 23660 12310 23716 12348
rect 22876 12066 22932 12078
rect 22876 12014 22878 12066
rect 22930 12014 22932 12066
rect 22764 11954 22820 11966
rect 22764 11902 22766 11954
rect 22818 11902 22820 11954
rect 22764 11732 22820 11902
rect 22764 11666 22820 11676
rect 22764 11396 22820 11406
rect 22484 11340 22596 11396
rect 22652 11340 22764 11396
rect 22428 11302 22484 11340
rect 22204 11172 22260 11182
rect 22204 11078 22260 11116
rect 22204 10724 22260 10734
rect 22204 10630 22260 10668
rect 22092 10498 22148 10510
rect 22092 10446 22094 10498
rect 22146 10446 22148 10498
rect 22092 10164 22148 10446
rect 22092 10098 22148 10108
rect 21868 9826 22036 9828
rect 21868 9774 21870 9826
rect 21922 9774 22036 9826
rect 21868 9772 22036 9774
rect 22428 10052 22484 10062
rect 21868 9762 21924 9772
rect 21196 9436 21812 9492
rect 20636 9156 20692 9166
rect 20524 9154 20692 9156
rect 20524 9102 20638 9154
rect 20690 9102 20692 9154
rect 20524 9100 20692 9102
rect 20636 9090 20692 9100
rect 20412 8820 20468 8830
rect 20300 8372 20356 8382
rect 20300 8278 20356 8316
rect 19964 8206 19966 8258
rect 20018 8206 20020 8258
rect 19964 8194 20020 8206
rect 20412 8258 20468 8764
rect 20412 8206 20414 8258
rect 20466 8206 20468 8258
rect 20412 8194 20468 8206
rect 21308 8596 21364 8606
rect 21308 8258 21364 8540
rect 21308 8206 21310 8258
rect 21362 8206 21364 8258
rect 21308 8194 21364 8206
rect 21420 8370 21476 8382
rect 21420 8318 21422 8370
rect 21474 8318 21476 8370
rect 21420 8260 21476 8318
rect 21420 8194 21476 8204
rect 21644 8260 21700 8270
rect 19740 8146 19796 8158
rect 19740 8094 19742 8146
rect 19794 8094 19796 8146
rect 19740 8036 19796 8094
rect 19404 7980 19684 8036
rect 19292 7364 19348 7980
rect 19516 7812 19572 7822
rect 19516 7698 19572 7756
rect 19516 7646 19518 7698
rect 19570 7646 19572 7698
rect 19516 7634 19572 7646
rect 19628 7700 19684 7980
rect 19740 7970 19796 7980
rect 20188 8034 20244 8046
rect 20188 7982 20190 8034
rect 20242 7982 20244 8034
rect 20188 7924 20244 7982
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20188 7858 20244 7868
rect 20748 8036 20804 8046
rect 19836 7802 20100 7812
rect 19740 7700 19796 7710
rect 19628 7698 19796 7700
rect 19628 7646 19742 7698
rect 19794 7646 19796 7698
rect 19628 7644 19796 7646
rect 19740 7634 19796 7644
rect 19292 7298 19348 7308
rect 19628 7474 19684 7486
rect 19628 7422 19630 7474
rect 19682 7422 19684 7474
rect 18396 6804 18452 6814
rect 18060 6626 18116 6636
rect 18284 6748 18396 6804
rect 17388 6402 17444 6412
rect 17612 6466 17668 6478
rect 17612 6414 17614 6466
rect 17666 6414 17668 6466
rect 17612 6244 17668 6414
rect 17612 6188 18228 6244
rect 18172 6130 18228 6188
rect 18172 6078 18174 6130
rect 18226 6078 18228 6130
rect 18172 6066 18228 6078
rect 17724 6020 17780 6030
rect 17724 5926 17780 5964
rect 17836 5908 17892 5918
rect 18284 5908 18340 6748
rect 18396 6738 18452 6748
rect 19628 6804 19684 7422
rect 19852 7474 19908 7486
rect 19852 7422 19854 7474
rect 19906 7422 19908 7474
rect 19852 7364 19908 7422
rect 19852 7298 19908 7308
rect 19964 7476 20020 7486
rect 19628 6738 19684 6748
rect 19964 6690 20020 7420
rect 19964 6638 19966 6690
rect 20018 6638 20020 6690
rect 19964 6626 20020 6638
rect 20300 6692 20356 6702
rect 20300 6598 20356 6636
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 18844 6132 18900 6142
rect 17836 5906 18340 5908
rect 17836 5854 17838 5906
rect 17890 5854 18340 5906
rect 17836 5852 18340 5854
rect 18396 5906 18452 5918
rect 18396 5854 18398 5906
rect 18450 5854 18452 5906
rect 16716 5796 16772 5806
rect 16604 5794 16772 5796
rect 16604 5742 16718 5794
rect 16770 5742 16772 5794
rect 16604 5740 16772 5742
rect 16716 5124 16772 5740
rect 16716 5058 16772 5068
rect 17388 5124 17444 5134
rect 17388 5030 17444 5068
rect 17836 5122 17892 5852
rect 17836 5070 17838 5122
rect 17890 5070 17892 5122
rect 17836 5058 17892 5070
rect 16492 4510 16494 4562
rect 16546 4510 16548 4562
rect 16492 4498 16548 4510
rect 16604 5010 16660 5022
rect 16604 4958 16606 5010
rect 16658 4958 16660 5010
rect 16604 4340 16660 4958
rect 17948 5012 18004 5022
rect 17388 4788 17444 4798
rect 16716 4340 16772 4350
rect 16604 4338 16772 4340
rect 16604 4286 16718 4338
rect 16770 4286 16772 4338
rect 16604 4284 16772 4286
rect 16716 4274 16772 4284
rect 17388 4338 17444 4732
rect 17948 4562 18004 4956
rect 17948 4510 17950 4562
rect 18002 4510 18004 4562
rect 17948 4498 18004 4510
rect 18396 4452 18452 5854
rect 18844 5012 18900 6076
rect 20188 6020 20244 6030
rect 20188 5906 20244 5964
rect 20188 5854 20190 5906
rect 20242 5854 20244 5906
rect 20188 5842 20244 5854
rect 20748 5906 20804 7980
rect 21532 8036 21588 8046
rect 21532 7942 21588 7980
rect 21644 7924 21700 8204
rect 21756 8258 21812 9436
rect 21756 8206 21758 8258
rect 21810 8206 21812 8258
rect 21756 8194 21812 8206
rect 22428 8258 22484 9996
rect 22652 9828 22708 11340
rect 22764 11302 22820 11340
rect 22876 11172 22932 12014
rect 23996 11396 24052 16604
rect 24332 15988 24388 15998
rect 24220 15652 24276 15662
rect 24220 15314 24276 15596
rect 24332 15426 24388 15932
rect 24332 15374 24334 15426
rect 24386 15374 24388 15426
rect 24332 15362 24388 15374
rect 24444 15874 24500 15886
rect 24444 15822 24446 15874
rect 24498 15822 24500 15874
rect 24220 15262 24222 15314
rect 24274 15262 24276 15314
rect 24220 15250 24276 15262
rect 24444 15204 24500 15822
rect 24444 14756 24500 15148
rect 24444 14690 24500 14700
rect 24556 14532 24612 17500
rect 25340 17106 25396 18396
rect 25452 18386 25508 18396
rect 25900 18340 25956 20078
rect 26796 20130 26852 20188
rect 26796 20078 26798 20130
rect 26850 20078 26852 20130
rect 26796 20066 26852 20078
rect 26908 20412 27076 20468
rect 27132 20802 27188 20814
rect 27132 20750 27134 20802
rect 27186 20750 27188 20802
rect 26124 20018 26180 20030
rect 26124 19966 26126 20018
rect 26178 19966 26180 20018
rect 26124 18900 26180 19966
rect 26124 18834 26180 18844
rect 26460 18450 26516 18462
rect 26908 18452 26964 20412
rect 26460 18398 26462 18450
rect 26514 18398 26516 18450
rect 26348 18340 26404 18350
rect 25900 18274 25956 18284
rect 26236 18338 26404 18340
rect 26236 18286 26350 18338
rect 26402 18286 26404 18338
rect 26236 18284 26404 18286
rect 26124 18226 26180 18238
rect 26124 18174 26126 18226
rect 26178 18174 26180 18226
rect 26124 17668 26180 18174
rect 25340 17054 25342 17106
rect 25394 17054 25396 17106
rect 25340 17042 25396 17054
rect 25900 17612 26124 17668
rect 25676 16996 25732 17006
rect 24780 16884 24836 16894
rect 24780 16790 24836 16828
rect 25676 16882 25732 16940
rect 25676 16830 25678 16882
rect 25730 16830 25732 16882
rect 25676 16818 25732 16830
rect 25340 16100 25396 16110
rect 25788 16100 25844 16110
rect 25340 16006 25396 16044
rect 25564 16044 25788 16100
rect 24892 15988 24948 15998
rect 24892 15894 24948 15932
rect 25228 15428 25284 15438
rect 25228 15334 25284 15372
rect 25452 15428 25508 15438
rect 25452 15148 25508 15372
rect 24556 14466 24612 14476
rect 25228 15092 25508 15148
rect 24780 13636 24836 13646
rect 24780 13542 24836 13580
rect 25228 13636 25284 15092
rect 25452 14644 25508 14654
rect 25452 14550 25508 14588
rect 25340 14308 25396 14318
rect 25340 13970 25396 14252
rect 25340 13918 25342 13970
rect 25394 13918 25396 13970
rect 25340 13906 25396 13918
rect 25564 13748 25620 16044
rect 25788 16006 25844 16044
rect 25676 15426 25732 15438
rect 25676 15374 25678 15426
rect 25730 15374 25732 15426
rect 25676 15092 25732 15374
rect 25676 15026 25732 15036
rect 25788 15092 25844 15102
rect 25900 15092 25956 17612
rect 26124 17602 26180 17612
rect 26124 17220 26180 17230
rect 26124 16996 26180 17164
rect 26124 15314 26180 16940
rect 26124 15262 26126 15314
rect 26178 15262 26180 15314
rect 26124 15250 26180 15262
rect 26236 15316 26292 18284
rect 26348 18274 26404 18284
rect 26460 17780 26516 18398
rect 26460 17714 26516 17724
rect 26572 18450 26964 18452
rect 26572 18398 26910 18450
rect 26962 18398 26964 18450
rect 26572 18396 26964 18398
rect 26460 16996 26516 17006
rect 26572 16996 26628 18396
rect 26908 18358 26964 18396
rect 27020 20018 27076 20030
rect 27020 19966 27022 20018
rect 27074 19966 27076 20018
rect 27020 19012 27076 19966
rect 27132 19460 27188 20750
rect 27580 20468 27636 26124
rect 27692 21588 27748 27692
rect 27804 27300 27860 28476
rect 27804 27206 27860 27244
rect 27916 25620 27972 29372
rect 28028 29540 28084 29934
rect 28028 28868 28084 29484
rect 28140 28980 28196 30046
rect 29596 30098 29652 30156
rect 29596 30046 29598 30098
rect 29650 30046 29652 30098
rect 29036 29764 29092 29774
rect 28588 29652 28644 29662
rect 28588 29204 28644 29596
rect 28700 29540 28756 29550
rect 28700 29446 28756 29484
rect 28812 29426 28868 29438
rect 28812 29374 28814 29426
rect 28866 29374 28868 29426
rect 28700 29204 28756 29214
rect 28588 29202 28756 29204
rect 28588 29150 28702 29202
rect 28754 29150 28756 29202
rect 28588 29148 28756 29150
rect 28700 29138 28756 29148
rect 28812 28980 28868 29374
rect 28140 28924 28868 28980
rect 28028 28812 28308 28868
rect 28028 28418 28084 28430
rect 28028 28366 28030 28418
rect 28082 28366 28084 28418
rect 28028 28082 28084 28366
rect 28028 28030 28030 28082
rect 28082 28030 28084 28082
rect 28028 28018 28084 28030
rect 28252 28084 28308 28812
rect 28252 27990 28308 28028
rect 28364 27972 28420 27982
rect 28476 27972 28532 28924
rect 28812 28756 28868 28766
rect 28700 28644 28756 28654
rect 28700 28550 28756 28588
rect 28420 27916 28532 27972
rect 28364 27878 28420 27916
rect 28028 25620 28084 25630
rect 27916 25618 28084 25620
rect 27916 25566 28030 25618
rect 28082 25566 28084 25618
rect 27916 25564 28084 25566
rect 27804 24836 27860 24846
rect 27804 23604 27860 24780
rect 27804 23538 27860 23548
rect 27916 22708 27972 25564
rect 28028 25554 28084 25564
rect 28588 25284 28644 25294
rect 28588 25190 28644 25228
rect 28140 23716 28196 23726
rect 28140 23622 28196 23660
rect 28812 23268 28868 28700
rect 29036 24836 29092 29708
rect 29260 29428 29316 29438
rect 29260 29334 29316 29372
rect 29596 28756 29652 30046
rect 29708 30100 29764 30110
rect 29764 30044 29876 30100
rect 29708 30034 29764 30044
rect 29708 29764 29764 29774
rect 29708 29426 29764 29708
rect 29820 29652 29876 30044
rect 29932 30098 29988 30940
rect 30268 30212 30324 31054
rect 30492 30322 30548 37212
rect 31052 36372 31108 36382
rect 31052 35026 31108 36316
rect 31836 36260 31892 37772
rect 31052 34974 31054 35026
rect 31106 34974 31108 35026
rect 31052 34962 31108 34974
rect 31500 36204 31892 36260
rect 31948 36482 32004 36494
rect 31948 36430 31950 36482
rect 32002 36430 32004 36482
rect 31164 34804 31220 34814
rect 31164 34710 31220 34748
rect 30940 34690 30996 34702
rect 30940 34638 30942 34690
rect 30994 34638 30996 34690
rect 30940 34354 30996 34638
rect 30940 34302 30942 34354
rect 30994 34302 30996 34354
rect 30940 34290 30996 34302
rect 31052 34244 31108 34254
rect 31052 34150 31108 34188
rect 30604 34130 30660 34142
rect 30604 34078 30606 34130
rect 30658 34078 30660 34130
rect 30604 33684 30660 34078
rect 30604 33618 30660 33628
rect 31276 34130 31332 34142
rect 31276 34078 31278 34130
rect 31330 34078 31332 34130
rect 31276 31948 31332 34078
rect 31500 31948 31556 36204
rect 31836 35812 31892 35822
rect 31948 35812 32004 36430
rect 32732 36372 32788 36382
rect 32732 36278 32788 36316
rect 31836 35810 32004 35812
rect 31836 35758 31838 35810
rect 31890 35758 32004 35810
rect 31836 35756 32004 35758
rect 31836 35364 31892 35756
rect 32172 35700 32228 35710
rect 32172 35698 32452 35700
rect 32172 35646 32174 35698
rect 32226 35646 32452 35698
rect 32172 35644 32452 35646
rect 32172 35634 32228 35644
rect 31612 34916 31668 34926
rect 31836 34916 31892 35308
rect 32284 35028 32340 35038
rect 32284 34934 32340 34972
rect 31612 34914 31892 34916
rect 31612 34862 31614 34914
rect 31666 34862 31892 34914
rect 31612 34860 31892 34862
rect 31612 33346 31668 34860
rect 32396 34356 32452 35644
rect 32284 34244 32340 34254
rect 32284 34150 32340 34188
rect 31948 34132 32004 34142
rect 31948 34038 32004 34076
rect 32060 34020 32116 34030
rect 32060 33926 32116 33964
rect 32396 33572 32452 34300
rect 32508 35588 32564 35598
rect 32508 34242 32564 35532
rect 32508 34190 32510 34242
rect 32562 34190 32564 34242
rect 32508 34178 32564 34190
rect 31612 33294 31614 33346
rect 31666 33294 31668 33346
rect 31612 33282 31668 33294
rect 32284 33516 32452 33572
rect 32508 33684 32564 33694
rect 32172 32562 32228 32574
rect 32172 32510 32174 32562
rect 32226 32510 32228 32562
rect 31836 32004 31892 32042
rect 32172 31948 32228 32510
rect 31052 31892 31108 31902
rect 31276 31892 31444 31948
rect 31500 31892 31668 31948
rect 31836 31938 31892 31948
rect 30940 31108 30996 31118
rect 31052 31108 31108 31836
rect 30940 31106 31108 31108
rect 30940 31054 30942 31106
rect 30994 31054 31108 31106
rect 30940 31052 31108 31054
rect 31276 31778 31332 31790
rect 31276 31726 31278 31778
rect 31330 31726 31332 31778
rect 30940 31042 30996 31052
rect 30604 30996 30660 31006
rect 30604 30994 30884 30996
rect 30604 30942 30606 30994
rect 30658 30942 30884 30994
rect 30604 30940 30884 30942
rect 30604 30930 30660 30940
rect 30492 30270 30494 30322
rect 30546 30270 30548 30322
rect 30492 30258 30548 30270
rect 30716 30324 30772 30334
rect 30268 30146 30324 30156
rect 30604 30210 30660 30222
rect 30604 30158 30606 30210
rect 30658 30158 30660 30210
rect 29932 30046 29934 30098
rect 29986 30046 29988 30098
rect 29932 30034 29988 30046
rect 30604 30100 30660 30158
rect 30604 30034 30660 30044
rect 29932 29652 29988 29662
rect 29820 29650 29988 29652
rect 29820 29598 29934 29650
rect 29986 29598 29988 29650
rect 29820 29596 29988 29598
rect 29932 29586 29988 29596
rect 30604 29652 30660 29662
rect 30716 29652 30772 30268
rect 30828 29876 30884 30940
rect 31276 30994 31332 31726
rect 31276 30942 31278 30994
rect 31330 30942 31332 30994
rect 31276 30436 31332 30942
rect 31388 30772 31444 31892
rect 31612 31444 31668 31892
rect 31948 31892 32228 31948
rect 31948 31780 32004 31892
rect 31612 30884 31668 31388
rect 31836 31724 32004 31780
rect 31724 31220 31780 31230
rect 31836 31220 31892 31724
rect 31724 31218 31892 31220
rect 31724 31166 31726 31218
rect 31778 31166 31892 31218
rect 31724 31164 31892 31166
rect 31724 31154 31780 31164
rect 31612 30818 31668 30828
rect 31724 30994 31780 31006
rect 31724 30942 31726 30994
rect 31778 30942 31780 30994
rect 31500 30772 31556 30782
rect 31388 30716 31500 30772
rect 31500 30678 31556 30716
rect 31276 30370 31332 30380
rect 31276 30098 31332 30110
rect 31276 30046 31278 30098
rect 31330 30046 31332 30098
rect 30828 29820 30996 29876
rect 30604 29650 30772 29652
rect 30604 29598 30606 29650
rect 30658 29598 30772 29650
rect 30604 29596 30772 29598
rect 30604 29586 30660 29596
rect 29708 29374 29710 29426
rect 29762 29374 29764 29426
rect 29708 29362 29764 29374
rect 30156 29428 30212 29438
rect 29596 28690 29652 28700
rect 29820 29092 29876 29102
rect 29708 28644 29764 28654
rect 29708 28550 29764 28588
rect 29820 28532 29876 29036
rect 30156 28532 30212 29372
rect 30268 29426 30324 29438
rect 30268 29374 30270 29426
rect 30322 29374 30324 29426
rect 30268 28868 30324 29374
rect 30268 28802 30324 28812
rect 30492 29426 30548 29438
rect 30492 29374 30494 29426
rect 30546 29374 30548 29426
rect 29820 28438 29876 28476
rect 30044 28530 30212 28532
rect 30044 28478 30158 28530
rect 30210 28478 30212 28530
rect 30044 28476 30212 28478
rect 29148 27972 29204 27982
rect 29148 27878 29204 27916
rect 29596 27860 29652 27870
rect 29596 27766 29652 27804
rect 29260 27748 29316 27758
rect 29260 27654 29316 27692
rect 30044 27524 30100 28476
rect 30156 28466 30212 28476
rect 30268 28644 30324 28654
rect 30492 28644 30548 29374
rect 30716 29426 30772 29438
rect 30716 29374 30718 29426
rect 30770 29374 30772 29426
rect 30716 29092 30772 29374
rect 30828 29428 30884 29438
rect 30828 29334 30884 29372
rect 30716 29026 30772 29036
rect 30716 28868 30772 28878
rect 30716 28774 30772 28812
rect 30940 28754 30996 29820
rect 31276 29540 31332 30046
rect 31276 29474 31332 29484
rect 31724 29988 31780 30942
rect 31948 30322 32004 30334
rect 31948 30270 31950 30322
rect 32002 30270 32004 30322
rect 31948 30100 32004 30270
rect 32284 30210 32340 33516
rect 32396 33234 32452 33246
rect 32396 33182 32398 33234
rect 32450 33182 32452 33234
rect 32396 32786 32452 33182
rect 32396 32734 32398 32786
rect 32450 32734 32452 32786
rect 32396 32722 32452 32734
rect 32508 32674 32564 33628
rect 32508 32622 32510 32674
rect 32562 32622 32564 32674
rect 32508 32610 32564 32622
rect 32844 31948 32900 41804
rect 33852 41300 33908 41918
rect 33852 41234 33908 41244
rect 34188 41970 34244 41982
rect 34188 41918 34190 41970
rect 34242 41918 34244 41970
rect 34188 40964 34244 41918
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 34636 41298 34692 41310
rect 34636 41246 34638 41298
rect 34690 41246 34692 41298
rect 34636 41188 34692 41246
rect 35532 41188 35588 41198
rect 34636 41132 35140 41188
rect 34860 40964 34916 40974
rect 34188 40962 34916 40964
rect 34188 40910 34862 40962
rect 34914 40910 34916 40962
rect 34188 40908 34916 40910
rect 33964 40514 34020 40526
rect 33964 40462 33966 40514
rect 34018 40462 34020 40514
rect 33068 40404 33124 40414
rect 33068 40310 33124 40348
rect 33516 40404 33572 40414
rect 33516 40310 33572 40348
rect 33740 40402 33796 40414
rect 33740 40350 33742 40402
rect 33794 40350 33796 40402
rect 33740 40292 33796 40350
rect 33740 40226 33796 40236
rect 33964 40180 34020 40462
rect 33964 40114 34020 40124
rect 34076 40290 34132 40302
rect 34076 40238 34078 40290
rect 34130 40238 34132 40290
rect 34076 39844 34132 40238
rect 34412 40292 34468 40302
rect 34412 40198 34468 40236
rect 34076 39778 34132 39788
rect 34524 40180 34580 40190
rect 33180 39506 33236 39518
rect 33180 39454 33182 39506
rect 33234 39454 33236 39506
rect 33068 38836 33124 38846
rect 33068 38742 33124 38780
rect 33180 38162 33236 39454
rect 33852 38722 33908 38734
rect 33852 38670 33854 38722
rect 33906 38670 33908 38722
rect 33852 38668 33908 38670
rect 34524 38724 34580 40124
rect 34860 39620 34916 40908
rect 34860 39554 34916 39564
rect 34972 40962 35028 40974
rect 34972 40910 34974 40962
rect 35026 40910 35028 40962
rect 34972 38668 35028 40910
rect 35084 40404 35140 41132
rect 35532 41186 35700 41188
rect 35532 41134 35534 41186
rect 35586 41134 35700 41186
rect 35532 41132 35700 41134
rect 35532 41122 35588 41132
rect 35084 40338 35140 40348
rect 35196 40962 35252 40974
rect 35196 40910 35198 40962
rect 35250 40910 35252 40962
rect 35196 40180 35252 40910
rect 35196 40114 35252 40124
rect 35644 40292 35700 41132
rect 38108 41186 38164 41198
rect 38108 41134 38110 41186
rect 38162 41134 38164 41186
rect 36092 41076 36148 41086
rect 36092 41074 36932 41076
rect 36092 41022 36094 41074
rect 36146 41022 36932 41074
rect 36092 41020 36932 41022
rect 36092 41010 36148 41020
rect 35868 40964 35924 40974
rect 35868 40870 35924 40908
rect 35980 40962 36036 40974
rect 35980 40910 35982 40962
rect 36034 40910 36036 40962
rect 35980 40628 36036 40910
rect 35980 40572 36596 40628
rect 36540 40514 36596 40572
rect 36540 40462 36542 40514
rect 36594 40462 36596 40514
rect 36540 40450 36596 40462
rect 36428 40404 36484 40414
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35308 39844 35364 39854
rect 35308 39730 35364 39788
rect 35308 39678 35310 39730
rect 35362 39678 35364 39730
rect 35308 38668 35364 39678
rect 35644 39618 35700 40236
rect 35980 40292 36036 40302
rect 36036 40236 36148 40292
rect 35980 40226 36036 40236
rect 36092 39730 36148 40236
rect 36092 39678 36094 39730
rect 36146 39678 36148 39730
rect 36092 39666 36148 39678
rect 35644 39566 35646 39618
rect 35698 39566 35700 39618
rect 35644 39554 35700 39566
rect 33180 38110 33182 38162
rect 33234 38110 33236 38162
rect 33180 38098 33236 38110
rect 33740 38612 33908 38668
rect 34412 38612 34580 38668
rect 34748 38612 35028 38668
rect 35084 38612 35364 38668
rect 35868 39506 35924 39518
rect 35868 39454 35870 39506
rect 35922 39454 35924 39506
rect 33292 38052 33348 38062
rect 33292 37958 33348 37996
rect 33628 37938 33684 37950
rect 33628 37886 33630 37938
rect 33682 37886 33684 37938
rect 33068 37826 33124 37838
rect 33068 37774 33070 37826
rect 33122 37774 33124 37826
rect 33068 37268 33124 37774
rect 33628 37378 33684 37886
rect 33740 37490 33796 38612
rect 34412 38162 34468 38612
rect 34412 38110 34414 38162
rect 34466 38110 34468 38162
rect 34412 38098 34468 38110
rect 34076 38052 34132 38062
rect 34076 37958 34132 37996
rect 34748 38052 34804 38612
rect 34748 37986 34804 37996
rect 35084 38050 35140 38612
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35084 37998 35086 38050
rect 35138 37998 35140 38050
rect 35084 37986 35140 37998
rect 35420 38052 35476 38062
rect 35868 38052 35924 39454
rect 36204 39506 36260 39518
rect 36204 39454 36206 39506
rect 36258 39454 36260 39506
rect 35980 38724 36036 38762
rect 36204 38724 36260 39454
rect 36316 39060 36372 39070
rect 36316 38966 36372 39004
rect 36428 38946 36484 40348
rect 36876 39844 36932 41020
rect 37548 40740 37604 40750
rect 37324 40402 37380 40414
rect 37324 40350 37326 40402
rect 37378 40350 37380 40402
rect 37100 39844 37156 39854
rect 36876 39842 37156 39844
rect 36876 39790 37102 39842
rect 37154 39790 37156 39842
rect 36876 39788 37156 39790
rect 37100 39778 37156 39788
rect 36988 39620 37044 39630
rect 36988 39526 37044 39564
rect 36428 38894 36430 38946
rect 36482 38894 36484 38946
rect 36428 38882 36484 38894
rect 37100 39394 37156 39406
rect 37100 39342 37102 39394
rect 37154 39342 37156 39394
rect 36036 38668 36260 38724
rect 35980 38658 36036 38668
rect 37100 38500 37156 39342
rect 37324 38724 37380 40350
rect 37548 39618 37604 40684
rect 38108 40740 38164 41134
rect 38780 41076 38836 41086
rect 38108 40674 38164 40684
rect 38220 41074 38836 41076
rect 38220 41022 38782 41074
rect 38834 41022 38836 41074
rect 38220 41020 38836 41022
rect 38220 40626 38276 41020
rect 38780 41010 38836 41020
rect 39340 41076 39396 41086
rect 38220 40574 38222 40626
rect 38274 40574 38276 40626
rect 38220 40562 38276 40574
rect 39116 40628 39172 40638
rect 39116 40534 39172 40572
rect 39340 40626 39396 41020
rect 39340 40574 39342 40626
rect 39394 40574 39396 40626
rect 39340 40562 39396 40574
rect 39564 40684 40180 40740
rect 37548 39566 37550 39618
rect 37602 39566 37604 39618
rect 37324 38658 37380 38668
rect 37436 38836 37492 38846
rect 37436 38500 37492 38780
rect 37548 38612 37604 39566
rect 37884 40516 37940 40526
rect 37884 38834 37940 40460
rect 39564 40514 39620 40684
rect 39564 40462 39566 40514
rect 39618 40462 39620 40514
rect 39564 40450 39620 40462
rect 39676 40516 39732 40526
rect 39676 40514 39844 40516
rect 39676 40462 39678 40514
rect 39730 40462 39844 40514
rect 39676 40460 39844 40462
rect 39676 40450 39732 40460
rect 39004 40402 39060 40414
rect 39004 40350 39006 40402
rect 39058 40350 39060 40402
rect 38108 40290 38164 40302
rect 38108 40238 38110 40290
rect 38162 40238 38164 40290
rect 38108 39172 38164 40238
rect 38668 40292 38724 40302
rect 38668 40290 38948 40292
rect 38668 40238 38670 40290
rect 38722 40238 38948 40290
rect 38668 40236 38948 40238
rect 38668 40226 38724 40236
rect 38556 40180 38612 40190
rect 38332 40178 38612 40180
rect 38332 40126 38558 40178
rect 38610 40126 38612 40178
rect 38332 40124 38612 40126
rect 38332 39730 38388 40124
rect 38556 40114 38612 40124
rect 38332 39678 38334 39730
rect 38386 39678 38388 39730
rect 38332 39666 38388 39678
rect 38892 39508 38948 40236
rect 39004 39732 39060 40350
rect 39788 40292 39844 40460
rect 39788 40226 39844 40236
rect 39900 40402 39956 40414
rect 39900 40350 39902 40402
rect 39954 40350 39956 40402
rect 39004 39666 39060 39676
rect 38892 39452 39620 39508
rect 38108 39116 38612 39172
rect 38556 39060 38612 39116
rect 38668 39060 38724 39070
rect 38892 39060 38948 39070
rect 38556 39058 38724 39060
rect 38556 39006 38670 39058
rect 38722 39006 38724 39058
rect 38556 39004 38724 39006
rect 38668 38994 38724 39004
rect 38780 39004 38892 39060
rect 37884 38782 37886 38834
rect 37938 38782 37940 38834
rect 37884 38770 37940 38782
rect 38220 38946 38276 38958
rect 38220 38894 38222 38946
rect 38274 38894 38276 38946
rect 37996 38612 38052 38622
rect 37548 38546 37604 38556
rect 37660 38610 38052 38612
rect 37660 38558 37998 38610
rect 38050 38558 38052 38610
rect 37660 38556 38052 38558
rect 37100 38444 37492 38500
rect 35476 37996 35924 38052
rect 36988 38164 37044 38174
rect 35420 37938 35476 37996
rect 35420 37886 35422 37938
rect 35474 37886 35476 37938
rect 35420 37874 35476 37886
rect 36988 37938 37044 38108
rect 37212 38052 37268 38062
rect 36988 37886 36990 37938
rect 37042 37886 37044 37938
rect 36988 37874 37044 37886
rect 37100 38050 37268 38052
rect 37100 37998 37214 38050
rect 37266 37998 37268 38050
rect 37100 37996 37268 37998
rect 37100 37604 37156 37996
rect 37212 37986 37268 37996
rect 33740 37438 33742 37490
rect 33794 37438 33796 37490
rect 33740 37426 33796 37438
rect 36764 37548 37156 37604
rect 33628 37326 33630 37378
rect 33682 37326 33684 37378
rect 33628 37314 33684 37326
rect 33068 37202 33124 37212
rect 33964 37268 34020 37278
rect 33964 37174 34020 37212
rect 35084 37268 35140 37278
rect 34860 36594 34916 36606
rect 34860 36542 34862 36594
rect 34914 36542 34916 36594
rect 32956 35812 33012 35822
rect 32956 35698 33012 35756
rect 34860 35812 34916 36542
rect 34860 35746 34916 35756
rect 32956 35646 32958 35698
rect 33010 35646 33012 35698
rect 32956 35634 33012 35646
rect 33404 35700 33460 35710
rect 33404 35698 33572 35700
rect 33404 35646 33406 35698
rect 33458 35646 33572 35698
rect 33404 35644 33572 35646
rect 33404 35634 33460 35644
rect 33180 35586 33236 35598
rect 33180 35534 33182 35586
rect 33234 35534 33236 35586
rect 33180 35028 33236 35534
rect 33180 34962 33236 34972
rect 33292 35364 33348 35374
rect 33068 34132 33124 34142
rect 33292 34132 33348 35308
rect 33068 34130 33348 34132
rect 33068 34078 33070 34130
rect 33122 34078 33348 34130
rect 33068 34076 33348 34078
rect 33516 34244 33572 35644
rect 33628 35698 33684 35710
rect 33628 35646 33630 35698
rect 33682 35646 33684 35698
rect 33628 35028 33684 35646
rect 33628 34962 33684 34972
rect 34412 35026 34468 35038
rect 34412 34974 34414 35026
rect 34466 34974 34468 35026
rect 34412 34692 34468 34974
rect 34412 34626 34468 34636
rect 33068 34066 33124 34076
rect 32732 31892 32900 31948
rect 33180 32562 33236 32574
rect 33180 32510 33182 32562
rect 33234 32510 33236 32562
rect 33180 32004 33236 32510
rect 33516 32562 33572 34188
rect 33852 34020 33908 34030
rect 33852 33926 33908 33964
rect 34524 33908 34580 33918
rect 34524 33458 34580 33852
rect 34524 33406 34526 33458
rect 34578 33406 34580 33458
rect 34524 33394 34580 33406
rect 33852 33124 33908 33134
rect 33852 32674 33908 33068
rect 33852 32622 33854 32674
rect 33906 32622 33908 32674
rect 33852 32610 33908 32622
rect 33516 32510 33518 32562
rect 33570 32510 33572 32562
rect 33516 32498 33572 32510
rect 33180 31938 33236 31948
rect 33404 32450 33460 32462
rect 33404 32398 33406 32450
rect 33458 32398 33460 32450
rect 33404 31948 33460 32398
rect 34972 32452 35028 32462
rect 34972 32358 35028 32396
rect 34636 32338 34692 32350
rect 34636 32286 34638 32338
rect 34690 32286 34692 32338
rect 34636 31948 34692 32286
rect 35084 31948 35140 37212
rect 35868 37268 35924 37278
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35532 35812 35588 35822
rect 35532 35718 35588 35756
rect 35756 35700 35812 35710
rect 35644 35698 35812 35700
rect 35644 35646 35758 35698
rect 35810 35646 35812 35698
rect 35644 35644 35812 35646
rect 35420 35588 35476 35598
rect 35420 35494 35476 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35420 35028 35476 35038
rect 35308 34916 35364 34926
rect 35308 34822 35364 34860
rect 35420 34914 35476 34972
rect 35644 35028 35700 35644
rect 35756 35634 35812 35644
rect 35420 34862 35422 34914
rect 35474 34862 35476 34914
rect 35420 34850 35476 34862
rect 35532 34916 35588 34926
rect 35644 34916 35700 34972
rect 35532 34914 35700 34916
rect 35532 34862 35534 34914
rect 35586 34862 35700 34914
rect 35532 34860 35700 34862
rect 35532 34850 35588 34860
rect 35868 34802 35924 37212
rect 36764 37268 36820 37548
rect 36764 37174 36820 37212
rect 36988 37378 37044 37390
rect 36988 37326 36990 37378
rect 37042 37326 37044 37378
rect 36988 37044 37044 37326
rect 37212 37044 37268 37054
rect 37324 37044 37380 38444
rect 37660 37492 37716 38556
rect 37996 38546 38052 38556
rect 38108 38612 38164 38622
rect 36988 37042 37380 37044
rect 36988 36990 37214 37042
rect 37266 36990 37380 37042
rect 36988 36988 37380 36990
rect 37436 37436 37716 37492
rect 37212 36978 37268 36988
rect 35980 35924 36036 35934
rect 35980 35830 36036 35868
rect 37212 35924 37268 35934
rect 36764 35812 36820 35822
rect 36764 35718 36820 35756
rect 36316 35700 36372 35710
rect 36316 35606 36372 35644
rect 36428 35474 36484 35486
rect 36428 35422 36430 35474
rect 36482 35422 36484 35474
rect 35868 34750 35870 34802
rect 35922 34750 35924 34802
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35420 33572 35476 33582
rect 35420 33478 35476 33516
rect 35756 33572 35812 33582
rect 35532 33348 35588 33358
rect 35532 33254 35588 33292
rect 35644 33236 35700 33246
rect 35196 32564 35252 32574
rect 35196 32470 35252 32508
rect 35644 32562 35700 33180
rect 35644 32510 35646 32562
rect 35698 32510 35700 32562
rect 35644 32498 35700 32510
rect 35532 32338 35588 32350
rect 35532 32286 35534 32338
rect 35586 32286 35588 32338
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35532 31948 35588 32286
rect 33404 31892 33572 31948
rect 34636 31892 34916 31948
rect 35084 31892 35252 31948
rect 32732 31778 32788 31892
rect 33516 31890 33572 31892
rect 33516 31838 33518 31890
rect 33570 31838 33572 31890
rect 33516 31826 33572 31838
rect 32732 31726 32734 31778
rect 32786 31726 32788 31778
rect 32284 30158 32286 30210
rect 32338 30158 32340 30210
rect 32284 30146 32340 30158
rect 32396 31556 32452 31566
rect 32732 31556 32788 31726
rect 32396 31554 32788 31556
rect 32396 31502 32398 31554
rect 32450 31502 32788 31554
rect 32396 31500 32788 31502
rect 31724 28868 31780 29932
rect 31836 30044 32228 30100
rect 31836 29204 31892 30044
rect 32172 29988 32228 30044
rect 32396 29988 32452 31500
rect 33068 31108 33124 31118
rect 34860 31108 34916 31892
rect 35084 31108 35140 31118
rect 34860 31106 35140 31108
rect 34860 31054 35086 31106
rect 35138 31054 35140 31106
rect 34860 31052 35140 31054
rect 32508 30996 32564 31006
rect 32620 30996 32676 31006
rect 32508 30994 32620 30996
rect 32508 30942 32510 30994
rect 32562 30942 32620 30994
rect 32508 30940 32620 30942
rect 32508 30930 32564 30940
rect 32172 29932 32452 29988
rect 31948 29876 32004 29886
rect 31948 29426 32004 29820
rect 32508 29652 32564 29662
rect 32508 29538 32564 29596
rect 32508 29486 32510 29538
rect 32562 29486 32564 29538
rect 32508 29474 32564 29486
rect 31948 29374 31950 29426
rect 32002 29374 32004 29426
rect 31948 29362 32004 29374
rect 32396 29204 32452 29214
rect 31836 29148 32004 29204
rect 31724 28802 31780 28812
rect 30940 28702 30942 28754
rect 30994 28702 30996 28754
rect 30940 28690 30996 28702
rect 30268 28642 30548 28644
rect 30268 28590 30270 28642
rect 30322 28590 30548 28642
rect 30268 28588 30548 28590
rect 31948 28644 32004 29148
rect 32396 29110 32452 29148
rect 30268 28420 30324 28588
rect 30268 27972 30324 28364
rect 30268 27906 30324 27916
rect 30380 27748 30436 27758
rect 30380 27654 30436 27692
rect 29596 27468 30100 27524
rect 29596 27186 29652 27468
rect 29596 27134 29598 27186
rect 29650 27134 29652 27186
rect 29596 27122 29652 27134
rect 30044 26404 30100 27468
rect 31724 26964 31780 26974
rect 30940 26962 31780 26964
rect 30940 26910 31726 26962
rect 31778 26910 31780 26962
rect 30940 26908 31780 26910
rect 30940 26514 30996 26908
rect 31724 26898 31780 26908
rect 30940 26462 30942 26514
rect 30994 26462 30996 26514
rect 30940 26450 30996 26462
rect 30044 26338 30100 26348
rect 30828 26404 30884 26414
rect 30828 26310 30884 26348
rect 31836 26068 31892 26078
rect 31724 26012 31836 26068
rect 29260 25284 29316 25294
rect 29260 25190 29316 25228
rect 31724 25284 31780 26012
rect 31836 26002 31892 26012
rect 31948 25508 32004 28588
rect 32508 28420 32564 28430
rect 32508 27746 32564 28364
rect 32508 27694 32510 27746
rect 32562 27694 32564 27746
rect 32508 27682 32564 27694
rect 31948 25442 32004 25452
rect 32396 27074 32452 27086
rect 32396 27022 32398 27074
rect 32450 27022 32452 27074
rect 29036 24780 30100 24836
rect 29036 24722 29092 24780
rect 29036 24670 29038 24722
rect 29090 24670 29092 24722
rect 29036 24658 29092 24670
rect 29708 24612 29764 24622
rect 29260 24610 29764 24612
rect 29260 24558 29710 24610
rect 29762 24558 29764 24610
rect 29260 24556 29764 24558
rect 29260 24050 29316 24556
rect 29708 24546 29764 24556
rect 29260 23998 29262 24050
rect 29314 23998 29316 24050
rect 29260 23986 29316 23998
rect 29484 23940 29540 23950
rect 29484 23846 29540 23884
rect 29596 23938 29652 23950
rect 29596 23886 29598 23938
rect 29650 23886 29652 23938
rect 29148 23826 29204 23838
rect 29148 23774 29150 23826
rect 29202 23774 29204 23826
rect 28812 23202 28868 23212
rect 28924 23716 28980 23726
rect 28476 23156 28532 23166
rect 28476 23062 28532 23100
rect 28700 23154 28756 23166
rect 28700 23102 28702 23154
rect 28754 23102 28756 23154
rect 27804 22652 27972 22708
rect 28140 23042 28196 23054
rect 28140 22990 28142 23042
rect 28194 22990 28196 23042
rect 28140 22708 28196 22990
rect 27804 22260 27860 22652
rect 28140 22642 28196 22652
rect 27804 22194 27860 22204
rect 27916 22484 27972 22494
rect 27972 22428 28308 22484
rect 27692 21522 27748 21532
rect 27804 21924 27860 21934
rect 27804 20804 27860 21868
rect 27916 20914 27972 22428
rect 28252 22370 28308 22428
rect 28252 22318 28254 22370
rect 28306 22318 28308 22370
rect 28252 22306 28308 22318
rect 28588 22260 28644 22270
rect 28588 22166 28644 22204
rect 28700 21924 28756 23102
rect 28924 23154 28980 23660
rect 28924 23102 28926 23154
rect 28978 23102 28980 23154
rect 28812 23044 28868 23054
rect 28812 22950 28868 22988
rect 28700 21858 28756 21868
rect 28140 21812 28196 21822
rect 28140 21474 28196 21756
rect 28588 21700 28644 21710
rect 28588 21606 28644 21644
rect 28140 21422 28142 21474
rect 28194 21422 28196 21474
rect 28140 21410 28196 21422
rect 28476 21586 28532 21598
rect 28476 21534 28478 21586
rect 28530 21534 28532 21586
rect 28476 20916 28532 21534
rect 28924 21476 28980 23102
rect 29036 23154 29092 23166
rect 29036 23102 29038 23154
rect 29090 23102 29092 23154
rect 29036 23044 29092 23102
rect 29036 22978 29092 22988
rect 29148 22260 29204 23774
rect 29260 23604 29316 23614
rect 29316 23548 29428 23604
rect 29260 23538 29316 23548
rect 29148 22194 29204 22204
rect 28812 21420 28980 21476
rect 29036 22036 29092 22046
rect 29036 21588 29092 21980
rect 29148 21588 29204 21598
rect 29036 21586 29204 21588
rect 29036 21534 29150 21586
rect 29202 21534 29204 21586
rect 29036 21532 29204 21534
rect 28588 21364 28644 21374
rect 28588 21270 28644 21308
rect 27916 20862 27918 20914
rect 27970 20862 27972 20914
rect 27916 20850 27972 20862
rect 28252 20860 28532 20916
rect 27580 20402 27636 20412
rect 27692 20802 27860 20804
rect 27692 20750 27806 20802
rect 27858 20750 27860 20802
rect 27692 20748 27860 20750
rect 27580 20018 27636 20030
rect 27580 19966 27582 20018
rect 27634 19966 27636 20018
rect 27580 19460 27636 19966
rect 27132 19458 27636 19460
rect 27132 19406 27134 19458
rect 27186 19406 27636 19458
rect 27132 19404 27636 19406
rect 27132 19394 27188 19404
rect 27692 19348 27748 20748
rect 27804 20738 27860 20748
rect 28140 20692 28196 20702
rect 28252 20692 28308 20860
rect 28476 20692 28532 20702
rect 28140 20690 28308 20692
rect 28140 20638 28142 20690
rect 28194 20638 28308 20690
rect 28140 20636 28308 20638
rect 28364 20636 28476 20692
rect 27916 20132 27972 20142
rect 27916 20038 27972 20076
rect 27244 19292 27748 19348
rect 27244 19234 27300 19292
rect 27244 19182 27246 19234
rect 27298 19182 27300 19234
rect 27244 19170 27300 19182
rect 27132 19012 27188 19022
rect 27020 19010 27188 19012
rect 27020 18958 27134 19010
rect 27186 18958 27188 19010
rect 27020 18956 27188 18958
rect 27020 18228 27076 18956
rect 27132 18946 27188 18956
rect 27580 19012 27636 19022
rect 26460 16994 26628 16996
rect 26460 16942 26462 16994
rect 26514 16942 26628 16994
rect 26460 16940 26628 16942
rect 26684 18172 27076 18228
rect 26460 16930 26516 16940
rect 26348 16882 26404 16894
rect 26348 16830 26350 16882
rect 26402 16830 26404 16882
rect 26348 15652 26404 16830
rect 26684 16212 26740 18172
rect 27580 17892 27636 18956
rect 27580 17826 27636 17836
rect 27692 18452 27748 19292
rect 27916 19124 27972 19134
rect 27916 19030 27972 19068
rect 27692 17890 27748 18396
rect 27692 17838 27694 17890
rect 27746 17838 27748 17890
rect 27692 17826 27748 17838
rect 27804 18564 27860 18574
rect 26796 17780 26852 17790
rect 26796 17220 26852 17724
rect 27132 17668 27188 17678
rect 26796 17154 26852 17164
rect 27020 17666 27188 17668
rect 27020 17614 27134 17666
rect 27186 17614 27188 17666
rect 27020 17612 27188 17614
rect 26404 15596 26516 15652
rect 26348 15586 26404 15596
rect 26348 15428 26404 15438
rect 26348 15334 26404 15372
rect 26236 15250 26292 15260
rect 26460 15148 26516 15596
rect 25788 15090 25956 15092
rect 25788 15038 25790 15090
rect 25842 15038 25956 15090
rect 25788 15036 25956 15038
rect 26236 15092 26516 15148
rect 25788 15026 25844 15036
rect 26012 14756 26068 14766
rect 25788 14644 25844 14654
rect 25788 14530 25844 14588
rect 25788 14478 25790 14530
rect 25842 14478 25844 14530
rect 25564 13746 25732 13748
rect 25564 13694 25566 13746
rect 25618 13694 25732 13746
rect 25564 13692 25732 13694
rect 25564 13682 25620 13692
rect 25228 13570 25284 13580
rect 25676 12740 25732 13692
rect 25788 12962 25844 14478
rect 26012 14530 26068 14700
rect 26012 14478 26014 14530
rect 26066 14478 26068 14530
rect 26012 14466 26068 14478
rect 26124 14420 26180 14430
rect 26124 14326 26180 14364
rect 26236 13970 26292 15092
rect 26236 13918 26238 13970
rect 26290 13918 26292 13970
rect 26236 13906 26292 13918
rect 26460 14756 26516 14766
rect 26460 13746 26516 14700
rect 26572 14756 26628 14766
rect 26684 14756 26740 16156
rect 26572 14754 26740 14756
rect 26572 14702 26574 14754
rect 26626 14702 26740 14754
rect 26572 14700 26740 14702
rect 26796 16884 26852 16894
rect 26796 15426 26852 16828
rect 26908 16772 26964 16782
rect 26908 16322 26964 16716
rect 26908 16270 26910 16322
rect 26962 16270 26964 16322
rect 26908 16258 26964 16270
rect 27020 16324 27076 17612
rect 27132 17602 27188 17612
rect 27356 17668 27412 17678
rect 27356 16884 27412 17612
rect 27804 17106 27860 18508
rect 27916 18338 27972 18350
rect 27916 18286 27918 18338
rect 27970 18286 27972 18338
rect 27916 18228 27972 18286
rect 27916 18162 27972 18172
rect 28140 17778 28196 20636
rect 28252 20132 28308 20142
rect 28252 19458 28308 20076
rect 28252 19406 28254 19458
rect 28306 19406 28308 19458
rect 28252 19394 28308 19406
rect 28364 19346 28420 20636
rect 28476 20626 28532 20636
rect 28476 20468 28532 20478
rect 28476 19796 28532 20412
rect 28588 20020 28644 20030
rect 28588 20018 28756 20020
rect 28588 19966 28590 20018
rect 28642 19966 28756 20018
rect 28588 19964 28756 19966
rect 28588 19954 28644 19964
rect 28476 19740 28644 19796
rect 28364 19294 28366 19346
rect 28418 19294 28420 19346
rect 28364 19282 28420 19294
rect 28588 19124 28644 19740
rect 28700 19460 28756 19964
rect 28700 19394 28756 19404
rect 28588 19068 28756 19124
rect 28476 19010 28532 19022
rect 28476 18958 28478 19010
rect 28530 18958 28532 19010
rect 28364 18564 28420 18574
rect 28364 18470 28420 18508
rect 28252 18452 28308 18462
rect 28252 18358 28308 18396
rect 28476 18228 28532 18958
rect 28476 18162 28532 18172
rect 28140 17726 28142 17778
rect 28194 17726 28196 17778
rect 28140 17714 28196 17726
rect 28252 17780 28308 17790
rect 28308 17724 28420 17780
rect 28252 17714 28308 17724
rect 27804 17054 27806 17106
rect 27858 17054 27860 17106
rect 27804 17042 27860 17054
rect 28028 17554 28084 17566
rect 28028 17502 28030 17554
rect 28082 17502 28084 17554
rect 27356 16818 27412 16828
rect 27468 16882 27524 16894
rect 27468 16830 27470 16882
rect 27522 16830 27524 16882
rect 26796 15374 26798 15426
rect 26850 15374 26852 15426
rect 26796 15092 26852 15374
rect 26908 15764 26964 15774
rect 26908 15428 26964 15708
rect 27020 15538 27076 16268
rect 27468 15540 27524 16830
rect 27020 15486 27022 15538
rect 27074 15486 27076 15538
rect 27020 15474 27076 15486
rect 27356 15484 27524 15540
rect 27580 16772 27636 16782
rect 26908 15362 26964 15372
rect 27132 15428 27188 15438
rect 26572 14690 26628 14700
rect 26796 14532 26852 15036
rect 26460 13694 26462 13746
rect 26514 13694 26516 13746
rect 26460 13682 26516 13694
rect 26572 14476 26852 14532
rect 27020 15316 27076 15326
rect 26572 13858 26628 14476
rect 27020 14308 27076 15260
rect 27132 15204 27188 15372
rect 27356 15148 27412 15484
rect 27580 15426 27636 16716
rect 27804 16770 27860 16782
rect 27804 16718 27806 16770
rect 27858 16718 27860 16770
rect 27580 15374 27582 15426
rect 27634 15374 27636 15426
rect 27580 15362 27636 15374
rect 27692 16100 27748 16110
rect 27692 15428 27748 16044
rect 27692 15314 27748 15372
rect 27692 15262 27694 15314
rect 27746 15262 27748 15314
rect 27692 15250 27748 15262
rect 27132 15138 27188 15148
rect 27020 13860 27076 14252
rect 27244 15092 27412 15148
rect 27804 15204 27860 16718
rect 27916 16098 27972 16110
rect 27916 16046 27918 16098
rect 27970 16046 27972 16098
rect 27916 15316 27972 16046
rect 27916 15250 27972 15260
rect 27804 15138 27860 15148
rect 27132 13972 27188 13982
rect 27244 13972 27300 15092
rect 27804 14532 27860 14542
rect 28028 14532 28084 17502
rect 28252 17444 28308 17454
rect 28140 17442 28308 17444
rect 28140 17390 28254 17442
rect 28306 17390 28308 17442
rect 28140 17388 28308 17390
rect 28140 16324 28196 17388
rect 28252 17378 28308 17388
rect 28252 16996 28308 17006
rect 28364 16996 28420 17724
rect 28252 16994 28420 16996
rect 28252 16942 28254 16994
rect 28306 16942 28420 16994
rect 28252 16940 28420 16942
rect 28588 17444 28644 17454
rect 28252 16930 28308 16940
rect 28476 16884 28532 16894
rect 28476 16790 28532 16828
rect 28588 16660 28644 17388
rect 28140 15988 28196 16268
rect 28140 15922 28196 15932
rect 28476 16604 28644 16660
rect 28476 16098 28532 16604
rect 28476 16046 28478 16098
rect 28530 16046 28532 16098
rect 28364 15874 28420 15886
rect 28364 15822 28366 15874
rect 28418 15822 28420 15874
rect 28140 15540 28196 15550
rect 28140 15426 28196 15484
rect 28140 15374 28142 15426
rect 28194 15374 28196 15426
rect 28140 15362 28196 15374
rect 28364 14756 28420 15822
rect 28476 15764 28532 16046
rect 28476 15698 28532 15708
rect 28588 16324 28644 16334
rect 28588 15426 28644 16268
rect 28700 15876 28756 19068
rect 28812 18116 28868 21420
rect 28924 18452 28980 18462
rect 28924 18338 28980 18396
rect 28924 18286 28926 18338
rect 28978 18286 28980 18338
rect 28924 18274 28980 18286
rect 28812 18060 28980 18116
rect 28700 15810 28756 15820
rect 28812 16658 28868 16670
rect 28812 16606 28814 16658
rect 28866 16606 28868 16658
rect 28588 15374 28590 15426
rect 28642 15374 28644 15426
rect 28588 15362 28644 15374
rect 28812 15428 28868 16606
rect 28476 15316 28532 15326
rect 28476 15222 28532 15260
rect 28364 14690 28420 14700
rect 28588 15204 28644 15214
rect 28588 15090 28644 15148
rect 28588 15038 28590 15090
rect 28642 15038 28644 15090
rect 28252 14644 28308 14654
rect 28252 14550 28308 14588
rect 28140 14532 28196 14542
rect 27804 14438 27860 14476
rect 27916 14530 28196 14532
rect 27916 14478 28142 14530
rect 28194 14478 28196 14530
rect 27916 14476 28196 14478
rect 27916 14308 27972 14476
rect 28140 14466 28196 14476
rect 27188 13916 27300 13972
rect 27356 14252 27972 14308
rect 28028 14306 28084 14318
rect 28028 14254 28030 14306
rect 28082 14254 28084 14306
rect 27356 13970 27412 14252
rect 27356 13918 27358 13970
rect 27410 13918 27412 13970
rect 27132 13878 27188 13916
rect 27356 13906 27412 13918
rect 26572 13806 26574 13858
rect 26626 13806 26628 13858
rect 26572 13748 26628 13806
rect 26572 13682 26628 13692
rect 26684 13858 27076 13860
rect 26684 13806 27022 13858
rect 27074 13806 27076 13858
rect 26684 13804 27076 13806
rect 26684 13186 26740 13804
rect 27020 13794 27076 13804
rect 27132 13748 27188 13758
rect 26684 13134 26686 13186
rect 26738 13134 26740 13186
rect 26684 13122 26740 13134
rect 26908 13636 26964 13646
rect 25788 12910 25790 12962
rect 25842 12910 25844 12962
rect 25788 12898 25844 12910
rect 26124 13074 26180 13086
rect 26124 13022 26126 13074
rect 26178 13022 26180 13074
rect 26124 12740 26180 13022
rect 25676 12684 26180 12740
rect 26908 12964 26964 13580
rect 27020 12964 27076 12974
rect 26908 12962 27076 12964
rect 26908 12910 27022 12962
rect 27074 12910 27076 12962
rect 26908 12908 27076 12910
rect 26908 11954 26964 12908
rect 27020 12898 27076 12908
rect 27132 12852 27188 13692
rect 27244 12852 27300 12862
rect 27132 12796 27244 12852
rect 27020 12404 27076 12414
rect 27132 12404 27188 12796
rect 27244 12758 27300 12796
rect 27020 12402 27188 12404
rect 27020 12350 27022 12402
rect 27074 12350 27188 12402
rect 27020 12348 27188 12350
rect 27692 12738 27748 12750
rect 27692 12686 27694 12738
rect 27746 12686 27748 12738
rect 27020 12338 27076 12348
rect 26908 11902 26910 11954
rect 26962 11902 26964 11954
rect 26908 11890 26964 11902
rect 27468 12066 27524 12078
rect 27468 12014 27470 12066
rect 27522 12014 27524 12066
rect 27468 11956 27524 12014
rect 27692 11956 27748 12686
rect 27916 12180 27972 12190
rect 27916 12086 27972 12124
rect 27468 11954 27860 11956
rect 27468 11902 27470 11954
rect 27522 11902 27860 11954
rect 27468 11900 27860 11902
rect 27468 11862 27524 11900
rect 27692 11620 27748 11630
rect 27692 11526 27748 11564
rect 23996 11330 24052 11340
rect 24556 11508 24612 11518
rect 22764 11116 22932 11172
rect 23548 11282 23604 11294
rect 23548 11230 23550 11282
rect 23602 11230 23604 11282
rect 22764 10610 22820 11116
rect 23548 10836 23604 11230
rect 23996 11172 24052 11182
rect 23660 10836 23716 10846
rect 23548 10834 23716 10836
rect 23548 10782 23662 10834
rect 23714 10782 23716 10834
rect 23548 10780 23716 10782
rect 23660 10770 23716 10780
rect 23212 10724 23268 10734
rect 23268 10668 23492 10724
rect 23212 10630 23268 10668
rect 22764 10558 22766 10610
rect 22818 10558 22820 10610
rect 22764 10546 22820 10558
rect 22876 10610 22932 10622
rect 22876 10558 22878 10610
rect 22930 10558 22932 10610
rect 22764 9828 22820 9838
rect 22652 9826 22820 9828
rect 22652 9774 22766 9826
rect 22818 9774 22820 9826
rect 22652 9772 22820 9774
rect 22764 9716 22820 9772
rect 22764 9650 22820 9660
rect 22876 9268 22932 10558
rect 23436 10610 23492 10668
rect 23436 10558 23438 10610
rect 23490 10558 23492 10610
rect 23436 10546 23492 10558
rect 23772 10610 23828 10622
rect 23772 10558 23774 10610
rect 23826 10558 23828 10610
rect 23100 10498 23156 10510
rect 23100 10446 23102 10498
rect 23154 10446 23156 10498
rect 22652 9212 22932 9268
rect 22988 10052 23044 10062
rect 23100 10052 23156 10446
rect 23772 10388 23828 10558
rect 23996 10610 24052 11116
rect 24556 10722 24612 11452
rect 24556 10670 24558 10722
rect 24610 10670 24612 10722
rect 24556 10658 24612 10670
rect 25676 11508 25732 11518
rect 23996 10558 23998 10610
rect 24050 10558 24052 10610
rect 23996 10546 24052 10558
rect 24444 10388 24500 10398
rect 23772 10386 24500 10388
rect 23772 10334 24446 10386
rect 24498 10334 24500 10386
rect 23772 10332 24500 10334
rect 23100 9996 23492 10052
rect 22988 9268 23044 9996
rect 23436 9938 23492 9996
rect 23436 9886 23438 9938
rect 23490 9886 23492 9938
rect 23436 9874 23492 9886
rect 23100 9268 23156 9278
rect 22988 9266 23156 9268
rect 22988 9214 23102 9266
rect 23154 9214 23156 9266
rect 22988 9212 23156 9214
rect 22652 8820 22708 9212
rect 23100 9202 23156 9212
rect 23212 9044 23268 9054
rect 22988 9042 23268 9044
rect 22988 8990 23214 9042
rect 23266 8990 23268 9042
rect 22988 8988 23268 8990
rect 22652 8754 22708 8764
rect 22764 8932 22820 8942
rect 22988 8932 23044 8988
rect 23212 8978 23268 8988
rect 22764 8930 23044 8932
rect 22764 8878 22766 8930
rect 22818 8878 23044 8930
rect 22764 8876 23044 8878
rect 22540 8708 22596 8718
rect 22540 8370 22596 8652
rect 22764 8596 22820 8876
rect 22764 8530 22820 8540
rect 23324 8708 23380 8718
rect 22540 8318 22542 8370
rect 22594 8318 22596 8370
rect 22540 8306 22596 8318
rect 22876 8484 22932 8494
rect 22428 8206 22430 8258
rect 22482 8206 22484 8258
rect 22428 8194 22484 8206
rect 22876 8258 22932 8428
rect 22876 8206 22878 8258
rect 22930 8206 22932 8258
rect 22876 8194 22932 8206
rect 21980 8148 22036 8158
rect 21980 8146 22260 8148
rect 21980 8094 21982 8146
rect 22034 8094 22260 8146
rect 21980 8092 22260 8094
rect 21980 8082 22036 8092
rect 21644 7858 21700 7868
rect 22092 7588 22148 7598
rect 22092 7252 22148 7532
rect 22204 7476 22260 8092
rect 22540 8146 22596 8158
rect 22540 8094 22542 8146
rect 22594 8094 22596 8146
rect 22316 8036 22372 8046
rect 22316 7700 22372 7980
rect 22540 8036 22596 8094
rect 22540 7970 22596 7980
rect 22764 8036 22820 8074
rect 22764 7970 22820 7980
rect 23324 8036 23380 8652
rect 23772 8708 23828 10332
rect 24444 10322 24500 10332
rect 25564 9938 25620 9950
rect 25564 9886 25566 9938
rect 25618 9886 25620 9938
rect 25564 9492 25620 9886
rect 25340 9436 25620 9492
rect 24332 9156 24388 9166
rect 24332 9062 24388 9100
rect 25340 9156 25396 9436
rect 25452 9268 25508 9278
rect 25676 9268 25732 11452
rect 26572 11284 26628 11294
rect 26572 11190 26628 11228
rect 27356 11284 27412 11294
rect 27356 11190 27412 11228
rect 26908 11172 26964 11182
rect 26908 11170 27300 11172
rect 26908 11118 26910 11170
rect 26962 11118 27300 11170
rect 26908 11116 27300 11118
rect 26908 11106 26964 11116
rect 27244 10052 27300 11116
rect 27692 10612 27748 10622
rect 27692 10518 27748 10556
rect 27244 9996 27748 10052
rect 25452 9266 25732 9268
rect 25452 9214 25454 9266
rect 25506 9214 25732 9266
rect 25452 9212 25732 9214
rect 26908 9716 26964 9726
rect 25452 9202 25508 9212
rect 25340 9090 25396 9100
rect 25788 9156 25844 9166
rect 25788 9062 25844 9100
rect 25228 9042 25284 9054
rect 25228 8990 25230 9042
rect 25282 8990 25284 9042
rect 24220 8820 24276 8830
rect 24220 8726 24276 8764
rect 23772 8642 23828 8652
rect 23324 7970 23380 7980
rect 25116 8260 25172 8270
rect 22764 7812 22820 7822
rect 22652 7700 22708 7710
rect 22316 7698 22708 7700
rect 22316 7646 22654 7698
rect 22706 7646 22708 7698
rect 22316 7644 22708 7646
rect 22652 7634 22708 7644
rect 22316 7476 22372 7486
rect 22204 7420 22316 7476
rect 22316 7382 22372 7420
rect 22764 7362 22820 7756
rect 24668 7700 24724 7710
rect 24668 7606 24724 7644
rect 22764 7310 22766 7362
rect 22818 7310 22820 7362
rect 22204 7252 22260 7262
rect 21868 7250 22260 7252
rect 21868 7198 22206 7250
rect 22258 7198 22260 7250
rect 21868 7196 22260 7198
rect 21420 6692 21476 6702
rect 21420 6598 21476 6636
rect 21868 6690 21924 7196
rect 22204 7186 22260 7196
rect 21868 6638 21870 6690
rect 21922 6638 21924 6690
rect 21868 6626 21924 6638
rect 22764 6692 22820 7310
rect 24556 7588 24612 7598
rect 24556 6804 24612 7532
rect 24892 7476 24948 7486
rect 24892 6914 24948 7420
rect 24892 6862 24894 6914
rect 24946 6862 24948 6914
rect 24892 6850 24948 6862
rect 24556 6738 24612 6748
rect 22428 6580 22484 6590
rect 20748 5854 20750 5906
rect 20802 5854 20804 5906
rect 20748 5842 20804 5854
rect 20860 6020 20916 6030
rect 18844 4946 18900 4956
rect 19292 5794 19348 5806
rect 19292 5742 19294 5794
rect 19346 5742 19348 5794
rect 19068 4452 19124 4462
rect 18396 4450 19124 4452
rect 18396 4398 19070 4450
rect 19122 4398 19124 4450
rect 18396 4396 19124 4398
rect 19068 4386 19124 4396
rect 19292 4452 19348 5742
rect 20860 5346 20916 5964
rect 20860 5294 20862 5346
rect 20914 5294 20916 5346
rect 20860 5282 20916 5294
rect 22428 6020 22484 6524
rect 22764 6132 22820 6636
rect 25116 6690 25172 8204
rect 25228 7700 25284 8990
rect 25676 9042 25732 9054
rect 25676 8990 25678 9042
rect 25730 8990 25732 9042
rect 25676 8482 25732 8990
rect 26908 9042 26964 9660
rect 27692 9154 27748 9996
rect 27804 9380 27860 11900
rect 28028 11396 28084 14254
rect 28364 13972 28420 13982
rect 28364 13746 28420 13916
rect 28364 13694 28366 13746
rect 28418 13694 28420 13746
rect 28364 13682 28420 13694
rect 28588 13746 28644 15038
rect 28812 14644 28868 15372
rect 28924 15148 28980 18060
rect 29036 16772 29092 21532
rect 29148 21522 29204 21532
rect 29148 21362 29204 21374
rect 29148 21310 29150 21362
rect 29202 21310 29204 21362
rect 29148 20468 29204 21310
rect 29260 20692 29316 20702
rect 29260 20598 29316 20636
rect 29148 20402 29204 20412
rect 29372 20356 29428 23548
rect 29596 22482 29652 23886
rect 30044 23938 30100 24780
rect 30044 23886 30046 23938
rect 30098 23886 30100 23938
rect 30044 23874 30100 23886
rect 30828 23826 30884 23838
rect 30828 23774 30830 23826
rect 30882 23774 30884 23826
rect 30828 23378 30884 23774
rect 30828 23326 30830 23378
rect 30882 23326 30884 23378
rect 30828 23314 30884 23326
rect 31612 23380 31668 23390
rect 30380 23268 30436 23278
rect 30044 23156 30100 23166
rect 29596 22430 29598 22482
rect 29650 22430 29652 22482
rect 29596 22418 29652 22430
rect 29708 23042 29764 23054
rect 29708 22990 29710 23042
rect 29762 22990 29764 23042
rect 29484 22260 29540 22270
rect 29484 22166 29540 22204
rect 29708 22146 29764 22990
rect 30044 22930 30100 23100
rect 30380 23154 30436 23212
rect 31052 23268 31108 23278
rect 31052 23174 31108 23212
rect 30380 23102 30382 23154
rect 30434 23102 30436 23154
rect 30380 23090 30436 23102
rect 30604 23156 30660 23166
rect 30604 23062 30660 23100
rect 31164 23154 31220 23166
rect 31164 23102 31166 23154
rect 31218 23102 31220 23154
rect 30044 22878 30046 22930
rect 30098 22878 30100 22930
rect 30044 22260 30100 22878
rect 30380 22932 30436 22942
rect 31164 22932 31220 23102
rect 31612 23044 31668 23324
rect 31612 22978 31668 22988
rect 31724 23156 31780 25228
rect 31836 24612 31892 24622
rect 32172 24612 32228 24622
rect 31836 24610 32228 24612
rect 31836 24558 31838 24610
rect 31890 24558 32174 24610
rect 32226 24558 32228 24610
rect 31836 24556 32228 24558
rect 31836 24546 31892 24556
rect 32172 24546 32228 24556
rect 32284 24498 32340 24510
rect 32284 24446 32286 24498
rect 32338 24446 32340 24498
rect 32284 23940 32340 24446
rect 32284 23874 32340 23884
rect 32396 23380 32452 27022
rect 32396 23314 32452 23324
rect 30380 22930 31220 22932
rect 30380 22878 30382 22930
rect 30434 22878 31220 22930
rect 30380 22876 31220 22878
rect 30380 22866 30436 22876
rect 30268 22372 30324 22382
rect 30268 22370 30436 22372
rect 30268 22318 30270 22370
rect 30322 22318 30436 22370
rect 30268 22316 30436 22318
rect 30268 22306 30324 22316
rect 30044 22194 30100 22204
rect 29708 22094 29710 22146
rect 29762 22094 29764 22146
rect 29596 21474 29652 21486
rect 29596 21422 29598 21474
rect 29650 21422 29652 21474
rect 29596 21362 29652 21422
rect 29596 21310 29598 21362
rect 29650 21310 29652 21362
rect 29596 21298 29652 21310
rect 29484 20692 29540 20702
rect 29484 20598 29540 20636
rect 29372 20290 29428 20300
rect 29596 20578 29652 20590
rect 29596 20526 29598 20578
rect 29650 20526 29652 20578
rect 29260 20244 29316 20254
rect 29148 20132 29204 20142
rect 29148 19796 29204 20076
rect 29260 20130 29316 20188
rect 29596 20244 29652 20526
rect 29596 20178 29652 20188
rect 29260 20078 29262 20130
rect 29314 20078 29316 20130
rect 29260 20066 29316 20078
rect 29148 19740 29316 19796
rect 29148 19236 29204 19246
rect 29148 19142 29204 19180
rect 29260 18450 29316 19740
rect 29708 19012 29764 22094
rect 29820 20804 29876 20814
rect 30044 20804 30100 20814
rect 29820 20802 30100 20804
rect 29820 20750 29822 20802
rect 29874 20750 30046 20802
rect 30098 20750 30100 20802
rect 29820 20748 30100 20750
rect 29820 20132 29876 20748
rect 30044 20738 30100 20748
rect 30268 20578 30324 20590
rect 30268 20526 30270 20578
rect 30322 20526 30324 20578
rect 30268 20244 30324 20526
rect 29820 20066 29876 20076
rect 29932 20188 30324 20244
rect 29932 19346 29988 20188
rect 30380 20132 30436 22316
rect 30940 22258 30996 22270
rect 30940 22206 30942 22258
rect 30994 22206 30996 22258
rect 30940 21810 30996 22206
rect 31724 21812 31780 23100
rect 31836 23154 31892 23166
rect 31836 23102 31838 23154
rect 31890 23102 31892 23154
rect 31836 22036 31892 23102
rect 32396 23156 32452 23166
rect 32396 23062 32452 23100
rect 31836 21970 31892 21980
rect 31948 22484 32004 22494
rect 31948 21812 32004 22428
rect 30940 21758 30942 21810
rect 30994 21758 30996 21810
rect 30940 21746 30996 21758
rect 31612 21756 31780 21812
rect 31836 21756 32004 21812
rect 30828 21588 30884 21598
rect 30604 20802 30660 20814
rect 30604 20750 30606 20802
rect 30658 20750 30660 20802
rect 29932 19294 29934 19346
rect 29986 19294 29988 19346
rect 29932 19282 29988 19294
rect 30044 20076 30436 20132
rect 30492 20690 30548 20702
rect 30492 20638 30494 20690
rect 30546 20638 30548 20690
rect 30044 19236 30100 20076
rect 30492 20020 30548 20638
rect 30492 19954 30548 19964
rect 30044 19170 30100 19180
rect 30156 19796 30212 19806
rect 29708 18946 29764 18956
rect 30156 19124 30212 19740
rect 29596 18676 29652 18686
rect 29260 18398 29262 18450
rect 29314 18398 29316 18450
rect 29260 18386 29316 18398
rect 29484 18562 29540 18574
rect 29484 18510 29486 18562
rect 29538 18510 29540 18562
rect 29484 18340 29540 18510
rect 29484 18004 29540 18284
rect 29596 18338 29652 18620
rect 29596 18286 29598 18338
rect 29650 18286 29652 18338
rect 29596 18274 29652 18286
rect 29932 18562 29988 18574
rect 29932 18510 29934 18562
rect 29986 18510 29988 18562
rect 29932 18228 29988 18510
rect 30156 18450 30212 19068
rect 30604 18676 30660 20750
rect 30604 18610 30660 18620
rect 30156 18398 30158 18450
rect 30210 18398 30212 18450
rect 30156 18386 30212 18398
rect 30716 18340 30772 18350
rect 30716 18246 30772 18284
rect 29932 18162 29988 18172
rect 29484 17948 29876 18004
rect 29372 17444 29428 17454
rect 29372 17350 29428 17388
rect 29148 16772 29204 16782
rect 29036 16716 29148 16772
rect 29148 16706 29204 16716
rect 29484 16772 29540 16782
rect 29540 16716 29652 16772
rect 29484 16678 29540 16716
rect 29148 16548 29204 16558
rect 29148 16322 29204 16492
rect 29148 16270 29150 16322
rect 29202 16270 29204 16322
rect 29148 16258 29204 16270
rect 29484 16100 29540 16110
rect 29484 16006 29540 16044
rect 29372 15316 29428 15326
rect 29372 15204 29428 15260
rect 29484 15204 29540 15214
rect 29372 15202 29540 15204
rect 29372 15150 29486 15202
rect 29538 15150 29540 15202
rect 29372 15148 29540 15150
rect 28924 15092 29092 15148
rect 29484 15138 29540 15148
rect 29036 14868 29092 15092
rect 29036 14812 29316 14868
rect 28868 14588 29092 14644
rect 28812 14578 28868 14588
rect 28700 13972 28756 13982
rect 28700 13970 28980 13972
rect 28700 13918 28702 13970
rect 28754 13918 28980 13970
rect 28700 13916 28980 13918
rect 28700 13906 28756 13916
rect 28588 13694 28590 13746
rect 28642 13694 28644 13746
rect 28588 13682 28644 13694
rect 28812 13076 28868 13086
rect 28140 12852 28196 12862
rect 28140 12740 28196 12796
rect 28588 12740 28644 12750
rect 28140 12738 28644 12740
rect 28140 12686 28142 12738
rect 28194 12686 28590 12738
rect 28642 12686 28644 12738
rect 28140 12684 28644 12686
rect 28140 12674 28196 12684
rect 28588 12628 28644 12684
rect 28588 12562 28644 12572
rect 28140 12292 28196 12302
rect 28812 12292 28868 13020
rect 28924 12404 28980 13916
rect 29036 13860 29092 14588
rect 29148 14532 29204 14542
rect 29148 14438 29204 14476
rect 29260 14420 29316 14812
rect 29260 14418 29428 14420
rect 29260 14366 29262 14418
rect 29314 14366 29428 14418
rect 29260 14364 29428 14366
rect 29260 14354 29316 14364
rect 29148 13860 29204 13870
rect 29036 13858 29204 13860
rect 29036 13806 29150 13858
rect 29202 13806 29204 13858
rect 29036 13804 29204 13806
rect 29148 13794 29204 13804
rect 29372 13074 29428 14364
rect 29596 14196 29652 16716
rect 29708 16212 29764 16222
rect 29708 16118 29764 16156
rect 29596 14130 29652 14140
rect 29820 13412 29876 17948
rect 30828 17108 30884 21532
rect 31276 21588 31332 21598
rect 31276 21586 31556 21588
rect 31276 21534 31278 21586
rect 31330 21534 31556 21586
rect 31276 21532 31556 21534
rect 31276 21522 31332 21532
rect 31500 21026 31556 21532
rect 31500 20974 31502 21026
rect 31554 20974 31556 21026
rect 31500 20962 31556 20974
rect 31612 20804 31668 21756
rect 31724 21588 31780 21598
rect 31724 21494 31780 21532
rect 31836 21026 31892 21756
rect 31836 20974 31838 21026
rect 31890 20974 31892 21026
rect 31836 20962 31892 20974
rect 32396 21588 32452 21598
rect 31612 20748 31892 20804
rect 31724 20130 31780 20142
rect 31724 20078 31726 20130
rect 31778 20078 31780 20130
rect 31052 20020 31108 20030
rect 31052 18450 31108 19964
rect 31388 19908 31444 19918
rect 31388 19814 31444 19852
rect 31052 18398 31054 18450
rect 31106 18398 31108 18450
rect 31052 18386 31108 18398
rect 31164 19348 31220 19358
rect 31164 18450 31220 19292
rect 31164 18398 31166 18450
rect 31218 18398 31220 18450
rect 31164 18386 31220 18398
rect 31724 18340 31780 20078
rect 31724 18274 31780 18284
rect 31836 18452 31892 20748
rect 32284 20802 32340 20814
rect 32284 20750 32286 20802
rect 32338 20750 32340 20802
rect 32060 20132 32116 20142
rect 32060 20038 32116 20076
rect 32060 19348 32116 19358
rect 32060 19254 32116 19292
rect 32284 18900 32340 20750
rect 32396 20690 32452 21532
rect 32396 20638 32398 20690
rect 32450 20638 32452 20690
rect 32396 20626 32452 20638
rect 32508 20692 32564 20702
rect 32508 20130 32564 20636
rect 32508 20078 32510 20130
rect 32562 20078 32564 20130
rect 32508 20066 32564 20078
rect 32396 19908 32452 19918
rect 32396 19814 32452 19852
rect 32508 19122 32564 19134
rect 32508 19070 32510 19122
rect 32562 19070 32564 19122
rect 32508 18900 32564 19070
rect 32284 18844 32564 18900
rect 32172 18452 32228 18462
rect 32284 18452 32340 18844
rect 31836 18450 32116 18452
rect 31836 18398 31838 18450
rect 31890 18398 32116 18450
rect 31836 18396 32116 18398
rect 31164 17444 31220 17454
rect 30884 17052 30996 17108
rect 30828 17014 30884 17052
rect 29932 16884 29988 16894
rect 29932 16790 29988 16828
rect 30716 16884 30772 16894
rect 30604 16212 30660 16222
rect 30044 15988 30100 15998
rect 30044 15894 30100 15932
rect 30380 15876 30436 15886
rect 30156 15820 30380 15876
rect 30044 15540 30100 15550
rect 30156 15540 30212 15820
rect 30380 15782 30436 15820
rect 30044 15538 30212 15540
rect 30044 15486 30046 15538
rect 30098 15486 30212 15538
rect 30044 15484 30212 15486
rect 30604 15538 30660 16156
rect 30716 15874 30772 16828
rect 30716 15822 30718 15874
rect 30770 15822 30772 15874
rect 30716 15764 30772 15822
rect 30716 15698 30772 15708
rect 30828 16324 30884 16334
rect 30604 15486 30606 15538
rect 30658 15486 30660 15538
rect 30044 15474 30100 15484
rect 30604 15474 30660 15486
rect 30380 15428 30436 15438
rect 30380 15334 30436 15372
rect 29820 13346 29876 13356
rect 30044 15316 30100 15326
rect 29372 13022 29374 13074
rect 29426 13022 29428 13074
rect 29372 13010 29428 13022
rect 30044 13076 30100 15260
rect 30492 15202 30548 15214
rect 30492 15150 30494 15202
rect 30546 15150 30548 15202
rect 30268 14308 30324 14318
rect 30268 14214 30324 14252
rect 30492 14306 30548 15150
rect 30604 14530 30660 14542
rect 30604 14478 30606 14530
rect 30658 14478 30660 14530
rect 30604 14418 30660 14478
rect 30604 14366 30606 14418
rect 30658 14366 30660 14418
rect 30604 14354 30660 14366
rect 30716 14532 30772 14542
rect 30492 14254 30494 14306
rect 30546 14254 30548 14306
rect 30492 14242 30548 14254
rect 30492 13860 30548 13870
rect 30044 12982 30100 13020
rect 30268 13858 30548 13860
rect 30268 13806 30494 13858
rect 30546 13806 30548 13858
rect 30268 13804 30548 13806
rect 28924 12348 29204 12404
rect 28140 12290 28420 12292
rect 28140 12238 28142 12290
rect 28194 12238 28420 12290
rect 28140 12236 28420 12238
rect 28140 12226 28196 12236
rect 28028 11282 28084 11340
rect 28028 11230 28030 11282
rect 28082 11230 28084 11282
rect 28028 11218 28084 11230
rect 28364 10722 28420 12236
rect 28588 12180 28644 12190
rect 28812 12180 28868 12236
rect 28924 12180 28980 12190
rect 28812 12178 28980 12180
rect 28812 12126 28926 12178
rect 28978 12126 28980 12178
rect 28812 12124 28980 12126
rect 28588 12086 28644 12124
rect 28924 12114 28980 12124
rect 28364 10670 28366 10722
rect 28418 10670 28420 10722
rect 28364 10658 28420 10670
rect 28476 11282 28532 11294
rect 28476 11230 28478 11282
rect 28530 11230 28532 11282
rect 27804 9314 27860 9324
rect 27692 9102 27694 9154
rect 27746 9102 27748 9154
rect 27692 9090 27748 9102
rect 26908 8990 26910 9042
rect 26962 8990 26964 9042
rect 26908 8978 26964 8990
rect 25676 8430 25678 8482
rect 25730 8430 25732 8482
rect 25564 8260 25620 8270
rect 25564 8166 25620 8204
rect 25284 7644 25620 7700
rect 25228 7634 25284 7644
rect 25228 7476 25284 7486
rect 25228 7382 25284 7420
rect 25116 6638 25118 6690
rect 25170 6638 25172 6690
rect 25116 6626 25172 6638
rect 25564 6690 25620 7644
rect 25676 7474 25732 8430
rect 25788 8930 25844 8942
rect 25788 8878 25790 8930
rect 25842 8878 25844 8930
rect 25788 8148 25844 8878
rect 28476 8932 28532 11230
rect 29036 9156 29092 12348
rect 29148 12290 29204 12348
rect 30268 12402 30324 13804
rect 30492 13794 30548 13804
rect 30268 12350 30270 12402
rect 30322 12350 30324 12402
rect 29148 12238 29150 12290
rect 29202 12238 29204 12290
rect 29148 12226 29204 12238
rect 29708 12292 29764 12302
rect 29708 12290 30100 12292
rect 29708 12238 29710 12290
rect 29762 12238 30100 12290
rect 29708 12236 30100 12238
rect 29708 12226 29764 12236
rect 29820 11396 29876 11406
rect 29820 11302 29876 11340
rect 29484 11284 29540 11294
rect 29484 11190 29540 11228
rect 29036 9090 29092 9100
rect 29148 11170 29204 11182
rect 29148 11118 29150 11170
rect 29202 11118 29204 11170
rect 29148 10612 29204 11118
rect 30044 10948 30100 12236
rect 30268 11620 30324 12350
rect 30604 12404 30660 12414
rect 30716 12404 30772 14476
rect 30828 13972 30884 16268
rect 30940 15428 30996 17052
rect 31052 15874 31108 15886
rect 31052 15822 31054 15874
rect 31106 15822 31108 15874
rect 31052 15652 31108 15822
rect 31052 15586 31108 15596
rect 30940 15362 30996 15372
rect 30940 14532 30996 14542
rect 31164 14532 31220 17388
rect 31612 15876 31668 15886
rect 31612 15782 31668 15820
rect 31388 15652 31444 15662
rect 31444 15596 31556 15652
rect 31388 15586 31444 15596
rect 30940 14530 31220 14532
rect 30940 14478 30942 14530
rect 30994 14478 31166 14530
rect 31218 14478 31220 14530
rect 30940 14476 31220 14478
rect 30940 14466 30996 14476
rect 31164 14466 31220 14476
rect 31276 15540 31332 15550
rect 31276 15314 31332 15484
rect 31388 15428 31444 15438
rect 31388 15334 31444 15372
rect 31276 15262 31278 15314
rect 31330 15262 31332 15314
rect 31276 13972 31332 15262
rect 31500 15148 31556 15596
rect 31836 15148 31892 18396
rect 32060 18228 32116 18396
rect 32228 18396 32340 18452
rect 32396 18562 32452 18574
rect 32396 18510 32398 18562
rect 32450 18510 32452 18562
rect 32172 18358 32228 18396
rect 32396 18228 32452 18510
rect 32508 18340 32564 18350
rect 32508 18246 32564 18284
rect 32060 18172 32452 18228
rect 32620 18228 32676 30940
rect 32956 30212 33012 30222
rect 33068 30212 33124 31052
rect 35084 31042 35140 31052
rect 33292 30996 33348 31006
rect 33292 30902 33348 30940
rect 34076 30884 34132 30894
rect 33740 30436 33796 30446
rect 33740 30342 33796 30380
rect 33404 30324 33460 30334
rect 33628 30324 33684 30334
rect 33404 30230 33460 30268
rect 33516 30268 33628 30324
rect 32844 30210 33124 30212
rect 32844 30158 32958 30210
rect 33010 30158 33124 30210
rect 32844 30156 33124 30158
rect 32732 29986 32788 29998
rect 32732 29934 32734 29986
rect 32786 29934 32788 29986
rect 32732 29764 32788 29934
rect 32732 29698 32788 29708
rect 32844 20804 32900 30156
rect 32956 30146 33012 30156
rect 33068 29540 33124 29550
rect 33068 29446 33124 29484
rect 33404 29428 33460 29438
rect 33516 29428 33572 30268
rect 33628 30258 33684 30268
rect 34076 30098 34132 30828
rect 35196 30772 35252 31892
rect 35084 30716 35252 30772
rect 35308 31892 35588 31948
rect 35644 31892 35700 31902
rect 35756 31892 35812 33516
rect 35868 33460 35924 34750
rect 35980 34916 36036 34926
rect 35980 34018 36036 34860
rect 36092 34914 36148 34926
rect 36092 34862 36094 34914
rect 36146 34862 36148 34914
rect 36092 34580 36148 34862
rect 36204 34914 36260 34926
rect 36204 34862 36206 34914
rect 36258 34862 36260 34914
rect 36204 34692 36260 34862
rect 36428 34916 36484 35422
rect 37100 35474 37156 35486
rect 37100 35422 37102 35474
rect 37154 35422 37156 35474
rect 36428 34850 36484 34860
rect 36988 35028 37044 35038
rect 36988 34804 37044 34972
rect 36204 34626 36260 34636
rect 36652 34802 37044 34804
rect 36652 34750 36990 34802
rect 37042 34750 37044 34802
rect 36652 34748 37044 34750
rect 36092 34514 36148 34524
rect 36204 34468 36260 34478
rect 36204 34356 36260 34412
rect 35980 33966 35982 34018
rect 36034 33966 36036 34018
rect 35980 33954 36036 33966
rect 36092 34300 36260 34356
rect 36092 33796 36148 34300
rect 36652 34242 36708 34748
rect 36988 34738 37044 34748
rect 37100 34804 37156 35422
rect 37100 34738 37156 34748
rect 37212 34580 37268 35868
rect 37436 35700 37492 37436
rect 38108 37380 38164 38556
rect 38220 38164 38276 38894
rect 38220 38098 38276 38108
rect 38444 38948 38500 38958
rect 38444 38836 38500 38892
rect 38780 38946 38836 39004
rect 38892 38994 38948 39004
rect 38780 38894 38782 38946
rect 38834 38894 38836 38946
rect 38780 38882 38836 38894
rect 38556 38836 38612 38846
rect 38444 38834 38612 38836
rect 38444 38782 38558 38834
rect 38610 38782 38612 38834
rect 38444 38780 38612 38782
rect 37884 37324 38164 37380
rect 38444 37380 38500 38780
rect 38556 38770 38612 38780
rect 39228 38836 39284 38846
rect 39228 38742 39284 38780
rect 38780 38724 38836 38734
rect 39564 38724 39620 39452
rect 39900 39172 39956 40350
rect 39900 39106 39956 39116
rect 39788 39060 39844 39070
rect 39788 38966 39844 39004
rect 39676 38948 39732 38958
rect 39676 38854 39732 38892
rect 40012 38836 40068 38846
rect 39788 38834 40068 38836
rect 39788 38782 40014 38834
rect 40066 38782 40068 38834
rect 39788 38780 40068 38782
rect 39676 38724 39732 38734
rect 39564 38722 39732 38724
rect 39564 38670 39678 38722
rect 39730 38670 39732 38722
rect 39564 38668 39732 38670
rect 38444 37378 38724 37380
rect 38444 37326 38446 37378
rect 38498 37326 38724 37378
rect 38444 37324 38724 37326
rect 37660 37266 37716 37278
rect 37660 37214 37662 37266
rect 37714 37214 37716 37266
rect 37660 37156 37716 37214
rect 37660 37090 37716 37100
rect 37548 37042 37604 37054
rect 37548 36990 37550 37042
rect 37602 36990 37604 37042
rect 37548 36260 37604 36990
rect 37884 36482 37940 37324
rect 38444 37314 38500 37324
rect 38220 37268 38276 37278
rect 38220 37174 38276 37212
rect 38332 37154 38388 37166
rect 38332 37102 38334 37154
rect 38386 37102 38388 37154
rect 37996 37044 38052 37054
rect 37996 37042 38276 37044
rect 37996 36990 37998 37042
rect 38050 36990 38276 37042
rect 37996 36988 38276 36990
rect 37996 36978 38052 36988
rect 37884 36430 37886 36482
rect 37938 36430 37940 36482
rect 37884 36418 37940 36430
rect 37548 36204 37940 36260
rect 37660 35924 37716 35934
rect 37492 35644 37604 35700
rect 37436 35606 37492 35644
rect 37548 34804 37604 35644
rect 37660 35698 37716 35868
rect 37660 35646 37662 35698
rect 37714 35646 37716 35698
rect 37660 35634 37716 35646
rect 37660 34804 37716 34814
rect 37548 34802 37716 34804
rect 37548 34750 37662 34802
rect 37714 34750 37716 34802
rect 37548 34748 37716 34750
rect 36652 34190 36654 34242
rect 36706 34190 36708 34242
rect 36428 34130 36484 34142
rect 36428 34078 36430 34130
rect 36482 34078 36484 34130
rect 35868 33234 35924 33404
rect 35868 33182 35870 33234
rect 35922 33182 35924 33234
rect 35868 33170 35924 33182
rect 35980 33740 36148 33796
rect 36204 34020 36260 34030
rect 35980 33124 36036 33740
rect 36092 33348 36148 33358
rect 36204 33348 36260 33964
rect 36092 33346 36260 33348
rect 36092 33294 36094 33346
rect 36146 33294 36260 33346
rect 36092 33292 36260 33294
rect 36316 33684 36372 33694
rect 36092 33282 36148 33292
rect 36204 33124 36260 33134
rect 35980 33068 36148 33124
rect 35980 32676 36036 32686
rect 36092 32676 36148 33068
rect 36316 33124 36372 33628
rect 36428 33572 36484 34078
rect 36540 34132 36596 34142
rect 36540 34038 36596 34076
rect 36652 34020 36708 34190
rect 36988 34524 37268 34580
rect 37324 34690 37380 34702
rect 37324 34638 37326 34690
rect 37378 34638 37380 34690
rect 36988 34242 37044 34524
rect 36988 34190 36990 34242
rect 37042 34190 37044 34242
rect 36988 34178 37044 34190
rect 36652 33954 36708 33964
rect 37100 33572 37156 34524
rect 37324 34468 37380 34638
rect 37324 34402 37380 34412
rect 37548 34244 37604 34748
rect 37660 34738 37716 34748
rect 37212 34188 37604 34244
rect 37772 34692 37828 34702
rect 37772 34242 37828 34636
rect 37772 34190 37774 34242
rect 37826 34190 37828 34242
rect 37212 34130 37268 34188
rect 37772 34178 37828 34190
rect 37212 34078 37214 34130
rect 37266 34078 37268 34130
rect 37212 34066 37268 34078
rect 37324 33908 37380 33918
rect 37324 33814 37380 33852
rect 37660 33906 37716 33918
rect 37660 33854 37662 33906
rect 37714 33854 37716 33906
rect 37660 33684 37716 33854
rect 37660 33618 37716 33628
rect 37100 33516 37604 33572
rect 36428 33506 36484 33516
rect 36428 33348 36484 33358
rect 37100 33348 37156 33358
rect 36428 33346 36932 33348
rect 36428 33294 36430 33346
rect 36482 33294 36932 33346
rect 36428 33292 36932 33294
rect 36428 33282 36484 33292
rect 36316 33068 36484 33124
rect 36204 33030 36260 33068
rect 36204 32676 36260 32686
rect 36092 32674 36260 32676
rect 36092 32622 36206 32674
rect 36258 32622 36260 32674
rect 36092 32620 36260 32622
rect 35980 32582 36036 32620
rect 36204 32610 36260 32620
rect 36428 32674 36484 33068
rect 36876 32786 36932 33292
rect 37100 33346 37492 33348
rect 37100 33294 37102 33346
rect 37154 33294 37492 33346
rect 37100 33292 37492 33294
rect 37100 33282 37156 33292
rect 37436 33236 37492 33292
rect 37324 33124 37380 33134
rect 36876 32734 36878 32786
rect 36930 32734 36932 32786
rect 36428 32622 36430 32674
rect 36482 32622 36484 32674
rect 36428 32610 36484 32622
rect 36764 32676 36820 32686
rect 36764 32582 36820 32620
rect 36316 32562 36372 32574
rect 36316 32510 36318 32562
rect 36370 32510 36372 32562
rect 36316 32452 36372 32510
rect 36316 32386 36372 32396
rect 35308 30772 35364 31836
rect 35644 31890 35812 31892
rect 35644 31838 35646 31890
rect 35698 31838 35812 31890
rect 35644 31836 35812 31838
rect 35644 31826 35700 31836
rect 35420 31108 35476 31118
rect 35420 31106 35588 31108
rect 35420 31054 35422 31106
rect 35474 31054 35588 31106
rect 35420 31052 35588 31054
rect 35420 31042 35476 31052
rect 35084 30324 35140 30716
rect 35308 30706 35364 30716
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34076 30046 34078 30098
rect 34130 30046 34132 30098
rect 34076 30034 34132 30046
rect 34300 30210 34356 30222
rect 34300 30158 34302 30210
rect 34354 30158 34356 30210
rect 33628 29988 33684 29998
rect 33628 29894 33684 29932
rect 34300 29988 34356 30158
rect 35084 30098 35140 30268
rect 35084 30046 35086 30098
rect 35138 30046 35140 30098
rect 35084 30034 35140 30046
rect 34748 29988 34804 29998
rect 34300 29986 34804 29988
rect 34300 29934 34750 29986
rect 34802 29934 34804 29986
rect 34300 29932 34804 29934
rect 34188 29652 34244 29662
rect 34300 29652 34356 29932
rect 34748 29922 34804 29932
rect 34244 29596 34356 29652
rect 34188 29558 34244 29596
rect 35420 29540 35476 29550
rect 35532 29540 35588 31052
rect 35420 29538 35588 29540
rect 35420 29486 35422 29538
rect 35474 29486 35588 29538
rect 35420 29484 35588 29486
rect 35756 30994 35812 31006
rect 35756 30942 35758 30994
rect 35810 30942 35812 30994
rect 35420 29474 35476 29484
rect 33404 29426 33572 29428
rect 33404 29374 33406 29426
rect 33458 29374 33572 29426
rect 33404 29372 33572 29374
rect 34748 29428 34804 29438
rect 33404 29362 33460 29372
rect 34748 29334 34804 29372
rect 35756 29428 35812 30942
rect 36540 30882 36596 30894
rect 36540 30830 36542 30882
rect 36594 30830 36596 30882
rect 36540 30100 36596 30830
rect 36876 30660 36932 32734
rect 37212 33122 37380 33124
rect 37212 33070 37326 33122
rect 37378 33070 37380 33122
rect 37212 33068 37380 33070
rect 37100 32562 37156 32574
rect 37100 32510 37102 32562
rect 37154 32510 37156 32562
rect 37100 32004 37156 32510
rect 36876 30594 36932 30604
rect 36988 31554 37044 31566
rect 36988 31502 36990 31554
rect 37042 31502 37044 31554
rect 36988 30884 37044 31502
rect 37100 31556 37156 31948
rect 37212 31892 37268 33068
rect 37324 33058 37380 33068
rect 37436 32562 37492 33180
rect 37436 32510 37438 32562
rect 37490 32510 37492 32562
rect 37436 32498 37492 32510
rect 37548 32788 37604 33516
rect 37660 33460 37716 33470
rect 37660 33234 37716 33404
rect 37660 33182 37662 33234
rect 37714 33182 37716 33234
rect 37660 33170 37716 33182
rect 37660 32788 37716 32798
rect 37548 32786 37716 32788
rect 37548 32734 37662 32786
rect 37714 32734 37716 32786
rect 37548 32732 37716 32734
rect 37548 32340 37604 32732
rect 37660 32722 37716 32732
rect 37884 32564 37940 36204
rect 38220 35140 38276 36988
rect 38332 36596 38388 37102
rect 38668 36820 38724 37324
rect 38780 37378 38836 38668
rect 39676 38658 39732 38668
rect 39116 38612 39172 38622
rect 39116 37490 39172 38556
rect 39116 37438 39118 37490
rect 39170 37438 39172 37490
rect 39116 37426 39172 37438
rect 38780 37326 38782 37378
rect 38834 37326 38836 37378
rect 38780 37314 38836 37326
rect 39452 37268 39508 37278
rect 39676 37268 39732 37278
rect 39452 37174 39508 37212
rect 39564 37212 39676 37268
rect 39564 37154 39620 37212
rect 39676 37202 39732 37212
rect 39564 37102 39566 37154
rect 39618 37102 39620 37154
rect 39564 37090 39620 37102
rect 38668 36764 38836 36820
rect 38668 36596 38724 36606
rect 38332 36594 38724 36596
rect 38332 36542 38670 36594
rect 38722 36542 38724 36594
rect 38332 36540 38724 36542
rect 38668 36530 38724 36540
rect 38780 35924 38836 36764
rect 39340 35924 39396 35934
rect 38780 35922 39396 35924
rect 38780 35870 39342 35922
rect 39394 35870 39396 35922
rect 38780 35868 39396 35870
rect 38780 35698 38836 35868
rect 39340 35858 39396 35868
rect 38780 35646 38782 35698
rect 38834 35646 38836 35698
rect 38780 35634 38836 35646
rect 39004 35700 39060 35710
rect 39004 35606 39060 35644
rect 39564 35698 39620 35710
rect 39564 35646 39566 35698
rect 39618 35646 39620 35698
rect 38332 35140 38388 35150
rect 38220 35138 38388 35140
rect 38220 35086 38334 35138
rect 38386 35086 38388 35138
rect 38220 35084 38388 35086
rect 38332 35074 38388 35084
rect 38332 34914 38388 34926
rect 38332 34862 38334 34914
rect 38386 34862 38388 34914
rect 37996 34692 38052 34702
rect 37996 34690 38164 34692
rect 37996 34638 37998 34690
rect 38050 34638 38164 34690
rect 37996 34636 38164 34638
rect 37996 34626 38052 34636
rect 38108 34580 38164 34636
rect 38108 33348 38164 34524
rect 38332 33908 38388 34862
rect 38668 34802 38724 34814
rect 38668 34750 38670 34802
rect 38722 34750 38724 34802
rect 38668 34468 38724 34750
rect 39452 34692 39508 34702
rect 39564 34692 39620 35646
rect 39788 35140 39844 38780
rect 40012 38770 40068 38780
rect 39340 34690 39620 34692
rect 39340 34638 39454 34690
rect 39506 34638 39620 34690
rect 39340 34636 39620 34638
rect 39676 35138 39844 35140
rect 39676 35086 39790 35138
rect 39842 35086 39844 35138
rect 39676 35084 39844 35086
rect 38668 34402 38724 34412
rect 39228 34468 39284 34478
rect 39340 34468 39396 34636
rect 39452 34626 39508 34636
rect 39284 34412 39396 34468
rect 39228 34402 39284 34412
rect 39452 34356 39508 34366
rect 39340 34244 39396 34254
rect 38332 33842 38388 33852
rect 38668 34132 38724 34142
rect 38444 33348 38500 33358
rect 38164 33346 38500 33348
rect 38164 33294 38446 33346
rect 38498 33294 38500 33346
rect 38164 33292 38500 33294
rect 38108 33254 38164 33292
rect 38444 33282 38500 33292
rect 37884 32498 37940 32508
rect 37996 33234 38052 33246
rect 37996 33182 37998 33234
rect 38050 33182 38052 33234
rect 37996 32786 38052 33182
rect 38668 33234 38724 34076
rect 38668 33182 38670 33234
rect 38722 33182 38724 33234
rect 38668 33170 38724 33182
rect 38780 33236 38836 33246
rect 38780 33142 38836 33180
rect 39340 33012 39396 34188
rect 37996 32734 37998 32786
rect 38050 32734 38052 32786
rect 37436 32284 37604 32340
rect 37268 31836 37380 31892
rect 37212 31826 37268 31836
rect 37324 31666 37380 31836
rect 37324 31614 37326 31666
rect 37378 31614 37380 31666
rect 37324 31602 37380 31614
rect 37436 31666 37492 32284
rect 37772 31892 37828 31902
rect 37436 31614 37438 31666
rect 37490 31614 37492 31666
rect 37436 31602 37492 31614
rect 37548 31890 37828 31892
rect 37548 31838 37774 31890
rect 37826 31838 37828 31890
rect 37548 31836 37828 31838
rect 37212 31556 37268 31566
rect 37100 31554 37268 31556
rect 37100 31502 37214 31554
rect 37266 31502 37268 31554
rect 37100 31500 37268 31502
rect 36988 30210 37044 30828
rect 36988 30158 36990 30210
rect 37042 30158 37044 30210
rect 36988 30146 37044 30158
rect 37212 30210 37268 31500
rect 37212 30158 37214 30210
rect 37266 30158 37268 30210
rect 37212 30146 37268 30158
rect 37436 30660 37492 30670
rect 36540 30034 36596 30044
rect 37100 30100 37156 30110
rect 37100 30006 37156 30044
rect 35756 29362 35812 29372
rect 33180 29314 33236 29326
rect 33180 29262 33182 29314
rect 33234 29262 33236 29314
rect 33068 28756 33124 28766
rect 33180 28756 33236 29262
rect 33964 29316 34020 29326
rect 34300 29316 34356 29326
rect 33964 29314 34300 29316
rect 33964 29262 33966 29314
rect 34018 29262 34300 29314
rect 33964 29260 34300 29262
rect 37436 29316 37492 30604
rect 37548 30210 37604 31836
rect 37772 31826 37828 31836
rect 37996 31892 38052 32734
rect 38780 32956 39396 33012
rect 38780 32674 38836 32956
rect 39004 32732 39284 32788
rect 38780 32622 38782 32674
rect 38834 32622 38836 32674
rect 38780 32610 38836 32622
rect 38892 32674 38948 32686
rect 38892 32622 38894 32674
rect 38946 32622 38948 32674
rect 38892 32564 38948 32622
rect 38892 32498 38948 32508
rect 39004 31948 39060 32732
rect 38668 31892 38724 31902
rect 38052 31836 38276 31892
rect 37996 31826 38052 31836
rect 37548 30158 37550 30210
rect 37602 30158 37604 30210
rect 37548 30146 37604 30158
rect 37996 30210 38052 30222
rect 37996 30158 37998 30210
rect 38050 30158 38052 30210
rect 37996 29988 38052 30158
rect 38220 30098 38276 31836
rect 38668 31666 38724 31836
rect 38668 31614 38670 31666
rect 38722 31614 38724 31666
rect 38668 31602 38724 31614
rect 38780 31892 39060 31948
rect 39116 32562 39172 32574
rect 39116 32510 39118 32562
rect 39170 32510 39172 32562
rect 39116 31948 39172 32510
rect 39228 32564 39284 32732
rect 39452 32676 39508 34300
rect 39676 34356 39732 35084
rect 39788 35074 39844 35084
rect 40012 38612 40068 38622
rect 40012 35922 40068 38556
rect 40124 38052 40180 40684
rect 40236 40516 40292 40526
rect 40236 40422 40292 40460
rect 40348 40514 40404 42028
rect 41804 42084 41860 42094
rect 40908 41300 40964 41310
rect 40348 40462 40350 40514
rect 40402 40462 40404 40514
rect 40348 40450 40404 40462
rect 40796 41298 40964 41300
rect 40796 41246 40910 41298
rect 40962 41246 40964 41298
rect 40796 41244 40964 41246
rect 40796 40516 40852 41244
rect 40908 41234 40964 41244
rect 41244 41186 41300 41198
rect 41244 41134 41246 41186
rect 41298 41134 41300 41186
rect 40796 40450 40852 40460
rect 40908 40740 40964 40750
rect 40908 40402 40964 40684
rect 40908 40350 40910 40402
rect 40962 40350 40964 40402
rect 40908 40338 40964 40350
rect 40236 40180 40292 40190
rect 40236 40086 40292 40124
rect 40460 39730 40516 39742
rect 40460 39678 40462 39730
rect 40514 39678 40516 39730
rect 40460 39060 40516 39678
rect 40460 38994 40516 39004
rect 40572 39732 40628 39742
rect 40180 37996 40404 38052
rect 40124 37958 40180 37996
rect 40236 37828 40292 37838
rect 40236 37734 40292 37772
rect 40348 37156 40404 37996
rect 40572 38050 40628 39676
rect 41132 39730 41188 39742
rect 41132 39678 41134 39730
rect 41186 39678 41188 39730
rect 41132 39396 41188 39678
rect 40572 37998 40574 38050
rect 40626 37998 40628 38050
rect 40572 37986 40628 37998
rect 40684 39340 41188 39396
rect 41244 39620 41300 41134
rect 41692 40292 41748 40302
rect 41580 40290 41748 40292
rect 41580 40238 41694 40290
rect 41746 40238 41748 40290
rect 41580 40236 41748 40238
rect 40460 37940 40516 37950
rect 40460 37846 40516 37884
rect 40684 37828 40740 39340
rect 41020 39172 41076 39182
rect 41076 39116 41188 39172
rect 41020 39106 41076 39116
rect 40796 38948 40852 38958
rect 40796 37938 40852 38892
rect 41020 38834 41076 38846
rect 41020 38782 41022 38834
rect 41074 38782 41076 38834
rect 40908 38052 40964 38062
rect 40908 37958 40964 37996
rect 40796 37886 40798 37938
rect 40850 37886 40852 37938
rect 40796 37874 40852 37886
rect 40684 37762 40740 37772
rect 41020 37604 41076 38782
rect 41132 38052 41188 39116
rect 41244 39058 41300 39564
rect 41244 39006 41246 39058
rect 41298 39006 41300 39058
rect 41244 38994 41300 39006
rect 41356 40180 41412 40190
rect 41244 38052 41300 38062
rect 41132 38050 41300 38052
rect 41132 37998 41246 38050
rect 41298 37998 41300 38050
rect 41132 37996 41300 37998
rect 41244 37986 41300 37996
rect 41356 37938 41412 40124
rect 41580 38050 41636 40236
rect 41692 40226 41748 40236
rect 41580 37998 41582 38050
rect 41634 37998 41636 38050
rect 41580 37986 41636 37998
rect 41804 38052 41860 42028
rect 41916 41858 41972 43036
rect 43596 42084 43652 42094
rect 43596 41990 43652 42028
rect 43708 42084 43764 42094
rect 43708 42082 43876 42084
rect 43708 42030 43710 42082
rect 43762 42030 43876 42082
rect 43708 42028 43876 42030
rect 43708 42018 43764 42028
rect 43036 41972 43092 41982
rect 43036 41878 43092 41916
rect 41916 41806 41918 41858
rect 41970 41806 41972 41858
rect 41916 41794 41972 41806
rect 43708 41746 43764 41758
rect 43708 41694 43710 41746
rect 43762 41694 43764 41746
rect 42028 41076 42084 41086
rect 42028 40982 42084 41020
rect 41916 40180 41972 40190
rect 41916 38948 41972 40124
rect 43148 39732 43204 39742
rect 43148 39058 43204 39676
rect 43148 39006 43150 39058
rect 43202 39006 43204 39058
rect 43148 38994 43204 39006
rect 43260 39506 43316 39518
rect 43260 39454 43262 39506
rect 43314 39454 43316 39506
rect 41916 38882 41972 38892
rect 43148 38276 43204 38286
rect 43260 38276 43316 39454
rect 43708 39060 43764 41694
rect 43820 41300 43876 42028
rect 44492 41972 44548 41982
rect 44156 41300 44212 41310
rect 43820 41298 44212 41300
rect 43820 41246 44158 41298
rect 44210 41246 44212 41298
rect 43820 41244 44212 41246
rect 44044 40628 44100 40638
rect 43148 38274 43316 38276
rect 43148 38222 43150 38274
rect 43202 38222 43316 38274
rect 43148 38220 43316 38222
rect 43372 39004 43764 39060
rect 43820 40292 43876 40302
rect 43148 38210 43204 38220
rect 41356 37886 41358 37938
rect 41410 37886 41412 37938
rect 41356 37874 41412 37886
rect 41804 37938 41860 37996
rect 42700 38052 42756 38062
rect 43372 38052 43428 39004
rect 41804 37886 41806 37938
rect 41858 37886 41860 37938
rect 41804 37874 41860 37886
rect 42476 37938 42532 37950
rect 42476 37886 42478 37938
rect 42530 37886 42532 37938
rect 42140 37828 42196 37838
rect 42476 37828 42532 37886
rect 42140 37826 42532 37828
rect 42140 37774 42142 37826
rect 42194 37774 42532 37826
rect 42140 37772 42532 37774
rect 42140 37762 42196 37772
rect 41020 37548 41300 37604
rect 41132 37378 41188 37390
rect 41132 37326 41134 37378
rect 41186 37326 41188 37378
rect 40796 37268 40852 37278
rect 41020 37268 41076 37278
rect 40348 37100 40516 37156
rect 40012 35870 40014 35922
rect 40066 35870 40068 35922
rect 40012 35140 40068 35870
rect 40236 35700 40292 35710
rect 40012 35074 40068 35084
rect 40124 35698 40292 35700
rect 40124 35646 40238 35698
rect 40290 35646 40292 35698
rect 40124 35644 40292 35646
rect 40012 34916 40068 34926
rect 39900 34914 40068 34916
rect 39900 34862 40014 34914
rect 40066 34862 40068 34914
rect 39900 34860 40068 34862
rect 39676 34354 39844 34356
rect 39676 34302 39678 34354
rect 39730 34302 39844 34354
rect 39676 34300 39844 34302
rect 39676 34290 39732 34300
rect 39676 33236 39732 33246
rect 39452 32610 39508 32620
rect 39564 33122 39620 33134
rect 39564 33070 39566 33122
rect 39618 33070 39620 33122
rect 39340 32564 39396 32574
rect 39228 32562 39396 32564
rect 39228 32510 39342 32562
rect 39394 32510 39396 32562
rect 39228 32508 39396 32510
rect 39340 32498 39396 32508
rect 39564 32004 39620 33070
rect 39676 32786 39732 33180
rect 39676 32734 39678 32786
rect 39730 32734 39732 32786
rect 39676 32722 39732 32734
rect 39116 31892 39508 31948
rect 38780 31666 38836 31892
rect 38780 31614 38782 31666
rect 38834 31614 38836 31666
rect 38444 31556 38500 31566
rect 38444 31462 38500 31500
rect 38780 31220 38836 31614
rect 39116 31778 39172 31790
rect 39340 31780 39396 31790
rect 39116 31726 39118 31778
rect 39170 31726 39172 31778
rect 38892 31220 38948 31230
rect 38780 31218 38948 31220
rect 38780 31166 38894 31218
rect 38946 31166 38948 31218
rect 38780 31164 38948 31166
rect 38892 31154 38948 31164
rect 39116 31106 39172 31726
rect 39116 31054 39118 31106
rect 39170 31054 39172 31106
rect 38668 30884 38724 30894
rect 38668 30790 38724 30828
rect 38220 30046 38222 30098
rect 38274 30046 38276 30098
rect 38220 30034 38276 30046
rect 39116 30100 39172 31054
rect 39228 31778 39396 31780
rect 39228 31726 39342 31778
rect 39394 31726 39396 31778
rect 39228 31724 39396 31726
rect 39228 30996 39284 31724
rect 39340 31714 39396 31724
rect 39228 30902 39284 30940
rect 39340 31108 39396 31118
rect 39340 30322 39396 31052
rect 39340 30270 39342 30322
rect 39394 30270 39396 30322
rect 39340 30258 39396 30270
rect 39452 30324 39508 31892
rect 39564 31780 39620 31948
rect 39676 32004 39732 32014
rect 39788 32004 39844 34300
rect 39900 34244 39956 34860
rect 40012 34850 40068 34860
rect 39900 33346 39956 34188
rect 40012 34692 40068 34702
rect 40012 34242 40068 34636
rect 40012 34190 40014 34242
rect 40066 34190 40068 34242
rect 40012 34178 40068 34190
rect 39900 33294 39902 33346
rect 39954 33294 39956 33346
rect 39900 33282 39956 33294
rect 40124 32900 40180 35644
rect 40236 35634 40292 35644
rect 40348 35364 40404 35374
rect 40348 34354 40404 35308
rect 40460 34916 40516 37100
rect 40796 36594 40852 37212
rect 40796 36542 40798 36594
rect 40850 36542 40852 36594
rect 40796 36530 40852 36542
rect 40908 37266 41076 37268
rect 40908 37214 41022 37266
rect 41074 37214 41076 37266
rect 40908 37212 41076 37214
rect 40908 35812 40964 37212
rect 41020 37202 41076 37212
rect 40460 34802 40516 34860
rect 40460 34750 40462 34802
rect 40514 34750 40516 34802
rect 40460 34738 40516 34750
rect 40796 35756 40964 35812
rect 41132 36594 41188 37326
rect 41132 36542 41134 36594
rect 41186 36542 41188 36594
rect 40796 34914 40852 35756
rect 41132 35700 41188 36542
rect 41132 35634 41188 35644
rect 40796 34862 40798 34914
rect 40850 34862 40852 34914
rect 40348 34302 40350 34354
rect 40402 34302 40404 34354
rect 40348 34290 40404 34302
rect 40348 34132 40404 34142
rect 39676 32002 39844 32004
rect 39676 31950 39678 32002
rect 39730 31950 39844 32002
rect 39676 31948 39844 31950
rect 39900 32844 40180 32900
rect 39676 31938 39732 31948
rect 39564 31714 39620 31724
rect 39900 31556 39956 32844
rect 40124 32788 40180 32844
rect 40124 32722 40180 32732
rect 40236 33348 40292 33358
rect 40348 33348 40404 34076
rect 40796 33572 40852 34862
rect 40908 35586 40964 35598
rect 40908 35534 40910 35586
rect 40962 35534 40964 35586
rect 40908 34244 40964 35534
rect 41244 35364 41300 37548
rect 41356 37266 41412 37278
rect 41356 37214 41358 37266
rect 41410 37214 41412 37266
rect 41356 35588 41412 37214
rect 41580 37268 41636 37278
rect 41580 37174 41636 37212
rect 41356 35522 41412 35532
rect 41244 34914 41300 35308
rect 41916 35026 41972 35038
rect 41916 34974 41918 35026
rect 41970 34974 41972 35026
rect 41244 34862 41246 34914
rect 41298 34862 41300 34914
rect 41244 34850 41300 34862
rect 41804 34916 41860 34926
rect 41916 34916 41972 34974
rect 41860 34860 41972 34916
rect 41804 34850 41860 34860
rect 41804 34356 41860 34366
rect 41804 34262 41860 34300
rect 40908 34150 40964 34188
rect 41244 34244 41300 34254
rect 41244 34150 41300 34188
rect 42140 34132 42196 34142
rect 42140 34038 42196 34076
rect 42476 34018 42532 37772
rect 42588 37828 42644 37838
rect 42588 37734 42644 37772
rect 42700 35924 42756 37996
rect 43148 37996 43428 38052
rect 43596 38052 43652 38062
rect 43036 37940 43092 37950
rect 43036 37846 43092 37884
rect 43148 37938 43204 37996
rect 43596 37958 43652 37996
rect 43148 37886 43150 37938
rect 43202 37886 43204 37938
rect 43148 37874 43204 37886
rect 43708 37940 43764 37950
rect 43820 37940 43876 40236
rect 43932 39620 43988 39630
rect 43932 39526 43988 39564
rect 43932 38052 43988 38062
rect 44044 38052 44100 40572
rect 44156 40180 44212 41244
rect 44156 40114 44212 40124
rect 43932 38050 44100 38052
rect 43932 37998 43934 38050
rect 43986 37998 44100 38050
rect 43932 37996 44100 37998
rect 44156 38834 44212 38846
rect 44156 38782 44158 38834
rect 44210 38782 44212 38834
rect 43932 37986 43988 37996
rect 43708 37938 43876 37940
rect 43708 37886 43710 37938
rect 43762 37886 43876 37938
rect 43708 37884 43876 37886
rect 43708 37874 43764 37884
rect 42812 37828 42868 37838
rect 42812 37826 42980 37828
rect 42812 37774 42814 37826
rect 42866 37774 42980 37826
rect 42812 37772 42980 37774
rect 42812 37762 42868 37772
rect 42924 36036 42980 37772
rect 43484 37044 43540 37054
rect 43484 36950 43540 36988
rect 43932 36484 43988 36494
rect 43820 36482 43988 36484
rect 43820 36430 43934 36482
rect 43986 36430 43988 36482
rect 43820 36428 43988 36430
rect 43260 36372 43316 36382
rect 43260 36370 43540 36372
rect 43260 36318 43262 36370
rect 43314 36318 43540 36370
rect 43260 36316 43540 36318
rect 43260 36306 43316 36316
rect 42924 35980 43316 36036
rect 42700 35868 43092 35924
rect 43036 35810 43092 35868
rect 43036 35758 43038 35810
rect 43090 35758 43092 35810
rect 43036 35746 43092 35758
rect 43148 35588 43204 35598
rect 42588 34244 42644 34254
rect 42588 34150 42644 34188
rect 43148 34242 43204 35532
rect 43260 34354 43316 35980
rect 43260 34302 43262 34354
rect 43314 34302 43316 34354
rect 43260 34290 43316 34302
rect 43484 34354 43540 36316
rect 43820 35700 43876 36428
rect 43932 36418 43988 36428
rect 44156 36372 44212 38782
rect 44156 36316 44436 36372
rect 43820 35606 43876 35644
rect 43932 36260 43988 36270
rect 43484 34302 43486 34354
rect 43538 34302 43540 34354
rect 43484 34290 43540 34302
rect 43148 34190 43150 34242
rect 43202 34190 43204 34242
rect 43148 34178 43204 34190
rect 42476 33966 42478 34018
rect 42530 33966 42532 34018
rect 42476 33954 42532 33966
rect 43820 34020 43876 34030
rect 43820 33926 43876 33964
rect 42812 33908 42868 33918
rect 42812 33906 42980 33908
rect 42812 33854 42814 33906
rect 42866 33854 42980 33906
rect 42812 33852 42980 33854
rect 42812 33842 42868 33852
rect 41020 33572 41076 33582
rect 40796 33570 41076 33572
rect 40796 33518 41022 33570
rect 41074 33518 41076 33570
rect 40796 33516 41076 33518
rect 41020 33506 41076 33516
rect 40236 33346 40404 33348
rect 40236 33294 40238 33346
rect 40290 33294 40404 33346
rect 40236 33292 40404 33294
rect 40012 32676 40068 32686
rect 40012 32582 40068 32620
rect 40236 32564 40292 33292
rect 40460 33234 40516 33246
rect 40460 33182 40462 33234
rect 40514 33182 40516 33234
rect 40348 32788 40404 32798
rect 40348 32694 40404 32732
rect 40124 32508 40292 32564
rect 39564 31500 39956 31556
rect 40012 31666 40068 31678
rect 40012 31614 40014 31666
rect 40066 31614 40068 31666
rect 39564 30660 39620 31500
rect 40012 31444 40068 31614
rect 39900 31388 40068 31444
rect 39676 31332 39732 31342
rect 39900 31332 39956 31388
rect 39676 31106 39732 31276
rect 39676 31054 39678 31106
rect 39730 31054 39732 31106
rect 39676 31042 39732 31054
rect 39788 31276 39956 31332
rect 40124 31332 40180 32508
rect 40236 32340 40292 32350
rect 40236 31554 40292 32284
rect 40460 32116 40516 33182
rect 40572 33236 40628 33246
rect 40572 33142 40628 33180
rect 41356 32788 41412 32798
rect 41020 32564 41076 32574
rect 40460 32050 40516 32060
rect 40572 32508 41020 32564
rect 40572 31892 40628 32508
rect 41020 32470 41076 32508
rect 41356 32562 41412 32732
rect 42924 32788 42980 33852
rect 43148 33124 43204 33134
rect 43148 33030 43204 33068
rect 42924 32694 42980 32732
rect 43372 32674 43428 32686
rect 43372 32622 43374 32674
rect 43426 32622 43428 32674
rect 41356 32510 41358 32562
rect 41410 32510 41412 32562
rect 41132 32340 41188 32350
rect 41132 32246 41188 32284
rect 41356 31948 41412 32510
rect 41804 32562 41860 32574
rect 41804 32510 41806 32562
rect 41858 32510 41860 32562
rect 40460 31836 40628 31892
rect 41020 31892 41412 31948
rect 41468 32338 41524 32350
rect 41468 32286 41470 32338
rect 41522 32286 41524 32338
rect 41468 31948 41524 32286
rect 41468 31892 41748 31948
rect 40348 31780 40404 31790
rect 40348 31686 40404 31724
rect 40236 31502 40238 31554
rect 40290 31502 40292 31554
rect 40236 31490 40292 31502
rect 39788 30994 39844 31276
rect 40124 31266 40180 31276
rect 40348 31220 40404 31230
rect 40460 31220 40516 31836
rect 40348 31218 40516 31220
rect 40348 31166 40350 31218
rect 40402 31166 40516 31218
rect 40348 31164 40516 31166
rect 40572 31666 40628 31678
rect 40572 31614 40574 31666
rect 40626 31614 40628 31666
rect 40348 31154 40404 31164
rect 39900 31108 39956 31118
rect 39900 31014 39956 31052
rect 40572 31108 40628 31614
rect 41020 31556 41076 31892
rect 41244 31666 41300 31678
rect 41244 31614 41246 31666
rect 41298 31614 41300 31666
rect 41020 31462 41076 31500
rect 41132 31554 41188 31566
rect 41132 31502 41134 31554
rect 41186 31502 41188 31554
rect 40572 31042 40628 31052
rect 39788 30942 39790 30994
rect 39842 30942 39844 30994
rect 39788 30884 39844 30942
rect 41020 30996 41076 31006
rect 39788 30818 39844 30828
rect 40908 30884 40964 30894
rect 40908 30790 40964 30828
rect 39564 30604 40292 30660
rect 39452 30258 39508 30268
rect 39116 30034 39172 30044
rect 37548 29316 37604 29326
rect 37436 29314 37604 29316
rect 37436 29262 37550 29314
rect 37602 29262 37604 29314
rect 37436 29260 37604 29262
rect 33964 29250 34020 29260
rect 34300 29222 34356 29260
rect 37548 29250 37604 29260
rect 37996 29316 38052 29932
rect 37996 29250 38052 29260
rect 38780 29988 38836 29998
rect 33068 28754 33236 28756
rect 33068 28702 33070 28754
rect 33122 28702 33236 28754
rect 33068 28700 33236 28702
rect 34748 29204 34804 29214
rect 33068 28690 33124 28700
rect 33740 28644 33796 28654
rect 33740 28550 33796 28588
rect 34300 28644 34356 28654
rect 34300 28550 34356 28588
rect 34748 26964 34804 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 38780 27748 38836 29932
rect 40012 29538 40068 29550
rect 40012 29486 40014 29538
rect 40066 29486 40068 29538
rect 40012 29428 40068 29486
rect 40012 29362 40068 29372
rect 40236 29426 40292 30604
rect 40236 29374 40238 29426
rect 40290 29374 40292 29426
rect 40236 29362 40292 29374
rect 40908 29428 40964 29438
rect 40908 29334 40964 29372
rect 41020 28644 41076 30940
rect 41132 29988 41188 31502
rect 41244 30212 41300 31614
rect 41244 30146 41300 30156
rect 41468 30212 41524 30222
rect 41692 30212 41748 31892
rect 41804 30884 41860 32510
rect 41804 30818 41860 30828
rect 42028 32562 42084 32574
rect 42028 32510 42030 32562
rect 42082 32510 42084 32562
rect 41468 30210 41748 30212
rect 41468 30158 41470 30210
rect 41522 30158 41748 30210
rect 41468 30156 41748 30158
rect 41916 30324 41972 30334
rect 41468 30146 41524 30156
rect 41132 29932 41748 29988
rect 41692 29538 41748 29932
rect 41692 29486 41694 29538
rect 41746 29486 41748 29538
rect 41692 29474 41748 29486
rect 41916 28754 41972 30268
rect 42028 30100 42084 32510
rect 42476 32564 42532 32574
rect 42532 32508 42868 32564
rect 42476 32470 42532 32508
rect 42252 32450 42308 32462
rect 42252 32398 42254 32450
rect 42306 32398 42308 32450
rect 42252 32340 42308 32398
rect 42700 32340 42756 32350
rect 42252 32338 42756 32340
rect 42252 32286 42702 32338
rect 42754 32286 42756 32338
rect 42252 32284 42756 32286
rect 42700 32274 42756 32284
rect 42028 30034 42084 30044
rect 42140 30210 42196 30222
rect 42140 30158 42142 30210
rect 42194 30158 42196 30210
rect 42140 29428 42196 30158
rect 42588 30212 42644 30222
rect 42588 30118 42644 30156
rect 42812 30210 42868 32508
rect 43036 32338 43092 32350
rect 43036 32286 43038 32338
rect 43090 32286 43092 32338
rect 43036 31106 43092 32286
rect 43036 31054 43038 31106
rect 43090 31054 43092 31106
rect 43036 31042 43092 31054
rect 43148 31554 43204 31566
rect 43148 31502 43150 31554
rect 43202 31502 43204 31554
rect 43148 30436 43204 31502
rect 43372 30996 43428 32622
rect 43596 32676 43652 32686
rect 43596 32562 43652 32620
rect 43596 32510 43598 32562
rect 43650 32510 43652 32562
rect 43596 32498 43652 32510
rect 43708 30996 43764 31006
rect 43372 30940 43708 30996
rect 43708 30902 43764 30940
rect 43148 30370 43204 30380
rect 42812 30158 42814 30210
rect 42866 30158 42868 30210
rect 42812 30146 42868 30158
rect 43484 30210 43540 30222
rect 43484 30158 43486 30210
rect 43538 30158 43540 30210
rect 42140 29362 42196 29372
rect 43484 30100 43540 30158
rect 43484 29316 43540 30044
rect 43820 29316 43876 29326
rect 43484 29314 43876 29316
rect 43484 29262 43822 29314
rect 43874 29262 43876 29314
rect 43484 29260 43876 29262
rect 43820 29250 43876 29260
rect 41916 28702 41918 28754
rect 41970 28702 41972 28754
rect 41916 28690 41972 28702
rect 41244 28644 41300 28654
rect 41020 28642 41300 28644
rect 41020 28590 41246 28642
rect 41298 28590 41300 28642
rect 41020 28588 41300 28590
rect 41244 28578 41300 28588
rect 43820 27970 43876 27982
rect 43820 27918 43822 27970
rect 43874 27918 43876 27970
rect 41804 27748 41860 27758
rect 38780 27692 39060 27748
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35084 27188 35140 27198
rect 35084 27094 35140 27132
rect 37100 27188 37156 27198
rect 37156 27132 37492 27188
rect 37100 27094 37156 27132
rect 34748 26870 34804 26908
rect 35644 26964 35700 26974
rect 35644 26870 35700 26908
rect 36092 26962 36148 26974
rect 36092 26910 36094 26962
rect 36146 26910 36148 26962
rect 35980 26850 36036 26862
rect 35980 26798 35982 26850
rect 36034 26798 36036 26850
rect 34188 26516 34244 26526
rect 34188 26514 35028 26516
rect 34188 26462 34190 26514
rect 34242 26462 35028 26514
rect 34188 26460 35028 26462
rect 34188 26450 34244 26460
rect 34636 26290 34692 26302
rect 34636 26238 34638 26290
rect 34690 26238 34692 26290
rect 34076 26180 34132 26190
rect 33068 25506 33124 25518
rect 33068 25454 33070 25506
rect 33122 25454 33124 25506
rect 33068 24724 33124 25454
rect 33068 24658 33124 24668
rect 33516 25506 33572 25518
rect 33516 25454 33518 25506
rect 33570 25454 33572 25506
rect 32956 24052 33012 24062
rect 33292 24052 33348 24062
rect 32956 24050 33348 24052
rect 32956 23998 32958 24050
rect 33010 23998 33294 24050
rect 33346 23998 33348 24050
rect 32956 23996 33348 23998
rect 32956 23986 33012 23996
rect 33292 23986 33348 23996
rect 33404 23714 33460 23726
rect 33404 23662 33406 23714
rect 33458 23662 33460 23714
rect 33068 23380 33124 23390
rect 33068 22484 33124 23324
rect 33404 23268 33460 23662
rect 33516 23604 33572 25454
rect 34076 24722 34132 26124
rect 34636 25620 34692 26238
rect 34972 26290 35028 26460
rect 34972 26238 34974 26290
rect 35026 26238 35028 26290
rect 34972 26226 35028 26238
rect 34076 24670 34078 24722
rect 34130 24670 34132 24722
rect 34076 24658 34132 24670
rect 34524 25564 34636 25620
rect 33740 24612 33796 24622
rect 33740 24518 33796 24556
rect 34188 23604 34244 23614
rect 33516 23548 34188 23604
rect 33404 23202 33460 23212
rect 33964 23268 34020 23278
rect 33964 22484 34020 23212
rect 33068 22390 33124 22428
rect 33852 22482 34020 22484
rect 33852 22430 33966 22482
rect 34018 22430 34020 22482
rect 33852 22428 34020 22430
rect 33740 22370 33796 22382
rect 33740 22318 33742 22370
rect 33794 22318 33796 22370
rect 33068 20804 33124 20814
rect 32844 20802 33124 20804
rect 32844 20750 33070 20802
rect 33122 20750 33124 20802
rect 32844 20748 33124 20750
rect 33068 20738 33124 20748
rect 33404 20580 33460 20590
rect 33292 20578 33460 20580
rect 33292 20526 33406 20578
rect 33458 20526 33460 20578
rect 33292 20524 33460 20526
rect 33740 20580 33796 22318
rect 33852 20802 33908 22428
rect 33964 22418 34020 22428
rect 34076 22372 34132 22382
rect 33964 21586 34020 21598
rect 33964 21534 33966 21586
rect 34018 21534 34020 21586
rect 33964 20914 34020 21534
rect 34076 21362 34132 22316
rect 34188 22370 34244 23548
rect 34188 22318 34190 22370
rect 34242 22318 34244 22370
rect 34188 22306 34244 22318
rect 34412 22708 34468 22718
rect 34412 22260 34468 22652
rect 34524 22484 34580 25564
rect 34636 25554 34692 25564
rect 35084 26180 35140 26190
rect 34972 24724 35028 24734
rect 34636 24612 34692 24622
rect 34636 24610 34916 24612
rect 34636 24558 34638 24610
rect 34690 24558 34916 24610
rect 34636 24556 34916 24558
rect 34636 24546 34692 24556
rect 34524 22418 34580 22428
rect 34860 22372 34916 24556
rect 34972 23938 35028 24668
rect 35084 24722 35140 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35868 25282 35924 25294
rect 35868 25230 35870 25282
rect 35922 25230 35924 25282
rect 35868 24948 35924 25230
rect 35868 24882 35924 24892
rect 35084 24670 35086 24722
rect 35138 24670 35140 24722
rect 35084 24658 35140 24670
rect 35532 24724 35588 24734
rect 35980 24724 36036 26798
rect 35532 24722 36036 24724
rect 35532 24670 35534 24722
rect 35586 24670 36036 24722
rect 35532 24668 36036 24670
rect 36092 24724 36148 26910
rect 35532 24658 35588 24668
rect 36092 24658 36148 24668
rect 36204 26964 36260 26974
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34972 23886 34974 23938
rect 35026 23886 35028 23938
rect 34972 23268 35028 23886
rect 35196 23940 35252 23950
rect 35084 23268 35140 23278
rect 34972 23266 35140 23268
rect 34972 23214 35086 23266
rect 35138 23214 35140 23266
rect 34972 23212 35140 23214
rect 35196 23268 35252 23884
rect 35420 23940 35476 23950
rect 36204 23940 36260 26908
rect 37436 25506 37492 27132
rect 38556 26962 38612 26974
rect 38556 26910 38558 26962
rect 38610 26910 38612 26962
rect 38220 26852 38276 26862
rect 37548 26850 38276 26852
rect 37548 26798 38222 26850
rect 38274 26798 38276 26850
rect 37548 26796 38276 26798
rect 37548 26514 37604 26796
rect 38220 26786 38276 26796
rect 37548 26462 37550 26514
rect 37602 26462 37604 26514
rect 37548 26450 37604 26462
rect 37996 26404 38052 26414
rect 37884 26180 37940 26190
rect 37884 26086 37940 26124
rect 37436 25454 37438 25506
rect 37490 25454 37492 25506
rect 37436 25442 37492 25454
rect 37548 25730 37604 25742
rect 37548 25678 37550 25730
rect 37602 25678 37604 25730
rect 35420 23938 35700 23940
rect 35420 23886 35422 23938
rect 35474 23886 35700 23938
rect 35420 23884 35700 23886
rect 35420 23874 35476 23884
rect 35308 23714 35364 23726
rect 35308 23662 35310 23714
rect 35362 23662 35364 23714
rect 35308 23380 35364 23662
rect 35532 23716 35588 23726
rect 35532 23622 35588 23660
rect 35532 23380 35588 23390
rect 35308 23378 35588 23380
rect 35308 23326 35534 23378
rect 35586 23326 35588 23378
rect 35308 23324 35588 23326
rect 35532 23314 35588 23324
rect 35196 23212 35364 23268
rect 35084 23202 35140 23212
rect 35308 23154 35364 23212
rect 35308 23102 35310 23154
rect 35362 23102 35364 23154
rect 35308 23090 35364 23102
rect 34972 23042 35028 23054
rect 34972 22990 34974 23042
rect 35026 22990 35028 23042
rect 34972 22594 35028 22990
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34972 22542 34974 22594
rect 35026 22542 35028 22594
rect 34972 22530 35028 22542
rect 35644 22596 35700 23884
rect 35644 22530 35700 22540
rect 35756 23884 36260 23940
rect 36540 25282 36596 25294
rect 36540 25230 36542 25282
rect 36594 25230 36596 25282
rect 35196 22372 35252 22382
rect 34860 22370 35252 22372
rect 34860 22318 35198 22370
rect 35250 22318 35252 22370
rect 34860 22316 35252 22318
rect 35196 22306 35252 22316
rect 35420 22372 35476 22382
rect 35420 22278 35476 22316
rect 35644 22372 35700 22382
rect 35644 22278 35700 22316
rect 34412 22166 34468 22204
rect 34300 22146 34356 22158
rect 34300 22094 34302 22146
rect 34354 22094 34356 22146
rect 34300 22036 34356 22094
rect 35084 22146 35140 22158
rect 35084 22094 35086 22146
rect 35138 22094 35140 22146
rect 35084 22036 35140 22094
rect 34300 21980 34692 22036
rect 34188 21924 34244 21934
rect 34636 21924 34692 21980
rect 35084 21970 35140 21980
rect 35196 22148 35252 22158
rect 34636 21868 35028 21924
rect 34188 21812 34244 21868
rect 34188 21756 34468 21812
rect 34412 21698 34468 21756
rect 34412 21646 34414 21698
rect 34466 21646 34468 21698
rect 34412 21634 34468 21646
rect 34748 21700 34804 21710
rect 34076 21310 34078 21362
rect 34130 21310 34132 21362
rect 34076 21298 34132 21310
rect 34188 21586 34244 21598
rect 34188 21534 34190 21586
rect 34242 21534 34244 21586
rect 33964 20862 33966 20914
rect 34018 20862 34020 20914
rect 33964 20850 34020 20862
rect 34188 20916 34244 21534
rect 34636 21588 34692 21598
rect 34748 21588 34804 21644
rect 34972 21698 35028 21868
rect 34972 21646 34974 21698
rect 35026 21646 35028 21698
rect 34972 21634 35028 21646
rect 35196 21700 35252 22092
rect 35644 21700 35700 21710
rect 35196 21634 35252 21644
rect 35420 21644 35644 21700
rect 34636 21586 34804 21588
rect 34636 21534 34638 21586
rect 34690 21534 34804 21586
rect 34636 21532 34804 21534
rect 35420 21586 35476 21644
rect 35644 21634 35700 21644
rect 35420 21534 35422 21586
rect 35474 21534 35476 21586
rect 34636 21522 34692 21532
rect 35420 21522 35476 21534
rect 35196 21364 35252 21374
rect 35644 21364 35700 21374
rect 35084 21362 35252 21364
rect 35084 21310 35198 21362
rect 35250 21310 35252 21362
rect 35084 21308 35252 21310
rect 34188 20850 34244 20860
rect 34300 21028 34356 21038
rect 35084 21028 35140 21308
rect 35196 21298 35252 21308
rect 35532 21362 35700 21364
rect 35532 21310 35646 21362
rect 35698 21310 35700 21362
rect 35532 21308 35700 21310
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 20972 35252 21028
rect 33852 20750 33854 20802
rect 33906 20750 33908 20802
rect 33852 20738 33908 20750
rect 34188 20692 34244 20702
rect 34188 20598 34244 20636
rect 33964 20580 34020 20590
rect 33740 20578 34020 20580
rect 33740 20526 33966 20578
rect 34018 20526 34020 20578
rect 33740 20524 34020 20526
rect 33068 20132 33124 20142
rect 32956 20130 33124 20132
rect 32956 20078 33070 20130
rect 33122 20078 33124 20130
rect 32956 20076 33124 20078
rect 32844 20020 32900 20030
rect 32844 19458 32900 19964
rect 32844 19406 32846 19458
rect 32898 19406 32900 19458
rect 32844 19394 32900 19406
rect 32844 19236 32900 19246
rect 32956 19236 33012 20076
rect 33068 20066 33124 20076
rect 32844 19234 33012 19236
rect 32844 19182 32846 19234
rect 32898 19182 33012 19234
rect 32844 19180 33012 19182
rect 32844 19170 32900 19180
rect 32620 18162 32676 18172
rect 32284 17668 32340 17678
rect 32284 17666 32676 17668
rect 32284 17614 32286 17666
rect 32338 17614 32676 17666
rect 32284 17612 32676 17614
rect 32284 17602 32340 17612
rect 32508 17444 32564 17454
rect 32620 17444 32676 17612
rect 32844 17444 32900 17454
rect 32620 17442 32900 17444
rect 32620 17390 32846 17442
rect 32898 17390 32900 17442
rect 32620 17388 32900 17390
rect 32508 17350 32564 17388
rect 31948 16324 32004 16334
rect 31948 16098 32004 16268
rect 32508 16100 32564 16110
rect 31948 16046 31950 16098
rect 32002 16046 32004 16098
rect 31948 16034 32004 16046
rect 32396 16098 32564 16100
rect 32396 16046 32510 16098
rect 32562 16046 32564 16098
rect 32396 16044 32564 16046
rect 32284 15876 32340 15886
rect 32060 15874 32340 15876
rect 32060 15822 32286 15874
rect 32338 15822 32340 15874
rect 32060 15820 32340 15822
rect 32060 15540 32116 15820
rect 32284 15810 32340 15820
rect 30828 13970 31108 13972
rect 30828 13918 30830 13970
rect 30882 13918 31108 13970
rect 30828 13916 31108 13918
rect 30828 13906 30884 13916
rect 31052 13076 31108 13916
rect 31276 13906 31332 13916
rect 31388 15092 31556 15148
rect 31724 15092 31892 15148
rect 31948 15484 32116 15540
rect 32396 15538 32452 16044
rect 32508 16034 32564 16044
rect 32396 15486 32398 15538
rect 32450 15486 32452 15538
rect 31276 13748 31332 13758
rect 31276 13654 31332 13692
rect 31164 13076 31220 13086
rect 31052 13074 31220 13076
rect 31052 13022 31166 13074
rect 31218 13022 31220 13074
rect 31052 13020 31220 13022
rect 31164 13010 31220 13020
rect 30604 12402 30772 12404
rect 30604 12350 30606 12402
rect 30658 12350 30772 12402
rect 30604 12348 30772 12350
rect 30604 12338 30660 12348
rect 30940 12292 30996 12302
rect 30940 12198 30996 12236
rect 31388 12068 31444 15092
rect 31500 13860 31556 13870
rect 31500 12740 31556 13804
rect 31724 13748 31780 15092
rect 31948 14642 32004 15484
rect 32396 15474 32452 15486
rect 32060 15092 32116 15102
rect 32060 14998 32116 15036
rect 31948 14590 31950 14642
rect 32002 14590 32004 14642
rect 31948 14578 32004 14590
rect 31836 13972 31892 13982
rect 31836 13858 31892 13916
rect 31836 13806 31838 13858
rect 31890 13806 31892 13858
rect 31836 13794 31892 13806
rect 32060 13860 32116 13870
rect 32060 13766 32116 13804
rect 32620 13860 32676 13870
rect 31724 13682 31780 13692
rect 31948 13748 32004 13758
rect 31948 13076 32004 13692
rect 32172 13522 32228 13534
rect 32172 13470 32174 13522
rect 32226 13470 32228 13522
rect 32060 13076 32116 13086
rect 31948 13074 32116 13076
rect 31948 13022 32062 13074
rect 32114 13022 32116 13074
rect 31948 13020 32116 13022
rect 32060 13010 32116 13020
rect 32172 12852 32228 13470
rect 31500 12646 31556 12684
rect 32060 12796 32228 12852
rect 32620 12962 32676 13804
rect 32620 12910 32622 12962
rect 32674 12910 32676 12962
rect 32060 12178 32116 12796
rect 32060 12126 32062 12178
rect 32114 12126 32116 12178
rect 32060 12114 32116 12126
rect 32284 12178 32340 12190
rect 32284 12126 32286 12178
rect 32338 12126 32340 12178
rect 30268 11554 30324 11564
rect 31164 12012 31444 12068
rect 31164 11508 31220 12012
rect 30604 11506 31220 11508
rect 30604 11454 31166 11506
rect 31218 11454 31220 11506
rect 30604 11452 31220 11454
rect 30492 11282 30548 11294
rect 30492 11230 30494 11282
rect 30546 11230 30548 11282
rect 30156 11172 30212 11182
rect 30492 11172 30548 11230
rect 30604 11282 30660 11452
rect 31164 11442 31220 11452
rect 30604 11230 30606 11282
rect 30658 11230 30660 11282
rect 30604 11218 30660 11230
rect 30156 11170 30548 11172
rect 30156 11118 30158 11170
rect 30210 11118 30548 11170
rect 30156 11116 30548 11118
rect 30156 11106 30212 11116
rect 30044 10892 30436 10948
rect 29148 9826 29204 10556
rect 29932 10500 29988 10510
rect 30380 10500 30436 10892
rect 30492 10724 30548 11116
rect 30828 11172 30884 11182
rect 30828 11170 31108 11172
rect 30828 11118 30830 11170
rect 30882 11118 31108 11170
rect 30828 11116 31108 11118
rect 30828 11106 30884 11116
rect 31052 10948 31108 11116
rect 31052 10892 31332 10948
rect 31276 10834 31332 10892
rect 31276 10782 31278 10834
rect 31330 10782 31332 10834
rect 31276 10770 31332 10782
rect 31052 10724 31108 10734
rect 30492 10668 30660 10724
rect 30604 10612 30660 10668
rect 31052 10630 31108 10668
rect 30828 10612 30884 10622
rect 30604 10610 30884 10612
rect 30604 10558 30830 10610
rect 30882 10558 30884 10610
rect 30604 10556 30884 10558
rect 30492 10500 30548 10510
rect 30380 10498 30548 10500
rect 30380 10446 30494 10498
rect 30546 10446 30548 10498
rect 30380 10444 30548 10446
rect 29932 9938 29988 10444
rect 30492 10052 30548 10444
rect 30492 9986 30548 9996
rect 29932 9886 29934 9938
rect 29986 9886 29988 9938
rect 29932 9874 29988 9886
rect 29148 9774 29150 9826
rect 29202 9774 29204 9826
rect 28476 8866 28532 8876
rect 25788 8082 25844 8092
rect 28812 7924 28868 7934
rect 28252 7700 28308 7710
rect 28252 7698 28532 7700
rect 28252 7646 28254 7698
rect 28306 7646 28532 7698
rect 28252 7644 28532 7646
rect 28252 7634 28308 7644
rect 25676 7422 25678 7474
rect 25730 7422 25732 7474
rect 25676 7410 25732 7422
rect 25564 6638 25566 6690
rect 25618 6638 25620 6690
rect 25564 6626 25620 6638
rect 25900 6804 25956 6814
rect 24332 6468 24388 6478
rect 24332 6374 24388 6412
rect 22764 6066 22820 6076
rect 23772 6132 23828 6142
rect 23772 6038 23828 6076
rect 22988 6020 23044 6030
rect 22428 5346 22484 5964
rect 22428 5294 22430 5346
rect 22482 5294 22484 5346
rect 22428 5282 22484 5294
rect 22876 6018 23044 6020
rect 22876 5966 22990 6018
rect 23042 5966 23044 6018
rect 22876 5964 23044 5966
rect 21644 5236 21700 5246
rect 20300 4900 20356 4910
rect 20300 4806 20356 4844
rect 21084 4900 21140 4910
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19292 4386 19348 4396
rect 19852 4452 19908 4462
rect 17388 4286 17390 4338
rect 17442 4286 17444 4338
rect 17388 4274 17444 4286
rect 19516 4338 19572 4350
rect 19516 4286 19518 4338
rect 19570 4286 19572 4338
rect 15372 4174 15374 4226
rect 15426 4174 15428 4226
rect 15372 4162 15428 4174
rect 14476 3726 14478 3778
rect 14530 3726 14532 3778
rect 14476 3714 14532 3726
rect 19516 4116 19572 4286
rect 19852 4226 19908 4396
rect 19852 4174 19854 4226
rect 19906 4174 19908 4226
rect 19852 4162 19908 4174
rect 14252 3614 14254 3666
rect 14306 3614 14308 3666
rect 14252 3602 14308 3614
rect 12684 3490 12740 3500
rect 14028 3556 14084 3566
rect 14028 3462 14084 3500
rect 19516 3556 19572 4060
rect 19516 3490 19572 3500
rect 21084 3442 21140 4844
rect 21532 4340 21588 4350
rect 21644 4340 21700 5180
rect 22204 5124 22260 5134
rect 22204 5030 22260 5068
rect 21532 4338 21644 4340
rect 21532 4286 21534 4338
rect 21586 4286 21644 4338
rect 21532 4284 21644 4286
rect 21532 4274 21588 4284
rect 21644 4246 21700 4284
rect 22316 4340 22372 4350
rect 22316 4246 22372 4284
rect 21420 4228 21476 4238
rect 21420 4134 21476 4172
rect 21196 4116 21252 4126
rect 21196 4114 21364 4116
rect 21196 4062 21198 4114
rect 21250 4062 21364 4114
rect 21196 4060 21364 4062
rect 21196 4050 21252 4060
rect 21308 3554 21364 4060
rect 21308 3502 21310 3554
rect 21362 3502 21364 3554
rect 21308 3490 21364 3502
rect 21084 3390 21086 3442
rect 21138 3390 21140 3442
rect 21084 3378 21140 3390
rect 22876 3442 22932 5964
rect 22988 5954 23044 5964
rect 25228 6020 25284 6030
rect 25228 5926 25284 5964
rect 24332 5908 24388 5918
rect 23996 5794 24052 5806
rect 23996 5742 23998 5794
rect 24050 5742 24052 5794
rect 23212 4900 23268 4910
rect 23212 4806 23268 4844
rect 23772 4340 23828 4350
rect 23996 4340 24052 5742
rect 23772 4338 24052 4340
rect 23772 4286 23774 4338
rect 23826 4286 24052 4338
rect 23772 4284 24052 4286
rect 24332 4452 24388 5852
rect 24444 5906 24500 5918
rect 24444 5854 24446 5906
rect 24498 5854 24500 5906
rect 24444 5124 24500 5854
rect 25340 5682 25396 5694
rect 25340 5630 25342 5682
rect 25394 5630 25396 5682
rect 25340 5124 25396 5630
rect 25452 5124 25508 5134
rect 25340 5122 25508 5124
rect 25340 5070 25454 5122
rect 25506 5070 25508 5122
rect 25340 5068 25508 5070
rect 24444 5058 24500 5068
rect 25452 5058 25508 5068
rect 25900 5122 25956 6748
rect 26908 6468 26964 6478
rect 26908 6130 26964 6412
rect 28140 6468 28196 6478
rect 28140 6374 28196 6412
rect 26908 6078 26910 6130
rect 26962 6078 26964 6130
rect 26908 6066 26964 6078
rect 28476 6130 28532 7644
rect 28812 7698 28868 7868
rect 28812 7646 28814 7698
rect 28866 7646 28868 7698
rect 28812 7634 28868 7646
rect 29148 7474 29204 9774
rect 30604 9604 30660 9614
rect 30604 9042 30660 9548
rect 30604 8990 30606 9042
rect 30658 8990 30660 9042
rect 30604 8978 30660 8990
rect 29820 8932 29876 8942
rect 29820 8838 29876 8876
rect 30268 8820 30324 8830
rect 29932 8818 30324 8820
rect 29932 8766 30270 8818
rect 30322 8766 30324 8818
rect 29932 8764 30324 8766
rect 29260 8372 29316 8382
rect 29260 8278 29316 8316
rect 29932 8258 29988 8764
rect 30268 8754 30324 8764
rect 30828 8428 30884 10556
rect 30940 10500 30996 10510
rect 30940 10406 30996 10444
rect 31388 9604 31444 12012
rect 32284 10836 32340 12126
rect 32620 12178 32676 12910
rect 32844 12964 32900 17388
rect 32956 15764 33012 19180
rect 33292 19236 33348 20524
rect 33404 20514 33460 20524
rect 33404 20132 33460 20142
rect 33404 20018 33460 20076
rect 33404 19966 33406 20018
rect 33458 19966 33460 20018
rect 33404 19460 33460 19966
rect 33404 19394 33460 19404
rect 33292 19142 33348 19180
rect 33404 18562 33460 18574
rect 33404 18510 33406 18562
rect 33458 18510 33460 18562
rect 33068 18452 33124 18462
rect 33068 18358 33124 18396
rect 33404 18340 33460 18510
rect 33628 18452 33684 18462
rect 33628 18340 33684 18396
rect 33404 18284 33684 18340
rect 33068 17666 33124 17678
rect 33516 17668 33572 17678
rect 33068 17614 33070 17666
rect 33122 17614 33124 17666
rect 33068 17556 33124 17614
rect 33068 17490 33124 17500
rect 33404 17666 33572 17668
rect 33404 17614 33518 17666
rect 33570 17614 33572 17666
rect 33404 17612 33572 17614
rect 33404 17444 33460 17612
rect 33516 17602 33572 17612
rect 33404 16882 33460 17388
rect 33404 16830 33406 16882
rect 33458 16830 33460 16882
rect 33404 16818 33460 16830
rect 33068 16324 33124 16334
rect 33628 16324 33684 18284
rect 33852 17780 33908 20524
rect 33964 20514 34020 20524
rect 34188 20132 34244 20142
rect 34300 20132 34356 20972
rect 35196 20916 35252 20972
rect 35308 20916 35364 20926
rect 35196 20914 35364 20916
rect 35196 20862 35310 20914
rect 35362 20862 35364 20914
rect 35196 20860 35364 20862
rect 35308 20850 35364 20860
rect 34748 20802 34804 20814
rect 34748 20750 34750 20802
rect 34802 20750 34804 20802
rect 34412 20692 34468 20702
rect 34748 20692 34804 20750
rect 34412 20690 34804 20692
rect 34412 20638 34414 20690
rect 34466 20638 34804 20690
rect 34412 20636 34804 20638
rect 34412 20626 34468 20636
rect 34188 20130 34356 20132
rect 34188 20078 34190 20130
rect 34242 20078 34356 20130
rect 34188 20076 34356 20078
rect 34188 20066 34244 20076
rect 33964 20020 34020 20030
rect 33964 19926 34020 19964
rect 34636 20018 34692 20030
rect 34636 19966 34638 20018
rect 34690 19966 34692 20018
rect 34412 19908 34468 19918
rect 34300 19906 34468 19908
rect 34300 19854 34414 19906
rect 34466 19854 34468 19906
rect 34300 19852 34468 19854
rect 34300 19460 34356 19852
rect 34412 19842 34468 19852
rect 33964 19404 34356 19460
rect 33964 19346 34020 19404
rect 33964 19294 33966 19346
rect 34018 19294 34020 19346
rect 33964 19282 34020 19294
rect 34076 18450 34132 18462
rect 34076 18398 34078 18450
rect 34130 18398 34132 18450
rect 34076 18340 34132 18398
rect 34076 18274 34132 18284
rect 34300 18450 34356 18462
rect 34300 18398 34302 18450
rect 34354 18398 34356 18450
rect 34300 18340 34356 18398
rect 34636 18452 34692 19966
rect 34748 19236 34804 20636
rect 34972 20802 35028 20814
rect 34972 20750 34974 20802
rect 35026 20750 35028 20802
rect 34972 20692 35028 20750
rect 34972 20626 35028 20636
rect 35196 20692 35252 20702
rect 35196 20598 35252 20636
rect 35420 20580 35476 20590
rect 35420 20486 35476 20524
rect 35532 20242 35588 21308
rect 35644 21298 35700 21308
rect 35532 20190 35534 20242
rect 35586 20190 35588 20242
rect 35532 20178 35588 20190
rect 35196 20132 35252 20142
rect 35196 20018 35252 20076
rect 35196 19966 35198 20018
rect 35250 19966 35252 20018
rect 35196 19954 35252 19966
rect 35420 20020 35476 20030
rect 35420 19926 35476 19964
rect 35644 20018 35700 20030
rect 35644 19966 35646 20018
rect 35698 19966 35700 20018
rect 34972 19908 35028 19918
rect 34972 19814 35028 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34748 19170 34804 19180
rect 35644 19124 35700 19966
rect 35644 19058 35700 19068
rect 34860 18452 34916 18462
rect 34692 18450 34916 18452
rect 34692 18398 34862 18450
rect 34914 18398 34916 18450
rect 34692 18396 34916 18398
rect 34636 18358 34692 18396
rect 34860 18386 34916 18396
rect 35308 18452 35364 18462
rect 35308 18358 35364 18396
rect 35532 18450 35588 18462
rect 35532 18398 35534 18450
rect 35586 18398 35588 18450
rect 34524 18340 34580 18350
rect 34300 18274 34356 18284
rect 34412 18338 34580 18340
rect 34412 18286 34526 18338
rect 34578 18286 34580 18338
rect 34412 18284 34580 18286
rect 33852 17714 33908 17724
rect 34300 17556 34356 17566
rect 34300 17462 34356 17500
rect 34188 16996 34244 17006
rect 34412 16996 34468 18284
rect 34524 18274 34580 18284
rect 35084 18338 35140 18350
rect 35084 18286 35086 18338
rect 35138 18286 35140 18338
rect 35084 17556 35140 18286
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35084 17490 35140 17500
rect 34188 16994 34468 16996
rect 34188 16942 34190 16994
rect 34242 16942 34468 16994
rect 34188 16940 34468 16942
rect 34188 16930 34244 16940
rect 35532 16884 35588 18398
rect 35532 16818 35588 16828
rect 34300 16772 34356 16782
rect 33964 16324 34020 16334
rect 33628 16322 34020 16324
rect 33628 16270 33966 16322
rect 34018 16270 34020 16322
rect 33628 16268 34020 16270
rect 33068 16210 33124 16268
rect 33964 16258 34020 16268
rect 34300 16322 34356 16716
rect 35756 16772 35812 23884
rect 36316 23826 36372 23838
rect 36316 23774 36318 23826
rect 36370 23774 36372 23826
rect 36204 23714 36260 23726
rect 36204 23662 36206 23714
rect 36258 23662 36260 23714
rect 36204 23604 36260 23662
rect 36204 23538 36260 23548
rect 36316 23492 36372 23774
rect 36540 23492 36596 25230
rect 37212 24948 37268 24958
rect 37212 23826 37268 24892
rect 37548 23938 37604 25678
rect 37884 25618 37940 25630
rect 37884 25566 37886 25618
rect 37938 25566 37940 25618
rect 37884 25284 37940 25566
rect 37884 25218 37940 25228
rect 37996 24946 38052 26348
rect 38556 25732 38612 26910
rect 38892 26850 38948 26862
rect 38892 26798 38894 26850
rect 38946 26798 38948 26850
rect 38892 26404 38948 26798
rect 38892 26338 38948 26348
rect 38892 26178 38948 26190
rect 38892 26126 38894 26178
rect 38946 26126 38948 26178
rect 38668 25732 38724 25742
rect 38556 25730 38724 25732
rect 38556 25678 38670 25730
rect 38722 25678 38724 25730
rect 38556 25676 38724 25678
rect 38668 25666 38724 25676
rect 38780 25508 38836 25518
rect 38892 25508 38948 26126
rect 39004 25844 39060 27692
rect 41020 27074 41076 27086
rect 41020 27022 41022 27074
rect 41074 27022 41076 27074
rect 39228 26962 39284 26974
rect 39228 26910 39230 26962
rect 39282 26910 39284 26962
rect 39228 26066 39284 26910
rect 40796 26964 40852 26974
rect 41020 26964 41076 27022
rect 40796 26962 41076 26964
rect 40796 26910 40798 26962
rect 40850 26910 41076 26962
rect 40796 26908 41076 26910
rect 41804 27074 41860 27692
rect 41804 27022 41806 27074
rect 41858 27022 41860 27074
rect 39228 26014 39230 26066
rect 39282 26014 39284 26066
rect 39228 26002 39284 26014
rect 39452 26290 39508 26302
rect 39452 26238 39454 26290
rect 39506 26238 39508 26290
rect 39004 25788 39284 25844
rect 38780 25506 38948 25508
rect 38780 25454 38782 25506
rect 38834 25454 38948 25506
rect 38780 25452 38948 25454
rect 37996 24894 37998 24946
rect 38050 24894 38052 24946
rect 37996 24882 38052 24894
rect 38444 25284 38500 25294
rect 38780 25284 38836 25452
rect 38500 25228 38836 25284
rect 38332 24724 38388 24734
rect 38332 24610 38388 24668
rect 38332 24558 38334 24610
rect 38386 24558 38388 24610
rect 38332 24546 38388 24558
rect 37548 23886 37550 23938
rect 37602 23886 37604 23938
rect 37548 23874 37604 23886
rect 37212 23774 37214 23826
rect 37266 23774 37268 23826
rect 37212 23762 37268 23774
rect 36988 23604 37044 23614
rect 37044 23548 37156 23604
rect 36988 23538 37044 23548
rect 36316 23436 36932 23492
rect 35980 23380 36036 23390
rect 35868 23156 35924 23166
rect 35868 22930 35924 23100
rect 35980 23154 36036 23324
rect 35980 23102 35982 23154
rect 36034 23102 36036 23154
rect 35980 23090 36036 23102
rect 36092 23268 36148 23278
rect 35868 22878 35870 22930
rect 35922 22878 35924 22930
rect 35868 21812 35924 22878
rect 36092 22708 36148 23212
rect 36540 23268 36596 23278
rect 36540 23174 36596 23212
rect 36092 22642 36148 22652
rect 36316 23154 36372 23166
rect 36316 23102 36318 23154
rect 36370 23102 36372 23154
rect 35980 22372 36036 22382
rect 36036 22316 36148 22372
rect 35980 22306 36036 22316
rect 35868 21746 35924 21756
rect 36092 21810 36148 22316
rect 36092 21758 36094 21810
rect 36146 21758 36148 21810
rect 36092 21746 36148 21758
rect 35868 21028 35924 21038
rect 36316 21028 36372 23102
rect 36764 23156 36820 23166
rect 36764 23062 36820 23100
rect 36428 23042 36484 23054
rect 36428 22990 36430 23042
rect 36482 22990 36484 23042
rect 36428 21924 36484 22990
rect 36876 22932 36932 23436
rect 36988 23380 37044 23390
rect 36988 23266 37044 23324
rect 36988 23214 36990 23266
rect 37042 23214 37044 23266
rect 36988 23202 37044 23214
rect 37100 23044 37156 23548
rect 37884 23268 37940 23278
rect 37772 23156 37828 23166
rect 36428 21858 36484 21868
rect 36764 22876 36932 22932
rect 36988 22988 37156 23044
rect 37436 23100 37772 23156
rect 36540 21700 36596 21738
rect 36540 21634 36596 21644
rect 35868 20934 35924 20972
rect 35980 20972 36372 21028
rect 36428 21586 36484 21598
rect 36428 21534 36430 21586
rect 36482 21534 36484 21586
rect 35980 20914 36036 20972
rect 35980 20862 35982 20914
rect 36034 20862 36036 20914
rect 35980 20850 36036 20862
rect 35980 20244 36036 20254
rect 35980 20018 36036 20188
rect 35980 19966 35982 20018
rect 36034 19966 36036 20018
rect 35980 19012 36036 19966
rect 36092 19346 36148 20972
rect 36428 20804 36484 21534
rect 36652 21588 36708 21598
rect 36652 21494 36708 21532
rect 36092 19294 36094 19346
rect 36146 19294 36148 19346
rect 36092 19282 36148 19294
rect 36316 20748 36484 20804
rect 36540 21476 36596 21486
rect 35980 18956 36148 19012
rect 35868 18562 35924 18574
rect 35868 18510 35870 18562
rect 35922 18510 35924 18562
rect 35868 17668 35924 18510
rect 35868 17602 35924 17612
rect 35756 16706 35812 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34300 16270 34302 16322
rect 34354 16270 34356 16322
rect 34300 16258 34356 16270
rect 33068 16158 33070 16210
rect 33122 16158 33124 16210
rect 33068 16146 33124 16158
rect 32956 15698 33012 15708
rect 34300 16098 34356 16110
rect 34300 16046 34302 16098
rect 34354 16046 34356 16098
rect 34300 15876 34356 16046
rect 34300 15148 34356 15820
rect 35532 15764 35588 15774
rect 34076 15092 34132 15102
rect 34300 15092 34692 15148
rect 34076 14644 34132 15036
rect 33964 14642 34132 14644
rect 33964 14590 34078 14642
rect 34130 14590 34132 14642
rect 33964 14588 34132 14590
rect 33068 13972 33124 13982
rect 33068 13858 33124 13916
rect 33068 13806 33070 13858
rect 33122 13806 33124 13858
rect 33068 13794 33124 13806
rect 33404 13860 33460 13870
rect 33404 13766 33460 13804
rect 32956 13748 33012 13758
rect 32956 13076 33012 13692
rect 33180 13524 33236 13534
rect 32956 13020 33124 13076
rect 32844 12898 32900 12908
rect 32956 12850 33012 12862
rect 32956 12798 32958 12850
rect 33010 12798 33012 12850
rect 32620 12126 32622 12178
rect 32674 12126 32676 12178
rect 32620 12114 32676 12126
rect 32844 12738 32900 12750
rect 32844 12686 32846 12738
rect 32898 12686 32900 12738
rect 32396 12068 32452 12078
rect 32396 11974 32452 12012
rect 32844 11508 32900 12686
rect 32956 11620 33012 12798
rect 33068 12404 33124 13020
rect 33180 12962 33236 13468
rect 33180 12910 33182 12962
rect 33234 12910 33236 12962
rect 33180 12898 33236 12910
rect 33516 12964 33572 12974
rect 33628 12964 33684 12974
rect 33572 12962 33684 12964
rect 33572 12910 33630 12962
rect 33682 12910 33684 12962
rect 33572 12908 33684 12910
rect 33068 12348 33236 12404
rect 32956 11554 33012 11564
rect 33068 12178 33124 12190
rect 33068 12126 33070 12178
rect 33122 12126 33124 12178
rect 32844 11442 32900 11452
rect 32620 11394 32676 11406
rect 32620 11342 32622 11394
rect 32674 11342 32676 11394
rect 32620 11284 32676 11342
rect 32620 11218 32676 11228
rect 33068 11394 33124 12126
rect 33068 11342 33070 11394
rect 33122 11342 33124 11394
rect 32284 10770 32340 10780
rect 32396 11170 32452 11182
rect 32396 11118 32398 11170
rect 32450 11118 32452 11170
rect 32396 11060 32452 11118
rect 33068 11060 33124 11342
rect 32396 11004 33124 11060
rect 31724 10724 31780 10734
rect 31724 10630 31780 10668
rect 31836 10498 31892 10510
rect 31836 10446 31838 10498
rect 31890 10446 31892 10498
rect 31836 9940 31892 10446
rect 32060 9940 32116 9950
rect 31836 9938 32116 9940
rect 31836 9886 32062 9938
rect 32114 9886 32116 9938
rect 31836 9884 32116 9886
rect 32060 9874 32116 9884
rect 32396 9716 32452 11004
rect 31388 9538 31444 9548
rect 32060 9660 32452 9716
rect 30940 9156 30996 9166
rect 30940 9062 30996 9100
rect 31388 9154 31444 9166
rect 31388 9102 31390 9154
rect 31442 9102 31444 9154
rect 29932 8206 29934 8258
rect 29986 8206 29988 8258
rect 29932 8194 29988 8206
rect 30044 8372 30100 8382
rect 29596 8036 29652 8046
rect 30044 8036 30100 8316
rect 30492 8372 30884 8428
rect 30268 8260 30324 8270
rect 30492 8260 30548 8372
rect 30268 8258 30548 8260
rect 30268 8206 30270 8258
rect 30322 8206 30548 8258
rect 30268 8204 30548 8206
rect 30268 8194 30324 8204
rect 30380 8036 30436 8046
rect 29596 8034 29876 8036
rect 29596 7982 29598 8034
rect 29650 7982 29876 8034
rect 29596 7980 29876 7982
rect 30044 8034 30436 8036
rect 30044 7982 30382 8034
rect 30434 7982 30436 8034
rect 30044 7980 30436 7982
rect 30492 8036 30548 8204
rect 30604 8260 30660 8270
rect 30604 8258 31332 8260
rect 30604 8206 30606 8258
rect 30658 8206 31332 8258
rect 30604 8204 31332 8206
rect 30604 8194 30660 8204
rect 31276 8146 31332 8204
rect 31276 8094 31278 8146
rect 31330 8094 31332 8146
rect 31276 8082 31332 8094
rect 30828 8036 30884 8046
rect 30492 8034 30884 8036
rect 30492 7982 30830 8034
rect 30882 7982 30884 8034
rect 30492 7980 30884 7982
rect 29596 7970 29652 7980
rect 29820 7586 29876 7980
rect 30380 7700 30436 7980
rect 30828 7970 30884 7980
rect 30940 8034 30996 8046
rect 30940 7982 30942 8034
rect 30994 7982 30996 8034
rect 30380 7634 30436 7644
rect 29820 7534 29822 7586
rect 29874 7534 29876 7586
rect 29820 7522 29876 7534
rect 29148 7422 29150 7474
rect 29202 7422 29204 7474
rect 28588 6804 28644 6814
rect 28588 6710 28644 6748
rect 29148 6692 29204 7422
rect 30828 6804 30884 6814
rect 30940 6804 30996 7982
rect 31052 8036 31108 8046
rect 31052 7942 31108 7980
rect 31388 7252 31444 9102
rect 31724 9156 31780 9166
rect 31780 9100 31892 9156
rect 31724 9090 31780 9100
rect 31836 9042 31892 9100
rect 31836 8990 31838 9042
rect 31890 8990 31892 9042
rect 31836 8978 31892 8990
rect 32060 8258 32116 9660
rect 32508 9604 32564 9614
rect 32508 9510 32564 9548
rect 33180 9268 33236 12348
rect 33516 11284 33572 12908
rect 33628 12898 33684 12908
rect 33964 12516 34020 14588
rect 34076 14578 34132 14588
rect 34412 14420 34468 14430
rect 34188 14418 34468 14420
rect 34188 14366 34414 14418
rect 34466 14366 34468 14418
rect 34188 14364 34468 14366
rect 34188 13860 34244 14364
rect 34412 14354 34468 14364
rect 34636 14418 34692 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34636 14366 34638 14418
rect 34690 14366 34692 14418
rect 34636 14354 34692 14366
rect 34748 14642 34804 14654
rect 34748 14590 34750 14642
rect 34802 14590 34804 14642
rect 34188 13766 34244 13804
rect 34748 13858 34804 14590
rect 34748 13806 34750 13858
rect 34802 13806 34804 13858
rect 34748 13794 34804 13806
rect 35084 13972 35140 13982
rect 35084 13858 35140 13916
rect 35084 13806 35086 13858
rect 35138 13806 35140 13858
rect 35084 13794 35140 13806
rect 34524 13746 34580 13758
rect 34524 13694 34526 13746
rect 34578 13694 34580 13746
rect 34300 13634 34356 13646
rect 34300 13582 34302 13634
rect 34354 13582 34356 13634
rect 34300 13074 34356 13582
rect 34524 13188 34580 13694
rect 35420 13748 35476 13758
rect 35532 13748 35588 15708
rect 36092 15148 36148 18956
rect 36316 18900 36372 20748
rect 36428 20580 36484 20590
rect 36540 20580 36596 21420
rect 36428 20578 36596 20580
rect 36428 20526 36430 20578
rect 36482 20526 36596 20578
rect 36428 20524 36596 20526
rect 36428 20244 36484 20524
rect 36428 20178 36484 20188
rect 36540 20020 36596 20030
rect 36540 19926 36596 19964
rect 36428 19124 36484 19134
rect 36484 19068 36708 19124
rect 36428 19058 36484 19068
rect 36316 18844 36596 18900
rect 36204 18450 36260 18462
rect 36204 18398 36206 18450
rect 36258 18398 36260 18450
rect 36204 18228 36260 18398
rect 36540 18452 36596 18844
rect 36540 18358 36596 18396
rect 36652 18562 36708 19068
rect 36652 18510 36654 18562
rect 36706 18510 36708 18562
rect 36652 18228 36708 18510
rect 36204 18162 36260 18172
rect 36428 18172 36708 18228
rect 36428 17778 36484 18172
rect 36428 17726 36430 17778
rect 36482 17726 36484 17778
rect 36428 17714 36484 17726
rect 36316 17556 36372 17566
rect 36316 16770 36372 17500
rect 36764 16882 36820 22876
rect 36876 22708 36932 22718
rect 36876 21586 36932 22652
rect 36988 22370 37044 22988
rect 36988 22318 36990 22370
rect 37042 22318 37044 22370
rect 36988 22306 37044 22318
rect 37100 22596 37156 22606
rect 36876 21534 36878 21586
rect 36930 21534 36932 21586
rect 36876 21522 36932 21534
rect 37100 21586 37156 22540
rect 37436 22370 37492 23100
rect 37772 23062 37828 23100
rect 37436 22318 37438 22370
rect 37490 22318 37492 22370
rect 37436 22306 37492 22318
rect 37884 22372 37940 23212
rect 37884 22306 37940 22316
rect 38444 23042 38500 25228
rect 38892 23492 38948 23502
rect 38892 23154 38948 23436
rect 38892 23102 38894 23154
rect 38946 23102 38948 23154
rect 38892 23090 38948 23102
rect 38444 22990 38446 23042
rect 38498 22990 38500 23042
rect 37212 22260 37268 22270
rect 37212 22166 37268 22204
rect 37324 22148 37380 22158
rect 37324 22054 37380 22092
rect 37548 22146 37604 22158
rect 37548 22094 37550 22146
rect 37602 22094 37604 22146
rect 37100 21534 37102 21586
rect 37154 21534 37156 21586
rect 37100 21522 37156 21534
rect 37548 21028 37604 22094
rect 38444 21812 38500 22990
rect 38556 22596 38612 22606
rect 38556 22036 38612 22540
rect 39116 22370 39172 22382
rect 39116 22318 39118 22370
rect 39170 22318 39172 22370
rect 38668 22260 38724 22270
rect 39116 22260 39172 22318
rect 38668 22258 39172 22260
rect 38668 22206 38670 22258
rect 38722 22206 39172 22258
rect 38668 22204 39172 22206
rect 38668 22194 38724 22204
rect 38556 21980 38724 22036
rect 38556 21812 38612 21822
rect 38444 21756 38556 21812
rect 38556 21746 38612 21756
rect 37548 20962 37604 20972
rect 38108 21588 38164 21598
rect 37100 20916 37156 20926
rect 37100 20822 37156 20860
rect 38108 20802 38164 21532
rect 38108 20750 38110 20802
rect 38162 20750 38164 20802
rect 37212 20692 37268 20702
rect 37212 20598 37268 20636
rect 37660 20690 37716 20702
rect 37660 20638 37662 20690
rect 37714 20638 37716 20690
rect 37100 20580 37156 20590
rect 37100 20244 37156 20524
rect 37436 20578 37492 20590
rect 37436 20526 37438 20578
rect 37490 20526 37492 20578
rect 37100 20188 37268 20244
rect 36876 20020 36932 20030
rect 37100 20020 37156 20030
rect 36932 19964 37044 20020
rect 36876 19954 36932 19964
rect 36988 19458 37044 19964
rect 36988 19406 36990 19458
rect 37042 19406 37044 19458
rect 36988 19394 37044 19406
rect 37100 19346 37156 19964
rect 37100 19294 37102 19346
rect 37154 19294 37156 19346
rect 37100 19282 37156 19294
rect 37100 18338 37156 18350
rect 37100 18286 37102 18338
rect 37154 18286 37156 18338
rect 37100 18228 37156 18286
rect 37100 18162 37156 18172
rect 37212 18340 37268 20188
rect 37436 20132 37492 20526
rect 37436 20066 37492 20076
rect 37660 19908 37716 20638
rect 38108 20020 38164 20750
rect 38668 20802 38724 21980
rect 39116 20916 39172 22204
rect 39116 20850 39172 20860
rect 38668 20750 38670 20802
rect 38722 20750 38724 20802
rect 38668 20738 38724 20750
rect 39228 20692 39284 25788
rect 39452 25506 39508 26238
rect 39452 25454 39454 25506
rect 39506 25454 39508 25506
rect 39452 24724 39508 25454
rect 39452 24658 39508 24668
rect 40684 23938 40740 23950
rect 40684 23886 40686 23938
rect 40738 23886 40740 23938
rect 39788 23492 39844 23502
rect 39788 23378 39844 23436
rect 39788 23326 39790 23378
rect 39842 23326 39844 23378
rect 39788 23314 39844 23326
rect 39900 23268 39956 23278
rect 39452 22372 39508 22382
rect 39452 22278 39508 22316
rect 39788 21812 39844 21822
rect 39788 21718 39844 21756
rect 38108 19954 38164 19964
rect 39004 20636 39284 20692
rect 37660 19124 37716 19852
rect 37660 19058 37716 19068
rect 37100 17892 37156 17902
rect 37212 17892 37268 18284
rect 37100 17890 37268 17892
rect 37100 17838 37102 17890
rect 37154 17838 37268 17890
rect 37100 17836 37268 17838
rect 37100 17826 37156 17836
rect 37548 17780 37604 17790
rect 37548 17686 37604 17724
rect 38892 17668 38948 17678
rect 36988 17556 37044 17566
rect 36988 17462 37044 17500
rect 37436 17442 37492 17454
rect 37436 17390 37438 17442
rect 37490 17390 37492 17442
rect 36764 16830 36766 16882
rect 36818 16830 36820 16882
rect 36764 16818 36820 16830
rect 37324 16884 37380 16894
rect 37436 16884 37492 17390
rect 38892 17108 38948 17612
rect 38892 17042 38948 17052
rect 37324 16882 37492 16884
rect 37324 16830 37326 16882
rect 37378 16830 37492 16882
rect 37324 16828 37492 16830
rect 37324 16818 37380 16828
rect 36316 16718 36318 16770
rect 36370 16718 36372 16770
rect 36316 16706 36372 16718
rect 36540 16772 36596 16782
rect 35980 15092 36148 15148
rect 36540 15204 36596 16716
rect 39004 16324 39060 20636
rect 39116 20242 39172 20254
rect 39116 20190 39118 20242
rect 39170 20190 39172 20242
rect 39116 20132 39172 20190
rect 39900 20188 39956 23212
rect 40684 23156 40740 23886
rect 40348 23044 40404 23054
rect 40348 22950 40404 22988
rect 40684 22484 40740 23100
rect 40684 22418 40740 22428
rect 39116 20066 39172 20076
rect 39788 20132 39956 20188
rect 40236 21474 40292 21486
rect 40236 21422 40238 21474
rect 40290 21422 40292 21474
rect 40012 20132 40068 20142
rect 39676 20020 39732 20030
rect 39676 19926 39732 19964
rect 39788 18452 39844 20132
rect 40012 20038 40068 20076
rect 40236 19348 40292 21422
rect 40348 20132 40404 20142
rect 40348 20038 40404 20076
rect 40236 19282 40292 19292
rect 40684 19236 40740 19246
rect 40684 19142 40740 19180
rect 40236 19124 40292 19134
rect 40236 19030 40292 19068
rect 40348 19012 40404 19022
rect 40348 19010 40740 19012
rect 40348 18958 40350 19010
rect 40402 18958 40740 19010
rect 40348 18956 40740 18958
rect 40348 18946 40404 18956
rect 40684 18676 40740 18956
rect 40796 18900 40852 26908
rect 41020 26290 41076 26302
rect 41020 26238 41022 26290
rect 41074 26238 41076 26290
rect 41020 21364 41076 26238
rect 41804 26290 41860 27022
rect 43148 27748 43204 27758
rect 43148 26964 43204 27692
rect 43596 27748 43652 27758
rect 43596 27654 43652 27692
rect 43148 26898 43204 26908
rect 41804 26238 41806 26290
rect 41858 26238 41860 26290
rect 41804 26226 41860 26238
rect 43820 26068 43876 27918
rect 43932 26852 43988 36204
rect 44044 35026 44100 35038
rect 44044 34974 44046 35026
rect 44098 34974 44100 35026
rect 44044 33346 44100 34974
rect 44044 33294 44046 33346
rect 44098 33294 44100 33346
rect 44044 33282 44100 33294
rect 44380 31948 44436 36316
rect 44492 36260 44548 41916
rect 44492 36194 44548 36204
rect 44268 31892 44436 31948
rect 44492 34020 44548 34030
rect 44044 31778 44100 31790
rect 44044 31726 44046 31778
rect 44098 31726 44100 31778
rect 44044 28754 44100 31726
rect 44044 28702 44046 28754
rect 44098 28702 44100 28754
rect 44044 28690 44100 28702
rect 44156 27858 44212 27870
rect 44156 27806 44158 27858
rect 44210 27806 44212 27858
rect 44156 27748 44212 27806
rect 44156 27682 44212 27692
rect 44268 27524 44324 31892
rect 44156 27468 44324 27524
rect 44156 27186 44212 27468
rect 44156 27134 44158 27186
rect 44210 27134 44212 27186
rect 44156 27122 44212 27134
rect 44268 26964 44324 26974
rect 43932 26796 44212 26852
rect 44156 26514 44212 26796
rect 44156 26462 44158 26514
rect 44210 26462 44212 26514
rect 44156 26450 44212 26462
rect 43820 26002 43876 26012
rect 41468 25620 41524 25630
rect 41468 25526 41524 25564
rect 44044 25620 44100 25630
rect 42252 25394 42308 25406
rect 42252 25342 42254 25394
rect 42306 25342 42308 25394
rect 41356 25284 41412 25294
rect 41244 25282 41412 25284
rect 41244 25230 41358 25282
rect 41410 25230 41412 25282
rect 41244 25228 41412 25230
rect 41244 23938 41300 25228
rect 41356 25218 41412 25228
rect 41916 25282 41972 25294
rect 41916 25230 41918 25282
rect 41970 25230 41972 25282
rect 41244 23886 41246 23938
rect 41298 23886 41300 23938
rect 41244 23874 41300 23886
rect 41468 24724 41524 24734
rect 41468 23156 41524 24668
rect 41692 24610 41748 24622
rect 41692 24558 41694 24610
rect 41746 24558 41748 24610
rect 41580 23156 41636 23166
rect 41468 23100 41580 23156
rect 41580 23062 41636 23100
rect 41020 21298 41076 21308
rect 41692 23044 41748 24558
rect 41692 21474 41748 22988
rect 41916 22146 41972 25230
rect 42252 24610 42308 25342
rect 43036 24834 43092 24846
rect 43036 24782 43038 24834
rect 43090 24782 43092 24834
rect 42252 24558 42254 24610
rect 42306 24558 42308 24610
rect 42252 24546 42308 24558
rect 42700 24722 42756 24734
rect 42700 24670 42702 24722
rect 42754 24670 42756 24722
rect 42476 23268 42532 23278
rect 42700 23268 42756 24670
rect 43036 23828 43092 24782
rect 44044 24050 44100 25564
rect 44044 23998 44046 24050
rect 44098 23998 44100 24050
rect 44044 23986 44100 23998
rect 44156 25284 44212 25294
rect 44268 25284 44324 26908
rect 44156 25282 44324 25284
rect 44156 25230 44158 25282
rect 44210 25230 44324 25282
rect 44156 25228 44324 25230
rect 43484 23828 43540 23838
rect 44156 23828 44212 25228
rect 43036 23826 43540 23828
rect 43036 23774 43486 23826
rect 43538 23774 43540 23826
rect 43036 23772 43540 23774
rect 43484 23762 43540 23772
rect 44044 23772 44212 23828
rect 43820 23268 43876 23278
rect 42476 23266 42756 23268
rect 42476 23214 42478 23266
rect 42530 23214 42756 23266
rect 42476 23212 42756 23214
rect 43708 23266 43876 23268
rect 43708 23214 43822 23266
rect 43874 23214 43876 23266
rect 43708 23212 43876 23214
rect 42476 23202 42532 23212
rect 42812 23156 42868 23166
rect 42812 23062 42868 23100
rect 43260 23154 43316 23166
rect 43260 23102 43262 23154
rect 43314 23102 43316 23154
rect 42364 22484 42420 22494
rect 42364 22390 42420 22428
rect 41916 22094 41918 22146
rect 41970 22094 41972 22146
rect 41916 22082 41972 22094
rect 41916 21588 41972 21598
rect 41916 21586 42084 21588
rect 41916 21534 41918 21586
rect 41970 21534 42084 21586
rect 41916 21532 42084 21534
rect 41916 21522 41972 21532
rect 41692 21422 41694 21474
rect 41746 21422 41748 21474
rect 41468 20916 41524 20926
rect 41468 20822 41524 20860
rect 41132 20580 41188 20590
rect 41132 20486 41188 20524
rect 40908 20132 40964 20142
rect 40908 20038 40964 20076
rect 41692 19906 41748 21422
rect 42028 21028 42084 21532
rect 42252 21364 42308 21374
rect 42252 21270 42308 21308
rect 42028 20972 42420 21028
rect 41804 20020 41860 20030
rect 42028 20020 42084 20972
rect 42364 20914 42420 20972
rect 42364 20862 42366 20914
rect 42418 20862 42420 20914
rect 42364 20850 42420 20862
rect 42924 20804 42980 20814
rect 43260 20804 43316 23102
rect 43372 21364 43428 21374
rect 43428 21308 43540 21364
rect 43372 21298 43428 21308
rect 42924 20802 43316 20804
rect 42924 20750 42926 20802
rect 42978 20750 43316 20802
rect 42924 20748 43316 20750
rect 43484 20802 43540 21308
rect 43484 20750 43486 20802
rect 43538 20750 43540 20802
rect 42924 20738 42980 20748
rect 43148 20188 43204 20748
rect 43484 20738 43540 20750
rect 43260 20580 43316 20590
rect 43260 20486 43316 20524
rect 43148 20132 43316 20188
rect 41804 20018 42028 20020
rect 41804 19966 41806 20018
rect 41858 19966 42028 20018
rect 41804 19964 42028 19966
rect 41804 19954 41860 19964
rect 41692 19854 41694 19906
rect 41746 19854 41748 19906
rect 41692 19842 41748 19854
rect 40796 18834 40852 18844
rect 41132 19234 41188 19246
rect 41132 19182 41134 19234
rect 41186 19182 41188 19234
rect 41132 18676 41188 19182
rect 40684 18620 41188 18676
rect 41244 19236 41300 19246
rect 41244 18562 41300 19180
rect 41244 18510 41246 18562
rect 41298 18510 41300 18562
rect 40012 18452 40068 18462
rect 39340 18450 40068 18452
rect 39340 18398 40014 18450
rect 40066 18398 40068 18450
rect 39340 18396 40068 18398
rect 39340 17666 39396 18396
rect 40012 18386 40068 18396
rect 40124 18340 40180 18350
rect 40124 18246 40180 18284
rect 40684 18340 40740 18350
rect 39340 17614 39342 17666
rect 39394 17614 39396 17666
rect 39340 17602 39396 17614
rect 39788 17106 39844 17118
rect 39788 17054 39790 17106
rect 39842 17054 39844 17106
rect 39004 16268 39620 16324
rect 39340 16098 39396 16110
rect 39340 16046 39342 16098
rect 39394 16046 39396 16098
rect 35420 13746 35588 13748
rect 35420 13694 35422 13746
rect 35474 13694 35588 13746
rect 35420 13692 35588 13694
rect 35756 14306 35812 14318
rect 35756 14254 35758 14306
rect 35810 14254 35812 14306
rect 35756 13748 35812 14254
rect 35980 13748 36036 15092
rect 35756 13746 36036 13748
rect 35756 13694 35982 13746
rect 36034 13694 36036 13746
rect 35756 13692 36036 13694
rect 35420 13682 35476 13692
rect 35980 13682 36036 13692
rect 35420 13524 35476 13562
rect 35420 13458 35476 13468
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 34524 13122 34580 13132
rect 34300 13022 34302 13074
rect 34354 13022 34356 13074
rect 34300 13010 34356 13022
rect 36428 13074 36484 13086
rect 36428 13022 36430 13074
rect 36482 13022 36484 13074
rect 36428 12852 36484 13022
rect 36540 13076 36596 15148
rect 38780 15876 38836 15886
rect 39340 15876 39396 16046
rect 38780 15874 39396 15876
rect 38780 15822 38782 15874
rect 38834 15822 39396 15874
rect 38780 15820 39396 15822
rect 36652 13746 36708 13758
rect 36652 13694 36654 13746
rect 36706 13694 36708 13746
rect 36652 13300 36708 13694
rect 38780 13524 38836 15820
rect 39228 15204 39284 15214
rect 39228 15110 39284 15148
rect 39116 13972 39172 13982
rect 39116 13878 39172 13916
rect 38780 13468 39172 13524
rect 36652 13234 36708 13244
rect 37436 13300 37492 13310
rect 36988 13188 37044 13198
rect 37436 13188 37492 13244
rect 36764 13076 36820 13086
rect 36540 13020 36708 13076
rect 36428 12786 36484 12796
rect 33852 12068 33908 12078
rect 33852 11974 33908 12012
rect 33852 11508 33908 11518
rect 33852 11414 33908 11452
rect 33516 11218 33572 11228
rect 33964 10834 34020 12460
rect 36540 12516 36596 12526
rect 33964 10782 33966 10834
rect 34018 10782 34020 10834
rect 33964 10770 34020 10782
rect 34076 12404 34132 12414
rect 34076 10834 34132 12348
rect 36316 12404 36372 12414
rect 36316 12178 36372 12348
rect 36316 12126 36318 12178
rect 36370 12126 36372 12178
rect 36316 12114 36372 12126
rect 36540 12178 36596 12460
rect 36540 12126 36542 12178
rect 36594 12126 36596 12178
rect 36540 12114 36596 12126
rect 35980 12068 36036 12078
rect 35980 12066 36260 12068
rect 35980 12014 35982 12066
rect 36034 12014 36260 12066
rect 35980 12012 36260 12014
rect 35980 12002 36036 12012
rect 36092 11844 36148 11854
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35980 11508 36036 11518
rect 35980 11414 36036 11452
rect 35532 11396 35588 11406
rect 34076 10782 34078 10834
rect 34130 10782 34132 10834
rect 34076 10770 34132 10782
rect 34636 11004 35252 11060
rect 34300 10610 34356 10622
rect 34300 10558 34302 10610
rect 34354 10558 34356 10610
rect 34188 10498 34244 10510
rect 34188 10446 34190 10498
rect 34242 10446 34244 10498
rect 33740 9268 33796 9278
rect 33180 9266 33796 9268
rect 33180 9214 33182 9266
rect 33234 9214 33742 9266
rect 33794 9214 33796 9266
rect 33180 9212 33796 9214
rect 33180 9202 33236 9212
rect 33740 9202 33796 9212
rect 32060 8206 32062 8258
rect 32114 8206 32116 8258
rect 31948 7700 32004 7710
rect 31388 7186 31444 7196
rect 31836 7644 31948 7700
rect 30828 6802 30996 6804
rect 30828 6750 30830 6802
rect 30882 6750 30996 6802
rect 30828 6748 30996 6750
rect 31836 6804 31892 7644
rect 31948 7634 32004 7644
rect 31948 7362 32004 7374
rect 31948 7310 31950 7362
rect 32002 7310 32004 7362
rect 31948 7252 32004 7310
rect 32060 7252 32116 8206
rect 32172 9156 32228 9166
rect 33068 9156 33124 9166
rect 32172 9154 33124 9156
rect 32172 9102 32174 9154
rect 32226 9102 33070 9154
rect 33122 9102 33124 9154
rect 32172 9100 33124 9102
rect 32172 7476 32228 9100
rect 33068 9090 33124 9100
rect 33404 9042 33460 9054
rect 33404 8990 33406 9042
rect 33458 8990 33460 9042
rect 32732 8148 32788 8158
rect 32732 8146 33236 8148
rect 32732 8094 32734 8146
rect 32786 8094 33236 8146
rect 32732 8092 33236 8094
rect 32732 8082 32788 8092
rect 32396 7700 32452 7710
rect 32396 7606 32452 7644
rect 33180 7698 33236 8092
rect 33180 7646 33182 7698
rect 33234 7646 33236 7698
rect 33180 7634 33236 7646
rect 33292 7700 33348 7710
rect 33292 7606 33348 7644
rect 32620 7588 32676 7598
rect 32620 7494 32676 7532
rect 32732 7532 33124 7588
rect 32284 7476 32340 7486
rect 32172 7474 32340 7476
rect 32172 7422 32286 7474
rect 32338 7422 32340 7474
rect 32172 7420 32340 7422
rect 32284 7364 32340 7420
rect 32732 7364 32788 7532
rect 33068 7474 33124 7532
rect 33068 7422 33070 7474
rect 33122 7422 33124 7474
rect 32284 7308 32788 7364
rect 32956 7364 33012 7374
rect 32060 7196 32452 7252
rect 31948 7186 32004 7196
rect 31836 6748 32228 6804
rect 30828 6738 30884 6748
rect 30044 6692 30100 6702
rect 29148 6690 30100 6692
rect 29148 6638 30046 6690
rect 30098 6638 30100 6690
rect 29148 6636 30100 6638
rect 30044 6626 30100 6636
rect 28476 6078 28478 6130
rect 28530 6078 28532 6130
rect 28476 6066 28532 6078
rect 29148 6468 29204 6478
rect 29148 6130 29204 6412
rect 29148 6078 29150 6130
rect 29202 6078 29204 6130
rect 29148 6066 29204 6078
rect 32172 6130 32228 6748
rect 32396 6692 32452 7196
rect 32956 6802 33012 7308
rect 32956 6750 32958 6802
rect 33010 6750 33012 6802
rect 32956 6738 33012 6750
rect 32396 6626 32452 6636
rect 32172 6078 32174 6130
rect 32226 6078 32228 6130
rect 32172 6066 32228 6078
rect 32620 6468 32676 6478
rect 32620 6132 32676 6412
rect 32620 6038 32676 6076
rect 33068 6130 33124 7422
rect 33404 7140 33460 8990
rect 34188 9044 34244 10446
rect 34300 9156 34356 10558
rect 34524 10610 34580 10622
rect 34524 10558 34526 10610
rect 34578 10558 34580 10610
rect 34524 10052 34580 10558
rect 34524 9986 34580 9996
rect 34524 9826 34580 9838
rect 34524 9774 34526 9826
rect 34578 9774 34580 9826
rect 34524 9492 34580 9774
rect 34636 9714 34692 11004
rect 34860 10836 34916 10846
rect 34860 10612 34916 10780
rect 35196 10834 35252 11004
rect 35196 10782 35198 10834
rect 35250 10782 35252 10834
rect 35196 10770 35252 10782
rect 35308 10724 35364 10734
rect 35308 10630 35364 10668
rect 35532 10722 35588 11340
rect 36092 10834 36148 11788
rect 36204 11620 36260 12012
rect 36204 11564 36484 11620
rect 36428 11506 36484 11564
rect 36428 11454 36430 11506
rect 36482 11454 36484 11506
rect 36428 11442 36484 11454
rect 36652 11284 36708 13020
rect 36764 12402 36820 13020
rect 36764 12350 36766 12402
rect 36818 12350 36820 12402
rect 36764 12338 36820 12350
rect 36988 12402 37044 13132
rect 37324 13186 37492 13188
rect 37324 13134 37438 13186
rect 37490 13134 37492 13186
rect 37324 13132 37492 13134
rect 36988 12350 36990 12402
rect 37042 12350 37044 12402
rect 36988 12338 37044 12350
rect 37100 12852 37156 12862
rect 36876 12066 36932 12078
rect 36876 12014 36878 12066
rect 36930 12014 36932 12066
rect 36428 11228 36708 11284
rect 36764 11396 36820 11406
rect 36316 11170 36372 11182
rect 36316 11118 36318 11170
rect 36370 11118 36372 11170
rect 36316 10948 36372 11118
rect 36316 10882 36372 10892
rect 36092 10782 36094 10834
rect 36146 10782 36148 10834
rect 36092 10770 36148 10782
rect 35532 10670 35534 10722
rect 35586 10670 35588 10722
rect 35532 10658 35588 10670
rect 35980 10722 36036 10734
rect 35980 10670 35982 10722
rect 36034 10670 36036 10722
rect 35084 10612 35140 10622
rect 34860 10610 35028 10612
rect 34860 10558 34862 10610
rect 34914 10558 35028 10610
rect 34860 10556 35028 10558
rect 34860 10546 34916 10556
rect 34748 10500 34804 10510
rect 34748 9828 34804 10444
rect 34972 10052 35028 10556
rect 35084 10518 35140 10556
rect 35868 10610 35924 10622
rect 35868 10558 35870 10610
rect 35922 10558 35924 10610
rect 35532 10388 35588 10398
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 34972 9996 35252 10052
rect 34748 9772 35028 9828
rect 34636 9662 34638 9714
rect 34690 9662 34692 9714
rect 34636 9650 34692 9662
rect 34524 9426 34580 9436
rect 34972 9266 35028 9772
rect 34972 9214 34974 9266
rect 35026 9214 35028 9266
rect 34972 9202 35028 9214
rect 35084 9268 35140 9278
rect 35084 9174 35140 9212
rect 35196 9266 35252 9996
rect 35308 9828 35364 9838
rect 35532 9828 35588 10332
rect 35308 9826 35588 9828
rect 35308 9774 35310 9826
rect 35362 9774 35588 9826
rect 35308 9772 35588 9774
rect 35644 9826 35700 9838
rect 35644 9774 35646 9826
rect 35698 9774 35700 9826
rect 35308 9762 35364 9772
rect 35644 9268 35700 9774
rect 35868 9714 35924 10558
rect 35980 9828 36036 10670
rect 35980 9762 36036 9772
rect 36316 10052 36372 10062
rect 35868 9662 35870 9714
rect 35922 9662 35924 9714
rect 35868 9650 35924 9662
rect 35196 9214 35198 9266
rect 35250 9214 35252 9266
rect 35196 9202 35252 9214
rect 35308 9212 35700 9268
rect 34300 9090 34356 9100
rect 34636 9100 34916 9156
rect 34188 8978 34244 8988
rect 34524 8818 34580 8830
rect 34524 8766 34526 8818
rect 34578 8766 34580 8818
rect 34076 8036 34132 8046
rect 34076 7698 34132 7980
rect 34076 7646 34078 7698
rect 34130 7646 34132 7698
rect 33516 7588 33572 7598
rect 33516 7494 33572 7532
rect 34076 7476 34132 7646
rect 34524 7476 34580 8766
rect 34636 7700 34692 9100
rect 34860 9044 34916 9100
rect 35308 9044 35364 9212
rect 34860 8988 35364 9044
rect 35868 9156 35924 9166
rect 35868 9042 35924 9100
rect 35868 8990 35870 9042
rect 35922 8990 35924 9042
rect 34748 8930 34804 8942
rect 34748 8878 34750 8930
rect 34802 8878 34804 8930
rect 34748 8036 34804 8878
rect 35756 8820 35812 8830
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34748 7970 34804 7980
rect 34860 8370 34916 8382
rect 34860 8318 34862 8370
rect 34914 8318 34916 8370
rect 34860 7924 34916 8318
rect 35756 8370 35812 8764
rect 35868 8428 35924 8990
rect 36316 9042 36372 9996
rect 36316 8990 36318 9042
rect 36370 8990 36372 9042
rect 36316 8708 36372 8990
rect 36316 8642 36372 8652
rect 36428 8428 36484 11228
rect 36540 10724 36596 10734
rect 36764 10724 36820 11340
rect 36876 10836 36932 12014
rect 37100 11394 37156 12796
rect 37100 11342 37102 11394
rect 37154 11342 37156 11394
rect 37100 11330 37156 11342
rect 37324 11394 37380 13132
rect 37436 13122 37492 13132
rect 37548 13076 37604 13086
rect 37548 12982 37604 13020
rect 38220 13076 38276 13086
rect 38220 12962 38276 13020
rect 38220 12910 38222 12962
rect 38274 12910 38276 12962
rect 38220 12898 38276 12910
rect 38668 12964 38724 12974
rect 38668 12962 38836 12964
rect 38668 12910 38670 12962
rect 38722 12910 38836 12962
rect 38668 12908 38836 12910
rect 38668 12898 38724 12908
rect 38780 12404 38836 12908
rect 38780 12310 38836 12348
rect 38892 12740 38948 12750
rect 38892 12290 38948 12684
rect 38892 12238 38894 12290
rect 38946 12238 38948 12290
rect 38108 12068 38164 12078
rect 37884 12066 38164 12068
rect 37884 12014 38110 12066
rect 38162 12014 38164 12066
rect 37884 12012 38164 12014
rect 37324 11342 37326 11394
rect 37378 11342 37380 11394
rect 37324 11330 37380 11342
rect 37548 11394 37604 11406
rect 37548 11342 37550 11394
rect 37602 11342 37604 11394
rect 37212 11170 37268 11182
rect 37212 11118 37214 11170
rect 37266 11118 37268 11170
rect 36876 10780 37156 10836
rect 36764 10668 36932 10724
rect 36540 9154 36596 10668
rect 36876 10164 36932 10668
rect 36988 10612 37044 10622
rect 36988 10518 37044 10556
rect 37100 10388 37156 10780
rect 37212 10500 37268 11118
rect 37548 10836 37604 11342
rect 37772 11396 37828 11406
rect 37772 11302 37828 11340
rect 37884 10836 37940 12012
rect 38108 12002 38164 12012
rect 38220 11956 38276 11966
rect 38220 11954 38388 11956
rect 38220 11902 38222 11954
rect 38274 11902 38388 11954
rect 38220 11900 38388 11902
rect 38220 11890 38276 11900
rect 38220 11620 38276 11630
rect 38220 11526 38276 11564
rect 38108 11508 38164 11518
rect 38108 11414 38164 11452
rect 37548 10770 37604 10780
rect 37772 10780 37940 10836
rect 38332 11396 38388 11900
rect 38556 11620 38612 11630
rect 38332 10834 38388 11340
rect 38332 10782 38334 10834
rect 38386 10782 38388 10834
rect 37436 10724 37492 10734
rect 37436 10630 37492 10668
rect 37212 10444 37716 10500
rect 37100 10332 37492 10388
rect 36876 10108 37380 10164
rect 37212 9826 37268 9838
rect 37212 9774 37214 9826
rect 37266 9774 37268 9826
rect 36540 9102 36542 9154
rect 36594 9102 36596 9154
rect 36540 9090 36596 9102
rect 36988 9714 37044 9726
rect 36988 9662 36990 9714
rect 37042 9662 37044 9714
rect 36652 9044 36708 9054
rect 36652 8950 36708 8988
rect 36988 8820 37044 9662
rect 37212 9268 37268 9774
rect 37212 9202 37268 9212
rect 37212 9042 37268 9054
rect 37212 8990 37214 9042
rect 37266 8990 37268 9042
rect 37212 8932 37268 8990
rect 37212 8866 37268 8876
rect 36988 8754 37044 8764
rect 35868 8372 36036 8428
rect 35756 8318 35758 8370
rect 35810 8318 35812 8370
rect 35756 8306 35812 8318
rect 34860 7858 34916 7868
rect 35196 8258 35252 8270
rect 35196 8206 35198 8258
rect 35250 8206 35252 8258
rect 35084 7700 35140 7710
rect 34636 7698 35140 7700
rect 34636 7646 35086 7698
rect 35138 7646 35140 7698
rect 34636 7644 35140 7646
rect 35084 7634 35140 7644
rect 34860 7476 34916 7486
rect 34524 7474 34916 7476
rect 34524 7422 34862 7474
rect 34914 7422 34916 7474
rect 34524 7420 34916 7422
rect 34076 7410 34132 7420
rect 33964 7364 34020 7374
rect 33964 7270 34020 7308
rect 33404 7084 33684 7140
rect 33292 6692 33348 6702
rect 33292 6598 33348 6636
rect 33068 6078 33070 6130
rect 33122 6078 33124 6130
rect 33068 6066 33124 6078
rect 33180 6580 33236 6590
rect 33180 6130 33236 6524
rect 33180 6078 33182 6130
rect 33234 6078 33236 6130
rect 33180 6066 33236 6078
rect 33292 6132 33348 6142
rect 33292 6038 33348 6076
rect 31276 6018 31332 6030
rect 31276 5966 31278 6018
rect 31330 5966 31332 6018
rect 25900 5070 25902 5122
rect 25954 5070 25956 5122
rect 25900 5058 25956 5070
rect 27244 5906 27300 5918
rect 27244 5854 27246 5906
rect 27298 5854 27300 5906
rect 27244 5124 27300 5854
rect 28028 5908 28084 5918
rect 28028 5814 28084 5852
rect 28700 5906 28756 5918
rect 28700 5854 28702 5906
rect 28754 5854 28756 5906
rect 27692 5794 27748 5806
rect 27692 5742 27694 5794
rect 27746 5742 27748 5794
rect 27692 5236 27748 5742
rect 28140 5236 28196 5246
rect 27692 5234 28196 5236
rect 27692 5182 28142 5234
rect 28194 5182 28196 5234
rect 27692 5180 28196 5182
rect 27468 5124 27524 5134
rect 27244 5122 27524 5124
rect 27244 5070 27470 5122
rect 27522 5070 27524 5122
rect 27244 5068 27524 5070
rect 27468 5058 27524 5068
rect 25228 4900 25284 4910
rect 25228 4562 25284 4844
rect 25228 4510 25230 4562
rect 25282 4510 25284 4562
rect 25228 4498 25284 4510
rect 22988 4228 23044 4238
rect 22988 4134 23044 4172
rect 23100 4114 23156 4126
rect 23100 4062 23102 4114
rect 23154 4062 23156 4114
rect 23100 3554 23156 4062
rect 23772 4116 23828 4284
rect 24332 4226 24388 4396
rect 24668 4340 24724 4350
rect 24668 4246 24724 4284
rect 25452 4340 25508 4350
rect 25452 4246 25508 4284
rect 24332 4174 24334 4226
rect 24386 4174 24388 4226
rect 24332 4162 24388 4174
rect 28140 4228 28196 5180
rect 28364 5122 28420 5134
rect 28364 5070 28366 5122
rect 28418 5070 28420 5122
rect 28364 4340 28420 5070
rect 28588 4340 28644 4350
rect 28364 4338 28644 4340
rect 28364 4286 28590 4338
rect 28642 4286 28644 4338
rect 28364 4284 28644 4286
rect 28140 4134 28196 4172
rect 28588 4228 28644 4284
rect 28588 4162 28644 4172
rect 23772 4050 23828 4060
rect 28700 4114 28756 5854
rect 29372 5906 29428 5918
rect 29372 5854 29374 5906
rect 29426 5854 29428 5906
rect 29372 5346 29428 5854
rect 29372 5294 29374 5346
rect 29426 5294 29428 5346
rect 29372 5282 29428 5294
rect 29484 5908 29540 5918
rect 29484 5234 29540 5852
rect 31276 5460 31332 5966
rect 31612 6020 31668 6030
rect 31612 5926 31668 5964
rect 33628 5906 33684 7084
rect 34300 6804 34356 6814
rect 34076 6580 34132 6590
rect 34076 6486 34132 6524
rect 34188 6132 34244 6142
rect 34188 6038 34244 6076
rect 34300 6018 34356 6748
rect 34300 5966 34302 6018
rect 34354 5966 34356 6018
rect 34300 5954 34356 5966
rect 34412 6356 34468 6366
rect 33628 5854 33630 5906
rect 33682 5854 33684 5906
rect 33628 5842 33684 5854
rect 30940 5404 31332 5460
rect 33068 5684 33124 5694
rect 29484 5182 29486 5234
rect 29538 5182 29540 5234
rect 29484 5170 29540 5182
rect 30604 5236 30660 5246
rect 30044 5124 30100 5134
rect 30044 5030 30100 5068
rect 30604 5124 30660 5180
rect 30940 5124 30996 5404
rect 30604 5122 30996 5124
rect 30604 5070 30606 5122
rect 30658 5070 30996 5122
rect 30604 5068 30996 5070
rect 31052 5234 31108 5246
rect 31052 5182 31054 5234
rect 31106 5182 31108 5234
rect 31052 5124 31108 5182
rect 33068 5234 33124 5628
rect 33068 5182 33070 5234
rect 33122 5182 33124 5234
rect 33068 5170 33124 5182
rect 30604 5058 30660 5068
rect 30828 4338 30884 5068
rect 31052 5058 31108 5068
rect 33628 4900 33684 4910
rect 33628 4806 33684 4844
rect 30828 4286 30830 4338
rect 30882 4286 30884 4338
rect 30828 4274 30884 4286
rect 34300 4340 34356 4350
rect 34412 4340 34468 6300
rect 34860 6356 34916 7420
rect 34972 7476 35028 7486
rect 35196 7476 35252 8206
rect 34972 7382 35028 7420
rect 35084 7474 35252 7476
rect 35084 7422 35198 7474
rect 35250 7422 35252 7474
rect 35084 7420 35252 7422
rect 34860 6290 34916 6300
rect 34748 5908 34804 5918
rect 35084 5908 35140 7420
rect 35196 7410 35252 7420
rect 35308 8260 35364 8270
rect 35308 7252 35364 8204
rect 35420 8258 35476 8270
rect 35420 8206 35422 8258
rect 35474 8206 35476 8258
rect 35420 7476 35476 8206
rect 35868 8260 35924 8270
rect 35868 8166 35924 8204
rect 35644 8034 35700 8046
rect 35644 7982 35646 8034
rect 35698 7982 35700 8034
rect 35644 7812 35700 7982
rect 35644 7746 35700 7756
rect 35756 7924 35812 7934
rect 35756 7586 35812 7868
rect 35868 7700 35924 7710
rect 35980 7700 36036 8372
rect 35924 7644 36036 7700
rect 36092 8372 36484 8428
rect 36876 8708 36932 8718
rect 35868 7606 35924 7644
rect 35756 7534 35758 7586
rect 35810 7534 35812 7586
rect 35756 7522 35812 7534
rect 35420 7474 35588 7476
rect 35420 7422 35422 7474
rect 35474 7422 35588 7474
rect 35420 7420 35588 7422
rect 35420 7410 35476 7420
rect 35308 7186 35364 7196
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34748 5906 35140 5908
rect 34748 5854 34750 5906
rect 34802 5854 35140 5906
rect 34748 5852 35140 5854
rect 35196 6692 35252 6702
rect 35196 5906 35252 6636
rect 35532 6132 35588 7420
rect 36092 6468 36148 8372
rect 36876 7474 36932 8652
rect 36876 7422 36878 7474
rect 36930 7422 36932 7474
rect 36876 7410 36932 7422
rect 36428 7252 36484 7262
rect 36204 6804 36260 6814
rect 36204 6710 36260 6748
rect 36092 6402 36148 6412
rect 35532 6066 35588 6076
rect 35196 5854 35198 5906
rect 35250 5854 35252 5906
rect 34748 5684 34804 5852
rect 35196 5842 35252 5854
rect 34748 5618 34804 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35980 5124 36036 5134
rect 35980 5030 36036 5068
rect 36428 5122 36484 7196
rect 36988 6692 37044 6702
rect 36988 6598 37044 6636
rect 36428 5070 36430 5122
rect 36482 5070 36484 5122
rect 36428 5058 36484 5070
rect 37100 6578 37156 6590
rect 37100 6526 37102 6578
rect 37154 6526 37156 6578
rect 37100 5796 37156 6526
rect 37100 5122 37156 5740
rect 37100 5070 37102 5122
rect 37154 5070 37156 5122
rect 37100 5058 37156 5070
rect 37324 4900 37380 10108
rect 37436 10050 37492 10332
rect 37436 9998 37438 10050
rect 37490 9998 37492 10050
rect 37436 9986 37492 9998
rect 37660 10050 37716 10444
rect 37660 9998 37662 10050
rect 37714 9998 37716 10050
rect 37660 9986 37716 9998
rect 37772 9044 37828 10780
rect 38332 10770 38388 10782
rect 38444 11508 38500 11518
rect 38444 10834 38500 11452
rect 38444 10782 38446 10834
rect 38498 10782 38500 10834
rect 38444 10770 38500 10782
rect 37772 8978 37828 8988
rect 37884 10610 37940 10622
rect 37884 10558 37886 10610
rect 37938 10558 37940 10610
rect 37884 9154 37940 10558
rect 38108 10610 38164 10622
rect 38108 10558 38110 10610
rect 38162 10558 38164 10610
rect 38108 10052 38164 10558
rect 38332 10612 38388 10622
rect 38556 10612 38612 11564
rect 38892 11394 38948 12238
rect 38892 11342 38894 11394
rect 38946 11342 38948 11394
rect 38892 11330 38948 11342
rect 38220 10498 38276 10510
rect 38220 10446 38222 10498
rect 38274 10446 38276 10498
rect 38220 10388 38276 10446
rect 38220 10322 38276 10332
rect 37884 9102 37886 9154
rect 37938 9102 37940 9154
rect 37884 8428 37940 9102
rect 37996 9996 38164 10052
rect 37996 8932 38052 9996
rect 38332 9938 38388 10556
rect 38332 9886 38334 9938
rect 38386 9886 38388 9938
rect 38332 9874 38388 9886
rect 38444 10556 38612 10612
rect 38108 9828 38164 9838
rect 38108 9734 38164 9772
rect 38444 9716 38500 10556
rect 38668 9940 38724 9950
rect 38668 9846 38724 9884
rect 38332 9660 38500 9716
rect 38892 9826 38948 9838
rect 38892 9774 38894 9826
rect 38946 9774 38948 9826
rect 38332 9042 38388 9660
rect 38444 9492 38500 9502
rect 38500 9436 38612 9492
rect 38444 9426 38500 9436
rect 38556 9268 38612 9436
rect 38668 9268 38724 9278
rect 38556 9266 38724 9268
rect 38556 9214 38670 9266
rect 38722 9214 38724 9266
rect 38556 9212 38724 9214
rect 38668 9202 38724 9212
rect 38332 8990 38334 9042
rect 38386 8990 38388 9042
rect 38332 8978 38388 8990
rect 38556 9044 38612 9054
rect 38556 8950 38612 8988
rect 38780 9042 38836 9054
rect 38780 8990 38782 9042
rect 38834 8990 38836 9042
rect 37996 8866 38052 8876
rect 38780 8428 38836 8990
rect 37772 8372 37940 8428
rect 38668 8372 38836 8428
rect 38892 8372 38948 9774
rect 37436 7812 37492 7822
rect 37436 7474 37492 7756
rect 37436 7422 37438 7474
rect 37490 7422 37492 7474
rect 37436 7410 37492 7422
rect 37772 6692 37828 8372
rect 38668 8260 38724 8372
rect 38668 8194 38724 8204
rect 38892 8258 38948 8316
rect 38892 8206 38894 8258
rect 38946 8206 38948 8258
rect 38892 8194 38948 8206
rect 39004 9042 39060 9054
rect 39004 8990 39006 9042
rect 39058 8990 39060 9042
rect 39004 7812 39060 8990
rect 39004 7746 39060 7756
rect 37772 6626 37828 6636
rect 38668 6802 38724 6814
rect 38668 6750 38670 6802
rect 38722 6750 38724 6802
rect 37436 6578 37492 6590
rect 37436 6526 37438 6578
rect 37490 6526 37492 6578
rect 37436 6356 37492 6526
rect 37436 6290 37492 6300
rect 37548 6466 37604 6478
rect 37548 6414 37550 6466
rect 37602 6414 37604 6466
rect 37548 5122 37604 6414
rect 37660 6132 37716 6142
rect 37660 6130 38164 6132
rect 37660 6078 37662 6130
rect 37714 6078 38164 6130
rect 37660 6076 38164 6078
rect 37660 6066 37716 6076
rect 37996 5796 38052 5806
rect 37996 5702 38052 5740
rect 37548 5070 37550 5122
rect 37602 5070 37604 5122
rect 37548 5058 37604 5070
rect 37324 4844 37828 4900
rect 37212 4564 37268 4574
rect 37212 4562 37604 4564
rect 37212 4510 37214 4562
rect 37266 4510 37604 4562
rect 37212 4508 37604 4510
rect 37212 4498 37268 4508
rect 34300 4338 34468 4340
rect 34300 4286 34302 4338
rect 34354 4286 34468 4338
rect 34300 4284 34468 4286
rect 34748 4340 34804 4350
rect 34748 4338 35140 4340
rect 34748 4286 34750 4338
rect 34802 4286 35140 4338
rect 34748 4284 35140 4286
rect 34300 4274 34356 4284
rect 34748 4274 34804 4284
rect 29484 4228 29540 4238
rect 29484 4134 29540 4172
rect 29932 4228 29988 4238
rect 29932 4134 29988 4172
rect 30492 4228 30548 4238
rect 30492 4134 30548 4172
rect 28700 4062 28702 4114
rect 28754 4062 28756 4114
rect 28700 4050 28756 4062
rect 35084 3778 35140 4284
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35084 3726 35086 3778
rect 35138 3726 35140 3778
rect 35084 3714 35140 3726
rect 35196 3668 35252 3678
rect 35196 3574 35252 3612
rect 23100 3502 23102 3554
rect 23154 3502 23156 3554
rect 23100 3490 23156 3502
rect 22876 3390 22878 3442
rect 22930 3390 22932 3442
rect 22876 3378 22932 3390
rect 37548 3442 37604 4508
rect 37772 4562 37828 4844
rect 37772 4510 37774 4562
rect 37826 4510 37828 4562
rect 37772 3668 37828 4510
rect 37772 3602 37828 3612
rect 37996 4338 38052 4350
rect 37996 4286 37998 4338
rect 38050 4286 38052 4338
rect 37884 3556 37940 3566
rect 37996 3556 38052 4286
rect 37884 3554 38052 3556
rect 37884 3502 37886 3554
rect 37938 3502 38052 3554
rect 37884 3500 38052 3502
rect 37884 3490 37940 3500
rect 37548 3390 37550 3442
rect 37602 3390 37604 3442
rect 37548 3378 37604 3390
rect 38108 3444 38164 6076
rect 38668 5908 38724 6750
rect 38444 5852 38668 5908
rect 38444 4226 38500 5852
rect 38668 5814 38724 5852
rect 38892 6690 38948 6702
rect 38892 6638 38894 6690
rect 38946 6638 38948 6690
rect 38892 5906 38948 6638
rect 38892 5854 38894 5906
rect 38946 5854 38948 5906
rect 38444 4174 38446 4226
rect 38498 4174 38500 4226
rect 38444 4162 38500 4174
rect 38556 5682 38612 5694
rect 38556 5630 38558 5682
rect 38610 5630 38612 5682
rect 38556 3554 38612 5630
rect 38668 5236 38724 5246
rect 38892 5236 38948 5854
rect 38724 5180 38948 5236
rect 38668 4338 38724 5180
rect 38668 4286 38670 4338
rect 38722 4286 38724 4338
rect 38668 4274 38724 4286
rect 39116 4228 39172 13468
rect 39228 11396 39284 11406
rect 39228 11302 39284 11340
rect 39452 8932 39508 8942
rect 39452 8838 39508 8876
rect 39340 8818 39396 8830
rect 39340 8766 39342 8818
rect 39394 8766 39396 8818
rect 39340 8258 39396 8766
rect 39340 8206 39342 8258
rect 39394 8206 39396 8258
rect 39340 8194 39396 8206
rect 39564 6692 39620 16268
rect 39788 15540 39844 17054
rect 40348 17108 40404 17118
rect 40348 17014 40404 17052
rect 40012 16100 40068 16110
rect 40012 16006 40068 16044
rect 40684 16098 40740 18284
rect 40684 16046 40686 16098
rect 40738 16046 40740 16098
rect 40684 16034 40740 16046
rect 41132 18226 41188 18238
rect 41132 18174 41134 18226
rect 41186 18174 41188 18226
rect 41132 16098 41188 18174
rect 41244 18116 41300 18510
rect 42028 18450 42084 19964
rect 42812 20020 42868 20030
rect 42812 19926 42868 19964
rect 42588 19906 42644 19918
rect 42588 19854 42590 19906
rect 42642 19854 42644 19906
rect 42028 18398 42030 18450
rect 42082 18398 42084 18450
rect 42028 18386 42084 18398
rect 42252 19348 42308 19358
rect 42588 19348 42644 19854
rect 42308 19292 42644 19348
rect 42700 19794 42756 19806
rect 42700 19742 42702 19794
rect 42754 19742 42756 19794
rect 41244 18050 41300 18060
rect 42140 18340 42196 18350
rect 42140 17778 42196 18284
rect 42140 17726 42142 17778
rect 42194 17726 42196 17778
rect 42140 17714 42196 17726
rect 42252 18338 42308 19292
rect 42700 18676 42756 19742
rect 42252 18286 42254 18338
rect 42306 18286 42308 18338
rect 41804 17442 41860 17454
rect 41804 17390 41806 17442
rect 41858 17390 41860 17442
rect 41804 17108 41860 17390
rect 41916 17108 41972 17118
rect 41804 17106 41972 17108
rect 41804 17054 41918 17106
rect 41970 17054 41972 17106
rect 41804 17052 41972 17054
rect 41916 17042 41972 17052
rect 42140 16884 42196 16894
rect 41132 16046 41134 16098
rect 41186 16046 41188 16098
rect 41132 16034 41188 16046
rect 41916 16882 42196 16884
rect 41916 16830 42142 16882
rect 42194 16830 42196 16882
rect 41916 16828 42196 16830
rect 39788 15474 39844 15484
rect 40236 15986 40292 15998
rect 40236 15934 40238 15986
rect 40290 15934 40292 15986
rect 39900 15426 39956 15438
rect 39900 15374 39902 15426
rect 39954 15374 39956 15426
rect 39676 15314 39732 15326
rect 39676 15262 39678 15314
rect 39730 15262 39732 15314
rect 39676 15204 39732 15262
rect 39900 15316 39956 15374
rect 40236 15428 40292 15934
rect 40908 15540 40964 15550
rect 40908 15446 40964 15484
rect 40236 15362 40292 15372
rect 41132 15428 41188 15438
rect 39900 15250 39956 15260
rect 40796 15316 40852 15326
rect 39676 15138 39732 15148
rect 40796 14530 40852 15260
rect 41132 15314 41188 15372
rect 41132 15262 41134 15314
rect 41186 15262 41188 15314
rect 41132 15250 41188 15262
rect 41916 15090 41972 16828
rect 42140 16818 42196 16828
rect 42028 16100 42084 16110
rect 42252 16100 42308 18286
rect 42588 18620 42756 18676
rect 42588 17666 42644 18620
rect 42700 18452 42756 18462
rect 43036 18452 43092 18462
rect 42700 18450 43092 18452
rect 42700 18398 42702 18450
rect 42754 18398 43038 18450
rect 43090 18398 43092 18450
rect 42700 18396 43092 18398
rect 42700 18386 42756 18396
rect 43036 18386 43092 18396
rect 42588 17614 42590 17666
rect 42642 17614 42644 17666
rect 42588 17602 42644 17614
rect 42084 16044 42308 16100
rect 42924 17442 42980 17454
rect 42924 17390 42926 17442
rect 42978 17390 42980 17442
rect 42028 15202 42084 16044
rect 42924 15988 42980 17390
rect 43260 16324 43316 20132
rect 43708 19460 43764 23212
rect 43820 23202 43876 23212
rect 44044 20188 44100 23772
rect 44156 23154 44212 23166
rect 44156 23102 44158 23154
rect 44210 23102 44212 23154
rect 44156 22932 44212 23102
rect 44212 22876 44324 22932
rect 44156 22866 44212 22876
rect 44268 22482 44324 22876
rect 44268 22430 44270 22482
rect 44322 22430 44324 22482
rect 44268 22418 44324 22430
rect 43820 20132 43876 20142
rect 43820 20038 43876 20076
rect 43932 20132 44100 20188
rect 44268 20578 44324 20590
rect 44268 20526 44270 20578
rect 44322 20526 44324 20578
rect 43708 19394 43764 19404
rect 43484 19010 43540 19022
rect 43484 18958 43486 19010
rect 43538 18958 43540 19010
rect 43372 18676 43428 18686
rect 43484 18676 43540 18958
rect 43372 18674 43540 18676
rect 43372 18622 43374 18674
rect 43426 18622 43540 18674
rect 43372 18620 43540 18622
rect 43372 18610 43428 18620
rect 43932 18340 43988 20132
rect 44156 20020 44212 20030
rect 44268 20020 44324 20526
rect 44156 20018 44324 20020
rect 44156 19966 44158 20018
rect 44210 19966 44324 20018
rect 44156 19964 44324 19966
rect 44156 19954 44212 19964
rect 44268 19572 44324 19964
rect 44268 19506 44324 19516
rect 44044 19348 44100 19358
rect 44044 19254 44100 19292
rect 43820 18284 43988 18340
rect 43820 17106 43876 18284
rect 43820 17054 43822 17106
rect 43874 17054 43876 17106
rect 43596 16884 43652 16894
rect 43596 16790 43652 16828
rect 43820 16324 43876 17054
rect 43260 16268 43540 16324
rect 43372 15988 43428 15998
rect 42924 15986 43428 15988
rect 42924 15934 43374 15986
rect 43426 15934 43428 15986
rect 42924 15932 43428 15934
rect 43372 15922 43428 15932
rect 42028 15150 42030 15202
rect 42082 15150 42084 15202
rect 42028 15138 42084 15150
rect 42476 15314 42532 15326
rect 42476 15262 42478 15314
rect 42530 15262 42532 15314
rect 42476 15204 42532 15262
rect 43484 15316 43540 16268
rect 43820 16258 43876 16268
rect 43932 18116 43988 18126
rect 43932 16210 43988 18060
rect 44156 16884 44212 16894
rect 44156 16790 44212 16828
rect 43932 16158 43934 16210
rect 43986 16158 43988 16210
rect 43932 16146 43988 16158
rect 43484 15222 43540 15260
rect 43036 15204 43092 15214
rect 42476 15202 43092 15204
rect 42476 15150 43038 15202
rect 43090 15150 43092 15202
rect 42476 15148 43092 15150
rect 41916 15038 41918 15090
rect 41970 15038 41972 15090
rect 41916 15026 41972 15038
rect 40796 14478 40798 14530
rect 40850 14478 40852 14530
rect 40796 14466 40852 14478
rect 41244 14532 41300 14542
rect 41244 14438 41300 14476
rect 41804 14530 41860 14542
rect 41804 14478 41806 14530
rect 41858 14478 41860 14530
rect 41580 14418 41636 14430
rect 41580 14366 41582 14418
rect 41634 14366 41636 14418
rect 41244 14308 41300 14318
rect 41300 14252 41412 14308
rect 41244 14242 41300 14252
rect 39788 13972 39844 13982
rect 40012 13972 40068 13982
rect 39844 13970 40068 13972
rect 39844 13918 40014 13970
rect 40066 13918 40068 13970
rect 39844 13916 40068 13918
rect 39788 13906 39844 13916
rect 40012 13906 40068 13916
rect 40348 13748 40404 13758
rect 40348 13654 40404 13692
rect 41244 13748 41300 13758
rect 41244 13654 41300 13692
rect 39676 13522 39732 13534
rect 39676 13470 39678 13522
rect 39730 13470 39732 13522
rect 39676 13076 39732 13470
rect 39676 13010 39732 13020
rect 41132 12738 41188 12750
rect 41132 12686 41134 12738
rect 41186 12686 41188 12738
rect 41132 12402 41188 12686
rect 41132 12350 41134 12402
rect 41186 12350 41188 12402
rect 41132 12338 41188 12350
rect 41356 10834 41412 14252
rect 41468 12292 41524 12302
rect 41580 12292 41636 14366
rect 41804 13636 41860 14478
rect 41804 13542 41860 13580
rect 42028 14532 42084 14542
rect 42028 13746 42084 14476
rect 42700 14308 42756 14318
rect 42700 13970 42756 14252
rect 42700 13918 42702 13970
rect 42754 13918 42756 13970
rect 42700 13906 42756 13918
rect 42028 13694 42030 13746
rect 42082 13694 42084 13746
rect 42028 12964 42084 13694
rect 42364 13636 42420 13646
rect 42364 13074 42420 13580
rect 43036 13076 43092 15148
rect 43148 13636 43204 13646
rect 43148 13542 43204 13580
rect 42364 13022 42366 13074
rect 42418 13022 42420 13074
rect 42140 12964 42196 12974
rect 42028 12962 42196 12964
rect 42028 12910 42142 12962
rect 42194 12910 42196 12962
rect 42028 12908 42196 12910
rect 41692 12740 41748 12750
rect 41692 12646 41748 12684
rect 41468 12290 41636 12292
rect 41468 12238 41470 12290
rect 41522 12238 41636 12290
rect 41468 12236 41636 12238
rect 41804 12292 41860 12302
rect 41468 12226 41524 12236
rect 41804 11170 41860 12236
rect 42028 12178 42084 12908
rect 42140 12898 42196 12908
rect 42028 12126 42030 12178
rect 42082 12126 42084 12178
rect 42028 12114 42084 12126
rect 42364 12066 42420 13022
rect 42364 12014 42366 12066
rect 42418 12014 42420 12066
rect 42364 12002 42420 12014
rect 42812 13020 43092 13076
rect 43708 13074 43764 13086
rect 43708 13022 43710 13074
rect 43762 13022 43764 13074
rect 42588 11954 42644 11966
rect 42588 11902 42590 11954
rect 42642 11902 42644 11954
rect 42588 11394 42644 11902
rect 42588 11342 42590 11394
rect 42642 11342 42644 11394
rect 42588 11330 42644 11342
rect 41804 11118 41806 11170
rect 41858 11118 41860 11170
rect 41804 11106 41860 11118
rect 42364 11170 42420 11182
rect 42364 11118 42366 11170
rect 42418 11118 42420 11170
rect 41356 10782 41358 10834
rect 41410 10782 41412 10834
rect 41356 10770 41412 10782
rect 41020 10722 41076 10734
rect 41020 10670 41022 10722
rect 41074 10670 41076 10722
rect 39564 6626 39620 6636
rect 39788 10276 39844 10286
rect 39788 6690 39844 10220
rect 40684 9828 40740 9838
rect 40684 9044 40740 9772
rect 41020 9156 41076 10670
rect 41804 10498 41860 10510
rect 41804 10446 41806 10498
rect 41858 10446 41860 10498
rect 41692 10388 41748 10398
rect 41244 10386 41748 10388
rect 41244 10334 41694 10386
rect 41746 10334 41748 10386
rect 41244 10332 41748 10334
rect 41244 9826 41300 10332
rect 41692 10322 41748 10332
rect 41804 10276 41860 10446
rect 41804 10210 41860 10220
rect 41244 9774 41246 9826
rect 41298 9774 41300 9826
rect 41244 9762 41300 9774
rect 42364 9828 42420 11118
rect 42364 9762 42420 9772
rect 42812 9604 42868 13020
rect 43036 12852 43092 12862
rect 43036 12850 43540 12852
rect 43036 12798 43038 12850
rect 43090 12798 43540 12850
rect 43036 12796 43540 12798
rect 43036 12786 43092 12796
rect 43260 12292 43316 12302
rect 43260 12198 43316 12236
rect 43484 12178 43540 12796
rect 43708 12628 43764 13022
rect 44156 12852 44212 12862
rect 44212 12796 44324 12852
rect 44156 12758 44212 12796
rect 43708 12562 43764 12572
rect 44268 12402 44324 12796
rect 44268 12350 44270 12402
rect 44322 12350 44324 12402
rect 44268 12338 44324 12350
rect 43484 12126 43486 12178
rect 43538 12126 43540 12178
rect 43484 12114 43540 12126
rect 42924 11170 42980 11182
rect 42924 11118 42926 11170
rect 42978 11118 42980 11170
rect 42924 9716 42980 11118
rect 44044 10276 44100 10286
rect 44044 9938 44100 10220
rect 44044 9886 44046 9938
rect 44098 9886 44100 9938
rect 44044 9874 44100 9886
rect 43484 9716 43540 9726
rect 42924 9714 43540 9716
rect 42924 9662 43486 9714
rect 43538 9662 43540 9714
rect 42924 9660 43540 9662
rect 43484 9650 43540 9660
rect 42812 9548 42980 9604
rect 41020 9090 41076 9100
rect 42028 9156 42084 9166
rect 40684 8978 40740 8988
rect 41020 8930 41076 8942
rect 41020 8878 41022 8930
rect 41074 8878 41076 8930
rect 40908 8818 40964 8830
rect 40908 8766 40910 8818
rect 40962 8766 40964 8818
rect 40908 8428 40964 8766
rect 40348 8372 40964 8428
rect 41020 8484 41076 8878
rect 41020 8418 41076 8428
rect 42028 8484 42084 9100
rect 42476 9154 42532 9166
rect 42476 9102 42478 9154
rect 42530 9102 42532 9154
rect 39900 7700 39956 7710
rect 39900 7606 39956 7644
rect 39788 6638 39790 6690
rect 39842 6638 39844 6690
rect 39788 6626 39844 6638
rect 40348 6690 40404 8372
rect 41804 8036 41860 8046
rect 41804 7942 41860 7980
rect 40908 7812 40964 7822
rect 40908 7698 40964 7756
rect 40908 7646 40910 7698
rect 40962 7646 40964 7698
rect 40908 7634 40964 7646
rect 41020 7362 41076 7374
rect 41020 7310 41022 7362
rect 41074 7310 41076 7362
rect 40460 7252 40516 7262
rect 40460 7158 40516 7196
rect 41020 7252 41076 7310
rect 42028 7364 42084 8428
rect 42140 8932 42196 8942
rect 42140 8370 42196 8876
rect 42476 8428 42532 9102
rect 42700 9042 42756 9054
rect 42700 8990 42702 9042
rect 42754 8990 42756 9042
rect 42700 8482 42756 8990
rect 42700 8430 42702 8482
rect 42754 8430 42756 8482
rect 42476 8372 42644 8428
rect 42700 8418 42756 8430
rect 42812 8484 42868 8494
rect 42140 8318 42142 8370
rect 42194 8318 42196 8370
rect 42140 8306 42196 8318
rect 42252 8260 42308 8270
rect 42252 7474 42308 8204
rect 42252 7422 42254 7474
rect 42306 7422 42308 7474
rect 42028 7362 42196 7364
rect 42028 7310 42030 7362
rect 42082 7310 42196 7362
rect 42028 7308 42196 7310
rect 42028 7298 42084 7308
rect 41020 7186 41076 7196
rect 40348 6638 40350 6690
rect 40402 6638 40404 6690
rect 40348 6626 40404 6638
rect 39452 6578 39508 6590
rect 39452 6526 39454 6578
rect 39506 6526 39508 6578
rect 39452 4450 39508 6526
rect 40348 6356 40404 6366
rect 40348 5234 40404 6300
rect 41468 6132 41524 6142
rect 41468 6038 41524 6076
rect 42140 6132 42196 7308
rect 40908 5908 40964 5918
rect 40908 5814 40964 5852
rect 41468 5908 41524 5918
rect 40348 5182 40350 5234
rect 40402 5182 40404 5234
rect 40348 5170 40404 5182
rect 41468 5234 41524 5852
rect 42140 5794 42196 6076
rect 42252 5906 42308 7422
rect 42588 6578 42644 8372
rect 42812 8370 42868 8428
rect 42924 8428 42980 9548
rect 43372 9492 43428 9502
rect 43372 9266 43428 9436
rect 44156 9492 44212 9502
rect 43372 9214 43374 9266
rect 43426 9214 43428 9266
rect 43372 9202 43428 9214
rect 43708 9380 43764 9390
rect 43708 8930 43764 9324
rect 44156 9266 44212 9436
rect 44156 9214 44158 9266
rect 44210 9214 44212 9266
rect 44156 9202 44212 9214
rect 43708 8878 43710 8930
rect 43762 8878 43764 8930
rect 43708 8866 43764 8878
rect 44492 8428 44548 33964
rect 44604 27748 44660 27758
rect 44604 26292 44660 27692
rect 44604 26226 44660 26236
rect 42924 8372 43204 8428
rect 42812 8318 42814 8370
rect 42866 8318 42868 8370
rect 42812 8306 42868 8318
rect 43148 8260 43204 8372
rect 43148 8166 43204 8204
rect 43372 8372 43428 8382
rect 43036 8036 43092 8046
rect 43036 7698 43092 7980
rect 43036 7646 43038 7698
rect 43090 7646 43092 7698
rect 43036 7634 43092 7646
rect 42700 7476 42756 7486
rect 42700 7474 42980 7476
rect 42700 7422 42702 7474
rect 42754 7422 42980 7474
rect 42700 7420 42980 7422
rect 42700 7410 42756 7420
rect 42924 7364 42980 7420
rect 43260 7474 43316 7486
rect 43260 7422 43262 7474
rect 43314 7422 43316 7474
rect 43260 7364 43316 7422
rect 42924 7308 43316 7364
rect 43372 6914 43428 8316
rect 44044 8372 44548 8428
rect 43372 6862 43374 6914
rect 43426 6862 43428 6914
rect 43372 6850 43428 6862
rect 43596 7700 43652 7710
rect 42588 6526 42590 6578
rect 42642 6526 42644 6578
rect 42588 6514 42644 6526
rect 43596 6578 43652 7644
rect 43596 6526 43598 6578
rect 43650 6526 43652 6578
rect 43596 6514 43652 6526
rect 43820 6692 43876 6702
rect 43596 6132 43652 6142
rect 43596 6038 43652 6076
rect 43820 6130 43876 6636
rect 43820 6078 43822 6130
rect 43874 6078 43876 6130
rect 43820 6066 43876 6078
rect 43932 6578 43988 6590
rect 43932 6526 43934 6578
rect 43986 6526 43988 6578
rect 42924 6020 42980 6030
rect 42924 5926 42980 5964
rect 43932 6020 43988 6526
rect 43932 5954 43988 5964
rect 42252 5854 42254 5906
rect 42306 5854 42308 5906
rect 42252 5842 42308 5854
rect 44044 5796 44100 8372
rect 44156 6132 44212 6142
rect 44156 6018 44212 6076
rect 44156 5966 44158 6018
rect 44210 5966 44212 6018
rect 44156 5954 44212 5966
rect 42140 5742 42142 5794
rect 42194 5742 42196 5794
rect 42140 5730 42196 5742
rect 43820 5740 44100 5796
rect 41468 5182 41470 5234
rect 41522 5182 41524 5234
rect 41468 5170 41524 5182
rect 41692 5684 41748 5694
rect 41244 5122 41300 5134
rect 41244 5070 41246 5122
rect 41298 5070 41300 5122
rect 39788 4898 39844 4910
rect 39788 4846 39790 4898
rect 39842 4846 39844 4898
rect 39788 4562 39844 4846
rect 39788 4510 39790 4562
rect 39842 4510 39844 4562
rect 39788 4498 39844 4510
rect 39452 4398 39454 4450
rect 39506 4398 39508 4450
rect 39452 4386 39508 4398
rect 39116 4162 39172 4172
rect 41020 4228 41076 4238
rect 41244 4228 41300 5070
rect 41580 5124 41636 5134
rect 41580 4562 41636 5068
rect 41580 4510 41582 4562
rect 41634 4510 41636 4562
rect 41580 4498 41636 4510
rect 41692 4450 41748 5628
rect 42140 5124 42196 5134
rect 42700 5124 42756 5134
rect 42140 5122 42756 5124
rect 42140 5070 42142 5122
rect 42194 5070 42702 5122
rect 42754 5070 42756 5122
rect 42140 5068 42756 5070
rect 42140 5058 42196 5068
rect 42700 5058 42756 5068
rect 42476 4900 42532 4910
rect 42476 4806 42532 4844
rect 41692 4398 41694 4450
rect 41746 4398 41748 4450
rect 41692 4386 41748 4398
rect 41076 4172 41300 4228
rect 41020 4134 41076 4172
rect 38556 3502 38558 3554
rect 38610 3502 38612 3554
rect 38556 3490 38612 3502
rect 38220 3444 38276 3454
rect 38108 3442 38276 3444
rect 38108 3390 38222 3442
rect 38274 3390 38276 3442
rect 38108 3388 38276 3390
rect 38220 3378 38276 3388
rect 43820 3442 43876 5740
rect 44268 4226 44324 4238
rect 44268 4174 44270 4226
rect 44322 4174 44324 4226
rect 43820 3390 43822 3442
rect 43874 3390 43876 3442
rect 43820 3378 43876 3390
rect 44156 3444 44212 3454
rect 44268 3444 44324 4174
rect 44156 3442 44324 3444
rect 44156 3390 44158 3442
rect 44210 3390 44324 3442
rect 44156 3388 44324 3390
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 44156 2772 44212 3388
rect 44156 2706 44212 2716
<< via2 >>
rect 41916 43036 41972 43092
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 32844 42082 32900 42084
rect 32844 42030 32846 42082
rect 32846 42030 32898 42082
rect 32898 42030 32900 42082
rect 32844 42028 32900 42030
rect 34076 42082 34132 42084
rect 34076 42030 34078 42082
rect 34078 42030 34130 42082
rect 34130 42030 34132 42082
rect 34076 42028 34132 42030
rect 40348 42028 40404 42084
rect 31612 41916 31668 41972
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 29932 41186 29988 41188
rect 29932 41134 29934 41186
rect 29934 41134 29986 41186
rect 29986 41134 29988 41186
rect 29932 41132 29988 41134
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 26908 40460 26964 40516
rect 27244 40460 27300 40516
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 26796 39730 26852 39732
rect 26796 39678 26798 39730
rect 26798 39678 26850 39730
rect 26850 39678 26852 39730
rect 26796 39676 26852 39678
rect 26684 39618 26740 39620
rect 26684 39566 26686 39618
rect 26686 39566 26738 39618
rect 26738 39566 26740 39618
rect 26684 39564 26740 39566
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 29260 40460 29316 40516
rect 28588 40348 28644 40404
rect 27692 40236 27748 40292
rect 28364 39618 28420 39620
rect 28364 39566 28366 39618
rect 28366 39566 28418 39618
rect 28418 39566 28420 39618
rect 28364 39564 28420 39566
rect 29708 40348 29764 40404
rect 31276 41132 31332 41188
rect 29932 39730 29988 39732
rect 29932 39678 29934 39730
rect 29934 39678 29986 39730
rect 29986 39678 29988 39730
rect 29932 39676 29988 39678
rect 30268 40402 30324 40404
rect 30268 40350 30270 40402
rect 30270 40350 30322 40402
rect 30322 40350 30324 40402
rect 30268 40348 30324 40350
rect 30156 40290 30212 40292
rect 30156 40238 30158 40290
rect 30158 40238 30210 40290
rect 30210 40238 30212 40290
rect 30156 40236 30212 40238
rect 30044 39564 30100 39620
rect 30380 39676 30436 39732
rect 28028 39394 28084 39396
rect 28028 39342 28030 39394
rect 28030 39342 28082 39394
rect 28082 39342 28084 39394
rect 28028 39340 28084 39342
rect 29036 39340 29092 39396
rect 27020 38556 27076 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 27916 38108 27972 38164
rect 30156 39228 30212 39284
rect 29820 39004 29876 39060
rect 29708 38892 29764 38948
rect 29036 38668 29092 38724
rect 29484 38780 29540 38836
rect 29260 38162 29316 38164
rect 29260 38110 29262 38162
rect 29262 38110 29314 38162
rect 29314 38110 29316 38162
rect 29260 38108 29316 38110
rect 29820 38668 29876 38724
rect 30044 38780 30100 38836
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 9436 36370 9492 36372
rect 9436 36318 9438 36370
rect 9438 36318 9490 36370
rect 9490 36318 9492 36370
rect 9436 36316 9492 36318
rect 7308 34972 7364 35028
rect 9324 35026 9380 35028
rect 9324 34974 9326 35026
rect 9326 34974 9378 35026
rect 9378 34974 9380 35026
rect 9324 34972 9380 34974
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 6972 33404 7028 33460
rect 7756 33404 7812 33460
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 7308 33234 7364 33236
rect 7308 33182 7310 33234
rect 7310 33182 7362 33234
rect 7362 33182 7364 33234
rect 7308 33180 7364 33182
rect 7980 32620 8036 32676
rect 8876 33404 8932 33460
rect 10444 36316 10500 36372
rect 10780 35698 10836 35700
rect 10780 35646 10782 35698
rect 10782 35646 10834 35698
rect 10834 35646 10836 35698
rect 10780 35644 10836 35646
rect 16156 35810 16212 35812
rect 16156 35758 16158 35810
rect 16158 35758 16210 35810
rect 16210 35758 16212 35810
rect 16156 35756 16212 35758
rect 15820 35196 15876 35252
rect 14588 34860 14644 34916
rect 11452 34300 11508 34356
rect 10108 33180 10164 33236
rect 9548 32674 9604 32676
rect 9548 32622 9550 32674
rect 9550 32622 9602 32674
rect 9602 32622 9604 32674
rect 9548 32620 9604 32622
rect 6076 31836 6132 31892
rect 7980 31890 8036 31892
rect 7980 31838 7982 31890
rect 7982 31838 8034 31890
rect 8034 31838 8036 31890
rect 7980 31836 8036 31838
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 10892 33180 10948 33236
rect 12684 34130 12740 34132
rect 12684 34078 12686 34130
rect 12686 34078 12738 34130
rect 12738 34078 12740 34130
rect 12684 34076 12740 34078
rect 13132 32508 13188 32564
rect 13468 34076 13524 34132
rect 11564 32284 11620 32340
rect 15932 34802 15988 34804
rect 15932 34750 15934 34802
rect 15934 34750 15986 34802
rect 15986 34750 15988 34802
rect 15932 34748 15988 34750
rect 17948 35868 18004 35924
rect 16716 35756 16772 35812
rect 16828 34914 16884 34916
rect 16828 34862 16830 34914
rect 16830 34862 16882 34914
rect 16882 34862 16884 34914
rect 16828 34860 16884 34862
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19404 35868 19460 35924
rect 17500 35196 17556 35252
rect 17388 34748 17444 34804
rect 16492 34076 16548 34132
rect 17276 34130 17332 34132
rect 17276 34078 17278 34130
rect 17278 34078 17330 34130
rect 17330 34078 17332 34130
rect 17276 34076 17332 34078
rect 17388 33292 17444 33348
rect 17724 34076 17780 34132
rect 14924 32674 14980 32676
rect 14924 32622 14926 32674
rect 14926 32622 14978 32674
rect 14978 32622 14980 32674
rect 14924 32620 14980 32622
rect 14588 32562 14644 32564
rect 14588 32510 14590 32562
rect 14590 32510 14642 32562
rect 14642 32510 14644 32562
rect 14588 32508 14644 32510
rect 8876 29426 8932 29428
rect 8876 29374 8878 29426
rect 8878 29374 8930 29426
rect 8930 29374 8932 29426
rect 8876 29372 8932 29374
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 6076 28700 6132 28756
rect 8316 28754 8372 28756
rect 8316 28702 8318 28754
rect 8318 28702 8370 28754
rect 8370 28702 8372 28754
rect 8316 28700 8372 28702
rect 7644 28642 7700 28644
rect 7644 28590 7646 28642
rect 7646 28590 7698 28642
rect 7698 28590 7700 28642
rect 7644 28588 7700 28590
rect 9548 29426 9604 29428
rect 9548 29374 9550 29426
rect 9550 29374 9602 29426
rect 9602 29374 9604 29426
rect 9548 29372 9604 29374
rect 15596 32674 15652 32676
rect 15596 32622 15598 32674
rect 15598 32622 15650 32674
rect 15650 32622 15652 32674
rect 15596 32620 15652 32622
rect 16156 32674 16212 32676
rect 16156 32622 16158 32674
rect 16158 32622 16210 32674
rect 16210 32622 16212 32674
rect 16156 32620 16212 32622
rect 17500 32620 17556 32676
rect 15036 31836 15092 31892
rect 17164 32284 17220 32340
rect 16268 31836 16324 31892
rect 18620 35810 18676 35812
rect 18620 35758 18622 35810
rect 18622 35758 18674 35810
rect 18674 35758 18676 35810
rect 18620 35756 18676 35758
rect 18284 35196 18340 35252
rect 18284 34748 18340 34804
rect 23548 35810 23604 35812
rect 23548 35758 23550 35810
rect 23550 35758 23602 35810
rect 23602 35758 23604 35810
rect 23548 35756 23604 35758
rect 17948 34636 18004 34692
rect 18620 34076 18676 34132
rect 18732 34748 18788 34804
rect 18172 33964 18228 34020
rect 17948 33292 18004 33348
rect 18620 33346 18676 33348
rect 18620 33294 18622 33346
rect 18622 33294 18674 33346
rect 18674 33294 18676 33346
rect 18620 33292 18676 33294
rect 18844 34300 18900 34356
rect 24220 35980 24276 36036
rect 23772 35644 23828 35700
rect 19964 34690 20020 34692
rect 19964 34638 19966 34690
rect 19966 34638 20018 34690
rect 20018 34638 20020 34690
rect 19964 34636 20020 34638
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 17836 31554 17892 31556
rect 17836 31502 17838 31554
rect 17838 31502 17890 31554
rect 17890 31502 17892 31554
rect 17836 31500 17892 31502
rect 18284 31554 18340 31556
rect 18284 31502 18286 31554
rect 18286 31502 18338 31554
rect 18338 31502 18340 31554
rect 18284 31500 18340 31502
rect 16716 30994 16772 30996
rect 16716 30942 16718 30994
rect 16718 30942 16770 30994
rect 16770 30942 16772 30994
rect 16716 30940 16772 30942
rect 18396 30940 18452 30996
rect 15148 30268 15204 30324
rect 11452 29596 11508 29652
rect 13244 29650 13300 29652
rect 13244 29598 13246 29650
rect 13246 29598 13298 29650
rect 13298 29598 13300 29650
rect 13244 29596 13300 29598
rect 10780 29372 10836 29428
rect 8876 28588 8932 28644
rect 13020 29260 13076 29316
rect 15932 30268 15988 30324
rect 13916 29314 13972 29316
rect 13916 29262 13918 29314
rect 13918 29262 13970 29314
rect 13970 29262 13972 29314
rect 13916 29260 13972 29262
rect 17052 30322 17108 30324
rect 17052 30270 17054 30322
rect 17054 30270 17106 30322
rect 17106 30270 17108 30322
rect 17052 30268 17108 30270
rect 17836 30210 17892 30212
rect 17836 30158 17838 30210
rect 17838 30158 17890 30210
rect 17890 30158 17892 30210
rect 17836 30156 17892 30158
rect 16268 29538 16324 29540
rect 16268 29486 16270 29538
rect 16270 29486 16322 29538
rect 16322 29486 16324 29538
rect 16268 29484 16324 29486
rect 17500 29538 17556 29540
rect 17500 29486 17502 29538
rect 17502 29486 17554 29538
rect 17554 29486 17556 29538
rect 17500 29484 17556 29486
rect 16828 29314 16884 29316
rect 16828 29262 16830 29314
rect 16830 29262 16882 29314
rect 16882 29262 16884 29314
rect 16828 29260 16884 29262
rect 14028 28476 14084 28532
rect 16044 28476 16100 28532
rect 11116 27916 11172 27972
rect 10780 27580 10836 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 8540 27244 8596 27300
rect 9212 27244 9268 27300
rect 8988 27132 9044 27188
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 8764 27020 8820 27076
rect 6972 25228 7028 25284
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 7196 24108 7252 24164
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4844 22370 4900 22372
rect 4844 22318 4846 22370
rect 4846 22318 4898 22370
rect 4898 22318 4900 22370
rect 4844 22316 4900 22318
rect 6412 23154 6468 23156
rect 6412 23102 6414 23154
rect 6414 23102 6466 23154
rect 6466 23102 6468 23154
rect 6412 23100 6468 23102
rect 6076 22988 6132 23044
rect 5516 22316 5572 22372
rect 5292 21644 5348 21700
rect 4396 21586 4452 21588
rect 4396 21534 4398 21586
rect 4398 21534 4450 21586
rect 4450 21534 4452 21586
rect 4396 21532 4452 21534
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 2604 19852 2660 19908
rect 6524 22428 6580 22484
rect 6636 21698 6692 21700
rect 6636 21646 6638 21698
rect 6638 21646 6690 21698
rect 6690 21646 6692 21698
rect 6636 21644 6692 21646
rect 4396 20076 4452 20132
rect 5628 20130 5684 20132
rect 5628 20078 5630 20130
rect 5630 20078 5682 20130
rect 5682 20078 5684 20130
rect 5628 20076 5684 20078
rect 4284 19852 4340 19908
rect 4956 19964 5012 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 3276 19234 3332 19236
rect 3276 19182 3278 19234
rect 3278 19182 3330 19234
rect 3330 19182 3332 19234
rect 3276 19180 3332 19182
rect 2044 19068 2100 19124
rect 3164 19122 3220 19124
rect 3164 19070 3166 19122
rect 3166 19070 3218 19122
rect 3218 19070 3220 19122
rect 3164 19068 3220 19070
rect 4620 19068 4676 19124
rect 4844 19180 4900 19236
rect 2380 18674 2436 18676
rect 2380 18622 2382 18674
rect 2382 18622 2434 18674
rect 2434 18622 2436 18674
rect 2380 18620 2436 18622
rect 4956 19292 5012 19348
rect 6076 19292 6132 19348
rect 6524 19346 6580 19348
rect 6524 19294 6526 19346
rect 6526 19294 6578 19346
rect 6578 19294 6580 19346
rect 6524 19292 6580 19294
rect 5068 19234 5124 19236
rect 5068 19182 5070 19234
rect 5070 19182 5122 19234
rect 5122 19182 5124 19234
rect 5068 19180 5124 19182
rect 5964 19234 6020 19236
rect 5964 19182 5966 19234
rect 5966 19182 6018 19234
rect 6018 19182 6020 19234
rect 5964 19180 6020 19182
rect 5628 18620 5684 18676
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 7756 25228 7812 25284
rect 10108 27132 10164 27188
rect 9660 27074 9716 27076
rect 9660 27022 9662 27074
rect 9662 27022 9714 27074
rect 9714 27022 9716 27074
rect 9660 27020 9716 27022
rect 10220 26908 10276 26964
rect 9772 26066 9828 26068
rect 9772 26014 9774 26066
rect 9774 26014 9826 26066
rect 9826 26014 9828 26066
rect 9772 26012 9828 26014
rect 10556 26348 10612 26404
rect 11004 27074 11060 27076
rect 11004 27022 11006 27074
rect 11006 27022 11058 27074
rect 11058 27022 11060 27074
rect 11004 27020 11060 27022
rect 12236 27916 12292 27972
rect 13804 27970 13860 27972
rect 13804 27918 13806 27970
rect 13806 27918 13858 27970
rect 13858 27918 13860 27970
rect 13804 27916 13860 27918
rect 17388 27970 17444 27972
rect 17388 27918 17390 27970
rect 17390 27918 17442 27970
rect 17442 27918 17444 27970
rect 17388 27916 17444 27918
rect 11564 27746 11620 27748
rect 11564 27694 11566 27746
rect 11566 27694 11618 27746
rect 11618 27694 11620 27746
rect 11564 27692 11620 27694
rect 11900 27634 11956 27636
rect 11900 27582 11902 27634
rect 11902 27582 11954 27634
rect 11954 27582 11956 27634
rect 11900 27580 11956 27582
rect 11228 27132 11284 27188
rect 12460 27692 12516 27748
rect 12236 26962 12292 26964
rect 12236 26910 12238 26962
rect 12238 26910 12290 26962
rect 12290 26910 12292 26962
rect 12236 26908 12292 26910
rect 15708 26962 15764 26964
rect 15708 26910 15710 26962
rect 15710 26910 15762 26962
rect 15762 26910 15764 26962
rect 15708 26908 15764 26910
rect 12348 26572 12404 26628
rect 13468 26572 13524 26628
rect 13132 26514 13188 26516
rect 13132 26462 13134 26514
rect 13134 26462 13186 26514
rect 13186 26462 13188 26514
rect 13132 26460 13188 26462
rect 12348 26012 12404 26068
rect 10332 25228 10388 25284
rect 9884 24892 9940 24948
rect 8540 23938 8596 23940
rect 8540 23886 8542 23938
rect 8542 23886 8594 23938
rect 8594 23886 8596 23938
rect 8540 23884 8596 23886
rect 7868 23826 7924 23828
rect 7868 23774 7870 23826
rect 7870 23774 7922 23826
rect 7922 23774 7924 23826
rect 7868 23772 7924 23774
rect 7756 23154 7812 23156
rect 7756 23102 7758 23154
rect 7758 23102 7810 23154
rect 7810 23102 7812 23154
rect 7756 23100 7812 23102
rect 7196 22988 7252 23044
rect 7420 22370 7476 22372
rect 7420 22318 7422 22370
rect 7422 22318 7474 22370
rect 7474 22318 7476 22370
rect 7420 22316 7476 22318
rect 9548 23826 9604 23828
rect 9548 23774 9550 23826
rect 9550 23774 9602 23826
rect 9602 23774 9604 23826
rect 9548 23772 9604 23774
rect 11676 25228 11732 25284
rect 10892 24946 10948 24948
rect 10892 24894 10894 24946
rect 10894 24894 10946 24946
rect 10946 24894 10948 24946
rect 10892 24892 10948 24894
rect 9212 22988 9268 23044
rect 10444 22594 10500 22596
rect 10444 22542 10446 22594
rect 10446 22542 10498 22594
rect 10498 22542 10500 22594
rect 10444 22540 10500 22542
rect 10444 22316 10500 22372
rect 9212 21868 9268 21924
rect 7756 21586 7812 21588
rect 7756 21534 7758 21586
rect 7758 21534 7810 21586
rect 7810 21534 7812 21586
rect 7756 21532 7812 21534
rect 10892 22988 10948 23044
rect 10892 22092 10948 22148
rect 10668 21868 10724 21924
rect 11340 22316 11396 22372
rect 10892 21308 10948 21364
rect 10444 20524 10500 20580
rect 8428 20076 8484 20132
rect 11900 22652 11956 22708
rect 13916 26514 13972 26516
rect 13916 26462 13918 26514
rect 13918 26462 13970 26514
rect 13970 26462 13972 26514
rect 13916 26460 13972 26462
rect 14140 26348 14196 26404
rect 12796 25228 12852 25284
rect 16716 26908 16772 26964
rect 16828 26290 16884 26292
rect 16828 26238 16830 26290
rect 16830 26238 16882 26290
rect 16882 26238 16884 26290
rect 16828 26236 16884 26238
rect 16268 25676 16324 25732
rect 16716 26012 16772 26068
rect 17388 26066 17444 26068
rect 17388 26014 17390 26066
rect 17390 26014 17442 26066
rect 17442 26014 17444 26066
rect 17388 26012 17444 26014
rect 17500 25676 17556 25732
rect 12796 23324 12852 23380
rect 12684 22652 12740 22708
rect 12348 22370 12404 22372
rect 12348 22318 12350 22370
rect 12350 22318 12402 22370
rect 12402 22318 12404 22370
rect 12348 22316 12404 22318
rect 12572 22316 12628 22372
rect 11564 21756 11620 21812
rect 12796 22258 12852 22260
rect 12796 22206 12798 22258
rect 12798 22206 12850 22258
rect 12850 22206 12852 22258
rect 12796 22204 12852 22206
rect 12460 21756 12516 21812
rect 13580 23378 13636 23380
rect 13580 23326 13582 23378
rect 13582 23326 13634 23378
rect 13634 23326 13636 23378
rect 13580 23324 13636 23326
rect 15820 24444 15876 24500
rect 16044 25228 16100 25284
rect 13692 22540 13748 22596
rect 13244 22092 13300 22148
rect 11676 21644 11732 21700
rect 11788 21586 11844 21588
rect 11788 21534 11790 21586
rect 11790 21534 11842 21586
rect 11842 21534 11844 21586
rect 11788 21532 11844 21534
rect 12012 21308 12068 21364
rect 11564 20860 11620 20916
rect 12348 21420 12404 21476
rect 12236 20748 12292 20804
rect 11340 20130 11396 20132
rect 11340 20078 11342 20130
rect 11342 20078 11394 20130
rect 11394 20078 11396 20130
rect 11340 20076 11396 20078
rect 11004 19180 11060 19236
rect 11116 19852 11172 19908
rect 6636 19068 6692 19124
rect 7196 18450 7252 18452
rect 7196 18398 7198 18450
rect 7198 18398 7250 18450
rect 7250 18398 7252 18450
rect 7196 18396 7252 18398
rect 5180 17724 5236 17780
rect 5964 17778 6020 17780
rect 5964 17726 5966 17778
rect 5966 17726 6018 17778
rect 6018 17726 6020 17778
rect 5964 17724 6020 17726
rect 6524 17554 6580 17556
rect 6524 17502 6526 17554
rect 6526 17502 6578 17554
rect 6578 17502 6580 17554
rect 6524 17500 6580 17502
rect 11116 18956 11172 19012
rect 8876 18508 8932 18564
rect 8540 18450 8596 18452
rect 8540 18398 8542 18450
rect 8542 18398 8594 18450
rect 8594 18398 8596 18450
rect 8540 18396 8596 18398
rect 7644 17500 7700 17556
rect 6076 17106 6132 17108
rect 6076 17054 6078 17106
rect 6078 17054 6130 17106
rect 6130 17054 6132 17106
rect 6076 17052 6132 17054
rect 9772 18508 9828 18564
rect 9660 17778 9716 17780
rect 9660 17726 9662 17778
rect 9662 17726 9714 17778
rect 9714 17726 9716 17778
rect 9660 17724 9716 17726
rect 8204 17052 8260 17108
rect 8988 17052 9044 17108
rect 7196 16940 7252 16996
rect 5292 16882 5348 16884
rect 5292 16830 5294 16882
rect 5294 16830 5346 16882
rect 5346 16830 5348 16882
rect 5292 16828 5348 16830
rect 7084 16828 7140 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 8316 16940 8372 16996
rect 9324 16828 9380 16884
rect 8428 15314 8484 15316
rect 8428 15262 8430 15314
rect 8430 15262 8482 15314
rect 8482 15262 8484 15314
rect 8428 15260 8484 15262
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 9548 15986 9604 15988
rect 9548 15934 9550 15986
rect 9550 15934 9602 15986
rect 9602 15934 9604 15986
rect 9548 15932 9604 15934
rect 8764 15820 8820 15876
rect 9436 15874 9492 15876
rect 9436 15822 9438 15874
rect 9438 15822 9490 15874
rect 9490 15822 9492 15874
rect 9436 15820 9492 15822
rect 8988 15426 9044 15428
rect 8988 15374 8990 15426
rect 8990 15374 9042 15426
rect 9042 15374 9044 15426
rect 8988 15372 9044 15374
rect 10668 18562 10724 18564
rect 10668 18510 10670 18562
rect 10670 18510 10722 18562
rect 10722 18510 10724 18562
rect 10668 18508 10724 18510
rect 10892 18450 10948 18452
rect 10892 18398 10894 18450
rect 10894 18398 10946 18450
rect 10946 18398 10948 18450
rect 10892 18396 10948 18398
rect 10556 18338 10612 18340
rect 10556 18286 10558 18338
rect 10558 18286 10610 18338
rect 10610 18286 10612 18338
rect 10556 18284 10612 18286
rect 10332 16716 10388 16772
rect 10444 16604 10500 16660
rect 10668 16716 10724 16772
rect 12460 20860 12516 20916
rect 12572 21084 12628 21140
rect 12684 20130 12740 20132
rect 12684 20078 12686 20130
rect 12686 20078 12738 20130
rect 12738 20078 12740 20130
rect 12684 20076 12740 20078
rect 12012 20018 12068 20020
rect 12012 19966 12014 20018
rect 12014 19966 12066 20018
rect 12066 19966 12068 20018
rect 12012 19964 12068 19966
rect 11900 19234 11956 19236
rect 11900 19182 11902 19234
rect 11902 19182 11954 19234
rect 11954 19182 11956 19234
rect 11900 19180 11956 19182
rect 12124 19122 12180 19124
rect 12124 19070 12126 19122
rect 12126 19070 12178 19122
rect 12178 19070 12180 19122
rect 12124 19068 12180 19070
rect 12348 19010 12404 19012
rect 12348 18958 12350 19010
rect 12350 18958 12402 19010
rect 12402 18958 12404 19010
rect 12348 18956 12404 18958
rect 12460 18396 12516 18452
rect 11900 18338 11956 18340
rect 11900 18286 11902 18338
rect 11902 18286 11954 18338
rect 11954 18286 11956 18338
rect 11900 18284 11956 18286
rect 11676 17778 11732 17780
rect 11676 17726 11678 17778
rect 11678 17726 11730 17778
rect 11730 17726 11732 17778
rect 11676 17724 11732 17726
rect 11900 16940 11956 16996
rect 11340 16604 11396 16660
rect 11788 16828 11844 16884
rect 11228 16210 11284 16212
rect 11228 16158 11230 16210
rect 11230 16158 11282 16210
rect 11282 16158 11284 16210
rect 11228 16156 11284 16158
rect 10556 16044 10612 16100
rect 10220 15932 10276 15988
rect 12572 18620 12628 18676
rect 12908 20636 12964 20692
rect 13692 21756 13748 21812
rect 13468 20690 13524 20692
rect 13468 20638 13470 20690
rect 13470 20638 13522 20690
rect 13522 20638 13524 20690
rect 13468 20636 13524 20638
rect 13916 21532 13972 21588
rect 13804 21084 13860 21140
rect 14588 22988 14644 23044
rect 14476 21698 14532 21700
rect 14476 21646 14478 21698
rect 14478 21646 14530 21698
rect 14530 21646 14532 21698
rect 14476 21644 14532 21646
rect 14140 21308 14196 21364
rect 14028 20748 14084 20804
rect 14364 21474 14420 21476
rect 14364 21422 14366 21474
rect 14366 21422 14418 21474
rect 14418 21422 14420 21474
rect 14364 21420 14420 21422
rect 13916 20076 13972 20132
rect 14252 20524 14308 20580
rect 13580 19852 13636 19908
rect 13804 19740 13860 19796
rect 13132 19516 13188 19572
rect 15260 22204 15316 22260
rect 15820 22204 15876 22260
rect 15484 21810 15540 21812
rect 15484 21758 15486 21810
rect 15486 21758 15538 21810
rect 15538 21758 15540 21810
rect 15484 21756 15540 21758
rect 14700 21644 14756 21700
rect 16492 21756 16548 21812
rect 15932 21698 15988 21700
rect 15932 21646 15934 21698
rect 15934 21646 15986 21698
rect 15986 21646 15988 21698
rect 15932 21644 15988 21646
rect 16380 21586 16436 21588
rect 16380 21534 16382 21586
rect 16382 21534 16434 21586
rect 16434 21534 16436 21586
rect 16380 21532 16436 21534
rect 16716 21474 16772 21476
rect 16716 21422 16718 21474
rect 16718 21422 16770 21474
rect 16770 21422 16772 21474
rect 16716 21420 16772 21422
rect 17276 21308 17332 21364
rect 17500 21420 17556 21476
rect 14476 20242 14532 20244
rect 14476 20190 14478 20242
rect 14478 20190 14530 20242
rect 14530 20190 14532 20242
rect 14476 20188 14532 20190
rect 14588 20018 14644 20020
rect 14588 19966 14590 20018
rect 14590 19966 14642 20018
rect 14642 19966 14644 20018
rect 14588 19964 14644 19966
rect 14140 19852 14196 19908
rect 14700 19628 14756 19684
rect 14140 19068 14196 19124
rect 15372 20188 15428 20244
rect 18284 29538 18340 29540
rect 18284 29486 18286 29538
rect 18286 29486 18338 29538
rect 18338 29486 18340 29538
rect 18284 29484 18340 29486
rect 17836 29426 17892 29428
rect 17836 29374 17838 29426
rect 17838 29374 17890 29426
rect 17890 29374 17892 29426
rect 17836 29372 17892 29374
rect 20412 34802 20468 34804
rect 20412 34750 20414 34802
rect 20414 34750 20466 34802
rect 20466 34750 20468 34802
rect 20412 34748 20468 34750
rect 20972 34636 21028 34692
rect 21084 35420 21140 35476
rect 23100 35420 23156 35476
rect 21084 34300 21140 34356
rect 22092 34300 22148 34356
rect 21980 34130 22036 34132
rect 21980 34078 21982 34130
rect 21982 34078 22034 34130
rect 22034 34078 22036 34130
rect 21980 34076 22036 34078
rect 20524 33292 20580 33348
rect 18620 30716 18676 30772
rect 18396 29372 18452 29428
rect 19180 29260 19236 29316
rect 19180 27858 19236 27860
rect 19180 27806 19182 27858
rect 19182 27806 19234 27858
rect 19234 27806 19236 27858
rect 19180 27804 19236 27806
rect 18284 26908 18340 26964
rect 18956 26962 19012 26964
rect 18956 26910 18958 26962
rect 18958 26910 19010 26962
rect 19010 26910 19012 26962
rect 18956 26908 19012 26910
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20860 32450 20916 32452
rect 20860 32398 20862 32450
rect 20862 32398 20914 32450
rect 20914 32398 20916 32450
rect 20860 32396 20916 32398
rect 24668 35868 24724 35924
rect 24444 35698 24500 35700
rect 24444 35646 24446 35698
rect 24446 35646 24498 35698
rect 24498 35646 24500 35698
rect 24444 35644 24500 35646
rect 24332 35586 24388 35588
rect 24332 35534 24334 35586
rect 24334 35534 24386 35586
rect 24386 35534 24388 35586
rect 24332 35532 24388 35534
rect 24444 35196 24500 35252
rect 24108 34188 24164 34244
rect 24220 33292 24276 33348
rect 22204 33180 22260 33236
rect 19852 30994 19908 30996
rect 19852 30942 19854 30994
rect 19854 30942 19906 30994
rect 19906 30942 19908 30994
rect 19852 30940 19908 30942
rect 20748 30940 20804 30996
rect 20412 30770 20468 30772
rect 20412 30718 20414 30770
rect 20414 30718 20466 30770
rect 20466 30718 20468 30770
rect 20412 30716 20468 30718
rect 21420 30882 21476 30884
rect 21420 30830 21422 30882
rect 21422 30830 21474 30882
rect 21474 30830 21476 30882
rect 21420 30828 21476 30830
rect 24556 34748 24612 34804
rect 26012 36204 26068 36260
rect 25452 35698 25508 35700
rect 25452 35646 25454 35698
rect 25454 35646 25506 35698
rect 25506 35646 25508 35698
rect 25452 35644 25508 35646
rect 26124 35980 26180 36036
rect 26236 36316 26292 36372
rect 25228 35420 25284 35476
rect 24892 35196 24948 35252
rect 26460 36482 26516 36484
rect 26460 36430 26462 36482
rect 26462 36430 26514 36482
rect 26514 36430 26516 36482
rect 26460 36428 26516 36430
rect 30380 39058 30436 39060
rect 30380 39006 30382 39058
rect 30382 39006 30434 39058
rect 30434 39006 30436 39058
rect 30380 39004 30436 39006
rect 30492 38946 30548 38948
rect 30492 38894 30494 38946
rect 30494 38894 30546 38946
rect 30546 38894 30548 38946
rect 30492 38892 30548 38894
rect 30268 38556 30324 38612
rect 30604 38834 30660 38836
rect 30604 38782 30606 38834
rect 30606 38782 30658 38834
rect 30658 38782 30660 38834
rect 30604 38780 30660 38782
rect 31276 40348 31332 40404
rect 32508 41244 32564 41300
rect 31612 40460 31668 40516
rect 31836 39564 31892 39620
rect 31276 39228 31332 39284
rect 32060 39730 32116 39732
rect 32060 39678 32062 39730
rect 32062 39678 32114 39730
rect 32114 39678 32116 39730
rect 32060 39676 32116 39678
rect 30828 38108 30884 38164
rect 32508 39618 32564 39620
rect 32508 39566 32510 39618
rect 32510 39566 32562 39618
rect 32562 39566 32564 39618
rect 32508 39564 32564 39566
rect 32620 38780 32676 38836
rect 31612 38722 31668 38724
rect 31612 38670 31614 38722
rect 31614 38670 31666 38722
rect 31666 38670 31668 38722
rect 31612 38668 31668 38670
rect 32284 38722 32340 38724
rect 32284 38670 32286 38722
rect 32286 38670 32338 38722
rect 32338 38670 32340 38722
rect 32284 38668 32340 38670
rect 26908 35868 26964 35924
rect 26460 35756 26516 35812
rect 26236 35420 26292 35476
rect 26348 35644 26404 35700
rect 26124 35026 26180 35028
rect 26124 34974 26126 35026
rect 26126 34974 26178 35026
rect 26178 34974 26180 35026
rect 26124 34972 26180 34974
rect 24780 34130 24836 34132
rect 24780 34078 24782 34130
rect 24782 34078 24834 34130
rect 24834 34078 24836 34130
rect 24780 34076 24836 34078
rect 25340 33516 25396 33572
rect 25004 33122 25060 33124
rect 25004 33070 25006 33122
rect 25006 33070 25058 33122
rect 25058 33070 25060 33122
rect 25004 33068 25060 33070
rect 24668 32956 24724 33012
rect 24668 32786 24724 32788
rect 24668 32734 24670 32786
rect 24670 32734 24722 32786
rect 24722 32734 24724 32786
rect 24668 32732 24724 32734
rect 24332 32674 24388 32676
rect 24332 32622 24334 32674
rect 24334 32622 24386 32674
rect 24386 32622 24388 32674
rect 24332 32620 24388 32622
rect 22988 32508 23044 32564
rect 25788 34242 25844 34244
rect 25788 34190 25790 34242
rect 25790 34190 25842 34242
rect 25842 34190 25844 34242
rect 25788 34188 25844 34190
rect 25564 33964 25620 34020
rect 26236 34690 26292 34692
rect 26236 34638 26238 34690
rect 26238 34638 26290 34690
rect 26290 34638 26292 34690
rect 26236 34636 26292 34638
rect 25788 33516 25844 33572
rect 25676 33068 25732 33124
rect 25788 33346 25844 33348
rect 25788 33294 25790 33346
rect 25790 33294 25842 33346
rect 25842 33294 25844 33346
rect 25788 33292 25844 33294
rect 25564 32732 25620 32788
rect 25900 33234 25956 33236
rect 25900 33182 25902 33234
rect 25902 33182 25954 33234
rect 25954 33182 25956 33234
rect 25900 33180 25956 33182
rect 27132 36482 27188 36484
rect 27132 36430 27134 36482
rect 27134 36430 27186 36482
rect 27186 36430 27188 36482
rect 27132 36428 27188 36430
rect 27468 36370 27524 36372
rect 27468 36318 27470 36370
rect 27470 36318 27522 36370
rect 27522 36318 27524 36370
rect 27468 36316 27524 36318
rect 27356 35980 27412 36036
rect 27916 36258 27972 36260
rect 27916 36206 27918 36258
rect 27918 36206 27970 36258
rect 27970 36206 27972 36258
rect 27916 36204 27972 36206
rect 30380 35756 30436 35812
rect 27804 35196 27860 35252
rect 26460 34802 26516 34804
rect 26460 34750 26462 34802
rect 26462 34750 26514 34802
rect 26514 34750 26516 34802
rect 26460 34748 26516 34750
rect 26460 34354 26516 34356
rect 26460 34302 26462 34354
rect 26462 34302 26514 34354
rect 26514 34302 26516 34354
rect 26460 34300 26516 34302
rect 26236 33180 26292 33236
rect 25340 32508 25396 32564
rect 22204 30828 22260 30884
rect 22764 30828 22820 30884
rect 20972 30156 21028 30212
rect 21644 30098 21700 30100
rect 21644 30046 21646 30098
rect 21646 30046 21698 30098
rect 21698 30046 21700 30098
rect 21644 30044 21700 30046
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 18732 26236 18788 26292
rect 18620 25340 18676 25396
rect 17948 24834 18004 24836
rect 17948 24782 17950 24834
rect 17950 24782 18002 24834
rect 18002 24782 18004 24834
rect 17948 24780 18004 24782
rect 18060 24722 18116 24724
rect 18060 24670 18062 24722
rect 18062 24670 18114 24722
rect 18114 24670 18116 24722
rect 18060 24668 18116 24670
rect 18284 24444 18340 24500
rect 18508 24108 18564 24164
rect 17836 22988 17892 23044
rect 18508 22428 18564 22484
rect 17724 21698 17780 21700
rect 17724 21646 17726 21698
rect 17726 21646 17778 21698
rect 17778 21646 17780 21698
rect 17724 21644 17780 21646
rect 17948 20972 18004 21028
rect 19292 25340 19348 25396
rect 19068 24780 19124 24836
rect 18844 24722 18900 24724
rect 18844 24670 18846 24722
rect 18846 24670 18898 24722
rect 18898 24670 18900 24722
rect 18844 24668 18900 24670
rect 19180 24444 19236 24500
rect 21308 29372 21364 29428
rect 20636 28642 20692 28644
rect 20636 28590 20638 28642
rect 20638 28590 20690 28642
rect 20690 28590 20692 28642
rect 20636 28588 20692 28590
rect 27244 34636 27300 34692
rect 26796 34018 26852 34020
rect 26796 33966 26798 34018
rect 26798 33966 26850 34018
rect 26850 33966 26852 34018
rect 26796 33964 26852 33966
rect 27132 33068 27188 33124
rect 26796 32732 26852 32788
rect 26684 32620 26740 32676
rect 26012 32450 26068 32452
rect 26012 32398 26014 32450
rect 26014 32398 26066 32450
rect 26066 32398 26068 32450
rect 26012 32396 26068 32398
rect 25900 31612 25956 31668
rect 26908 32956 26964 33012
rect 27020 32562 27076 32564
rect 27020 32510 27022 32562
rect 27022 32510 27074 32562
rect 27074 32510 27076 32562
rect 27020 32508 27076 32510
rect 27468 34188 27524 34244
rect 27692 34860 27748 34916
rect 28140 34802 28196 34804
rect 28140 34750 28142 34802
rect 28142 34750 28194 34802
rect 28194 34750 28196 34802
rect 28140 34748 28196 34750
rect 28700 35586 28756 35588
rect 28700 35534 28702 35586
rect 28702 35534 28754 35586
rect 28754 35534 28756 35586
rect 28700 35532 28756 35534
rect 28364 34636 28420 34692
rect 28700 34748 28756 34804
rect 28588 34300 28644 34356
rect 28252 34130 28308 34132
rect 28252 34078 28254 34130
rect 28254 34078 28306 34130
rect 28306 34078 28308 34130
rect 28252 34076 28308 34078
rect 28028 33628 28084 33684
rect 28700 32620 28756 32676
rect 29708 34972 29764 35028
rect 29372 34860 29428 34916
rect 29148 34300 29204 34356
rect 28924 34130 28980 34132
rect 28924 34078 28926 34130
rect 28926 34078 28978 34130
rect 28978 34078 28980 34130
rect 28924 34076 28980 34078
rect 29036 32674 29092 32676
rect 29036 32622 29038 32674
rect 29038 32622 29090 32674
rect 29090 32622 29092 32674
rect 29036 32620 29092 32622
rect 27916 32450 27972 32452
rect 27916 32398 27918 32450
rect 27918 32398 27970 32450
rect 27970 32398 27972 32450
rect 27916 32396 27972 32398
rect 29932 34802 29988 34804
rect 29932 34750 29934 34802
rect 29934 34750 29986 34802
rect 29986 34750 29988 34802
rect 29932 34748 29988 34750
rect 30156 33234 30212 33236
rect 30156 33182 30158 33234
rect 30158 33182 30210 33234
rect 30210 33182 30212 33234
rect 30156 33180 30212 33182
rect 26236 31500 26292 31556
rect 24556 29596 24612 29652
rect 24780 29708 24836 29764
rect 21308 28588 21364 28644
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20188 27804 20244 27860
rect 20300 27692 20356 27748
rect 20412 26796 20468 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19628 26236 19684 26292
rect 19852 26178 19908 26180
rect 19852 26126 19854 26178
rect 19854 26126 19906 26178
rect 19906 26126 19908 26178
rect 19852 26124 19908 26126
rect 19740 25730 19796 25732
rect 19740 25678 19742 25730
rect 19742 25678 19794 25730
rect 19794 25678 19796 25730
rect 19740 25676 19796 25678
rect 20860 27692 20916 27748
rect 21980 27746 22036 27748
rect 21980 27694 21982 27746
rect 21982 27694 22034 27746
rect 22034 27694 22036 27746
rect 21980 27692 22036 27694
rect 21308 26796 21364 26852
rect 21308 26290 21364 26292
rect 21308 26238 21310 26290
rect 21310 26238 21362 26290
rect 21362 26238 21364 26290
rect 21308 26236 21364 26238
rect 20412 26124 20468 26180
rect 22540 26348 22596 26404
rect 23548 26402 23604 26404
rect 23548 26350 23550 26402
rect 23550 26350 23602 26402
rect 23602 26350 23604 26402
rect 23548 26348 23604 26350
rect 21420 25618 21476 25620
rect 21420 25566 21422 25618
rect 21422 25566 21474 25618
rect 21474 25566 21476 25618
rect 21420 25564 21476 25566
rect 22428 25618 22484 25620
rect 22428 25566 22430 25618
rect 22430 25566 22482 25618
rect 22482 25566 22484 25618
rect 22428 25564 22484 25566
rect 19964 25394 20020 25396
rect 19964 25342 19966 25394
rect 19966 25342 20018 25394
rect 20018 25342 20020 25394
rect 19964 25340 20020 25342
rect 19628 25228 19684 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 24892 20356 24948
rect 21980 24946 22036 24948
rect 21980 24894 21982 24946
rect 21982 24894 22034 24946
rect 22034 24894 22036 24946
rect 21980 24892 22036 24894
rect 22540 24834 22596 24836
rect 22540 24782 22542 24834
rect 22542 24782 22594 24834
rect 22594 24782 22596 24834
rect 22540 24780 22596 24782
rect 24668 29426 24724 29428
rect 24668 29374 24670 29426
rect 24670 29374 24722 29426
rect 24722 29374 24724 29426
rect 24668 29372 24724 29374
rect 25228 29708 25284 29764
rect 26012 31106 26068 31108
rect 26012 31054 26014 31106
rect 26014 31054 26066 31106
rect 26066 31054 26068 31106
rect 26012 31052 26068 31054
rect 25676 29708 25732 29764
rect 25340 29650 25396 29652
rect 25340 29598 25342 29650
rect 25342 29598 25394 29650
rect 25394 29598 25396 29650
rect 25340 29596 25396 29598
rect 26236 29708 26292 29764
rect 26460 29986 26516 29988
rect 26460 29934 26462 29986
rect 26462 29934 26514 29986
rect 26514 29934 26516 29986
rect 26460 29932 26516 29934
rect 26348 29596 26404 29652
rect 29708 31836 29764 31892
rect 27244 31612 27300 31668
rect 27132 31554 27188 31556
rect 27132 31502 27134 31554
rect 27134 31502 27186 31554
rect 27186 31502 27188 31554
rect 27132 31500 27188 31502
rect 27020 31388 27076 31444
rect 27804 31666 27860 31668
rect 27804 31614 27806 31666
rect 27806 31614 27858 31666
rect 27858 31614 27860 31666
rect 27804 31612 27860 31614
rect 27916 31388 27972 31444
rect 26684 29484 26740 29540
rect 27132 29708 27188 29764
rect 25116 28588 25172 28644
rect 23996 27746 24052 27748
rect 23996 27694 23998 27746
rect 23998 27694 24050 27746
rect 24050 27694 24052 27746
rect 23996 27692 24052 27694
rect 24444 27858 24500 27860
rect 24444 27806 24446 27858
rect 24446 27806 24498 27858
rect 24498 27806 24500 27858
rect 24444 27804 24500 27806
rect 23996 26236 24052 26292
rect 23996 25730 24052 25732
rect 23996 25678 23998 25730
rect 23998 25678 24050 25730
rect 24050 25678 24052 25730
rect 23996 25676 24052 25678
rect 25116 25676 25172 25732
rect 23660 24780 23716 24836
rect 24108 24780 24164 24836
rect 19628 24444 19684 24500
rect 18172 21420 18228 21476
rect 17388 20636 17444 20692
rect 15260 19906 15316 19908
rect 15260 19854 15262 19906
rect 15262 19854 15314 19906
rect 15314 19854 15316 19906
rect 15260 19852 15316 19854
rect 14812 19516 14868 19572
rect 14028 18620 14084 18676
rect 17052 19234 17108 19236
rect 17052 19182 17054 19234
rect 17054 19182 17106 19234
rect 17106 19182 17108 19234
rect 17052 19180 17108 19182
rect 18732 21586 18788 21588
rect 18732 21534 18734 21586
rect 18734 21534 18786 21586
rect 18786 21534 18788 21586
rect 18732 21532 18788 21534
rect 18620 21362 18676 21364
rect 18620 21310 18622 21362
rect 18622 21310 18674 21362
rect 18674 21310 18676 21362
rect 18620 21308 18676 21310
rect 19068 23660 19124 23716
rect 22428 24498 22484 24500
rect 22428 24446 22430 24498
rect 22430 24446 22482 24498
rect 22482 24446 22484 24498
rect 22428 24444 22484 24446
rect 23772 24444 23828 24500
rect 19740 24162 19796 24164
rect 19740 24110 19742 24162
rect 19742 24110 19794 24162
rect 19794 24110 19796 24162
rect 19740 24108 19796 24110
rect 19852 23660 19908 23716
rect 20300 23714 20356 23716
rect 20300 23662 20302 23714
rect 20302 23662 20354 23714
rect 20354 23662 20356 23714
rect 20300 23660 20356 23662
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19292 22988 19348 23044
rect 19180 22092 19236 22148
rect 19068 21868 19124 21924
rect 18956 21196 19012 21252
rect 19068 21644 19124 21700
rect 18172 20636 18228 20692
rect 17612 20018 17668 20020
rect 17612 19966 17614 20018
rect 17614 19966 17666 20018
rect 17666 19966 17668 20018
rect 17612 19964 17668 19966
rect 15372 18620 15428 18676
rect 12796 18508 12852 18564
rect 13692 18508 13748 18564
rect 13804 18226 13860 18228
rect 13804 18174 13806 18226
rect 13806 18174 13858 18226
rect 13858 18174 13860 18226
rect 13804 18172 13860 18174
rect 14476 17836 14532 17892
rect 13804 17724 13860 17780
rect 14028 17612 14084 17668
rect 12460 16828 12516 16884
rect 13132 16716 13188 16772
rect 14252 16604 14308 16660
rect 12124 16156 12180 16212
rect 11900 15932 11956 15988
rect 10108 15820 10164 15876
rect 11116 15484 11172 15540
rect 9100 13692 9156 13748
rect 10332 15202 10388 15204
rect 10332 15150 10334 15202
rect 10334 15150 10386 15202
rect 10386 15150 10388 15202
rect 10332 15148 10388 15150
rect 12236 15820 12292 15876
rect 12236 15372 12292 15428
rect 12460 16210 12516 16212
rect 12460 16158 12462 16210
rect 12462 16158 12514 16210
rect 12514 16158 12516 16210
rect 12460 16156 12516 16158
rect 14252 16156 14308 16212
rect 13132 15538 13188 15540
rect 13132 15486 13134 15538
rect 13134 15486 13186 15538
rect 13186 15486 13188 15538
rect 13132 15484 13188 15486
rect 13356 15426 13412 15428
rect 13356 15374 13358 15426
rect 13358 15374 13410 15426
rect 13410 15374 13412 15426
rect 13356 15372 13412 15374
rect 13244 15202 13300 15204
rect 13244 15150 13246 15202
rect 13246 15150 13298 15202
rect 13298 15150 13300 15202
rect 13244 15148 13300 15150
rect 13468 15260 13524 15316
rect 14140 15986 14196 15988
rect 14140 15934 14142 15986
rect 14142 15934 14194 15986
rect 14194 15934 14196 15986
rect 14140 15932 14196 15934
rect 13804 15874 13860 15876
rect 13804 15822 13806 15874
rect 13806 15822 13858 15874
rect 13858 15822 13860 15874
rect 13804 15820 13860 15822
rect 14140 15538 14196 15540
rect 14140 15486 14142 15538
rect 14142 15486 14194 15538
rect 14194 15486 14196 15538
rect 14140 15484 14196 15486
rect 9884 13692 9940 13748
rect 10892 13746 10948 13748
rect 10892 13694 10894 13746
rect 10894 13694 10946 13746
rect 10946 13694 10948 13746
rect 10892 13692 10948 13694
rect 12348 13468 12404 13524
rect 12796 14252 12852 14308
rect 15820 18674 15876 18676
rect 15820 18622 15822 18674
rect 15822 18622 15874 18674
rect 15874 18622 15876 18674
rect 15820 18620 15876 18622
rect 15036 18562 15092 18564
rect 15036 18510 15038 18562
rect 15038 18510 15090 18562
rect 15090 18510 15092 18562
rect 15036 18508 15092 18510
rect 15596 18562 15652 18564
rect 15596 18510 15598 18562
rect 15598 18510 15650 18562
rect 15650 18510 15652 18562
rect 15596 18508 15652 18510
rect 16940 18508 16996 18564
rect 16268 18450 16324 18452
rect 16268 18398 16270 18450
rect 16270 18398 16322 18450
rect 16322 18398 16324 18450
rect 16268 18396 16324 18398
rect 14812 18172 14868 18228
rect 14924 17724 14980 17780
rect 15596 17778 15652 17780
rect 15596 17726 15598 17778
rect 15598 17726 15650 17778
rect 15650 17726 15652 17778
rect 15596 17724 15652 17726
rect 16268 17666 16324 17668
rect 16268 17614 16270 17666
rect 16270 17614 16322 17666
rect 16322 17614 16324 17666
rect 16268 17612 16324 17614
rect 16604 17666 16660 17668
rect 16604 17614 16606 17666
rect 16606 17614 16658 17666
rect 16658 17614 16660 17666
rect 16604 17612 16660 17614
rect 17276 18450 17332 18452
rect 17276 18398 17278 18450
rect 17278 18398 17330 18450
rect 17330 18398 17332 18450
rect 17276 18396 17332 18398
rect 17612 18562 17668 18564
rect 17612 18510 17614 18562
rect 17614 18510 17666 18562
rect 17666 18510 17668 18562
rect 17612 18508 17668 18510
rect 14588 16716 14644 16772
rect 14588 15538 14644 15540
rect 14588 15486 14590 15538
rect 14590 15486 14642 15538
rect 14642 15486 14644 15538
rect 14588 15484 14644 15486
rect 13356 13692 13412 13748
rect 13356 13468 13412 13524
rect 11676 12796 11732 12852
rect 12460 12850 12516 12852
rect 12460 12798 12462 12850
rect 12462 12798 12514 12850
rect 12514 12798 12516 12850
rect 12460 12796 12516 12798
rect 11004 10722 11060 10724
rect 11004 10670 11006 10722
rect 11006 10670 11058 10722
rect 11058 10670 11060 10722
rect 11004 10668 11060 10670
rect 9436 9826 9492 9828
rect 9436 9774 9438 9826
rect 9438 9774 9490 9826
rect 9490 9774 9492 9826
rect 9436 9772 9492 9774
rect 12236 11170 12292 11172
rect 12236 11118 12238 11170
rect 12238 11118 12290 11170
rect 12290 11118 12292 11170
rect 12236 11116 12292 11118
rect 11900 10722 11956 10724
rect 11900 10670 11902 10722
rect 11902 10670 11954 10722
rect 11954 10670 11956 10722
rect 11900 10668 11956 10670
rect 12796 11170 12852 11172
rect 12796 11118 12798 11170
rect 12798 11118 12850 11170
rect 12850 11118 12852 11170
rect 12796 11116 12852 11118
rect 13356 11116 13412 11172
rect 13132 10892 13188 10948
rect 12348 10668 12404 10724
rect 12796 10722 12852 10724
rect 12796 10670 12798 10722
rect 12798 10670 12850 10722
rect 12850 10670 12852 10722
rect 12796 10668 12852 10670
rect 11228 9212 11284 9268
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 9548 8316 9604 8372
rect 11228 8370 11284 8372
rect 11228 8318 11230 8370
rect 11230 8318 11282 8370
rect 11282 8318 11284 8370
rect 11228 8316 11284 8318
rect 11900 8316 11956 8372
rect 11340 8258 11396 8260
rect 11340 8206 11342 8258
rect 11342 8206 11394 8258
rect 11394 8206 11396 8258
rect 11340 8204 11396 8206
rect 12124 8652 12180 8708
rect 12012 8204 12068 8260
rect 12460 9772 12516 9828
rect 13468 9826 13524 9828
rect 13468 9774 13470 9826
rect 13470 9774 13522 9826
rect 13522 9774 13524 9826
rect 13468 9772 13524 9774
rect 13580 13580 13636 13636
rect 12796 9714 12852 9716
rect 12796 9662 12798 9714
rect 12798 9662 12850 9714
rect 12850 9662 12852 9714
rect 12796 9660 12852 9662
rect 13580 9660 13636 9716
rect 13804 13634 13860 13636
rect 13804 13582 13806 13634
rect 13806 13582 13858 13634
rect 13858 13582 13860 13634
rect 13804 13580 13860 13582
rect 12796 9212 12852 9268
rect 10892 8146 10948 8148
rect 10892 8094 10894 8146
rect 10894 8094 10946 8146
rect 10946 8094 10948 8146
rect 10892 8092 10948 8094
rect 9324 7980 9380 8036
rect 10780 8034 10836 8036
rect 10780 7982 10782 8034
rect 10782 7982 10834 8034
rect 10834 7982 10836 8034
rect 10780 7980 10836 7982
rect 13132 9042 13188 9044
rect 13132 8990 13134 9042
rect 13134 8990 13186 9042
rect 13186 8990 13188 9042
rect 13132 8988 13188 8990
rect 13244 8876 13300 8932
rect 13020 8092 13076 8148
rect 14140 13468 14196 13524
rect 14364 13468 14420 13524
rect 14812 15986 14868 15988
rect 14812 15934 14814 15986
rect 14814 15934 14866 15986
rect 14866 15934 14868 15986
rect 14812 15932 14868 15934
rect 16828 16770 16884 16772
rect 16828 16718 16830 16770
rect 16830 16718 16882 16770
rect 16882 16718 16884 16770
rect 16828 16716 16884 16718
rect 16604 16380 16660 16436
rect 15932 16322 15988 16324
rect 15932 16270 15934 16322
rect 15934 16270 15986 16322
rect 15986 16270 15988 16322
rect 15932 16268 15988 16270
rect 15148 16098 15204 16100
rect 15148 16046 15150 16098
rect 15150 16046 15202 16098
rect 15202 16046 15204 16098
rect 15148 16044 15204 16046
rect 17276 16380 17332 16436
rect 17836 17052 17892 17108
rect 17500 16268 17556 16324
rect 16604 15484 16660 15540
rect 17724 15484 17780 15540
rect 14812 14306 14868 14308
rect 14812 14254 14814 14306
rect 14814 14254 14866 14306
rect 14866 14254 14868 14306
rect 14812 14252 14868 14254
rect 15148 13580 15204 13636
rect 15372 13804 15428 13860
rect 15708 14252 15764 14308
rect 15484 13580 15540 13636
rect 15596 13522 15652 13524
rect 15596 13470 15598 13522
rect 15598 13470 15650 13522
rect 15650 13470 15652 13522
rect 15596 13468 15652 13470
rect 15932 14028 15988 14084
rect 16492 13804 16548 13860
rect 17164 14306 17220 14308
rect 17164 14254 17166 14306
rect 17166 14254 17218 14306
rect 17218 14254 17220 14306
rect 17164 14252 17220 14254
rect 18284 20018 18340 20020
rect 18284 19966 18286 20018
rect 18286 19966 18338 20018
rect 18338 19966 18340 20018
rect 18284 19964 18340 19966
rect 18508 18956 18564 19012
rect 18284 18562 18340 18564
rect 18284 18510 18286 18562
rect 18286 18510 18338 18562
rect 18338 18510 18340 18562
rect 18284 18508 18340 18510
rect 18396 17836 18452 17892
rect 18620 18450 18676 18452
rect 18620 18398 18622 18450
rect 18622 18398 18674 18450
rect 18674 18398 18676 18450
rect 18620 18396 18676 18398
rect 18508 15372 18564 15428
rect 19404 21586 19460 21588
rect 19404 21534 19406 21586
rect 19406 21534 19458 21586
rect 19458 21534 19460 21586
rect 19404 21532 19460 21534
rect 19292 21308 19348 21364
rect 19180 20972 19236 21028
rect 19628 21868 19684 21924
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19180 19740 19236 19796
rect 20300 22092 20356 22148
rect 19964 21420 20020 21476
rect 19740 21308 19796 21364
rect 20188 21308 20244 21364
rect 20076 20690 20132 20692
rect 20076 20638 20078 20690
rect 20078 20638 20130 20690
rect 20130 20638 20132 20690
rect 20076 20636 20132 20638
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19628 20076 19684 20132
rect 19964 20188 20020 20244
rect 21196 23266 21252 23268
rect 21196 23214 21198 23266
rect 21198 23214 21250 23266
rect 21250 23214 21252 23266
rect 21196 23212 21252 23214
rect 20524 21308 20580 21364
rect 21532 21532 21588 21588
rect 20412 20188 20468 20244
rect 20636 20130 20692 20132
rect 20636 20078 20638 20130
rect 20638 20078 20690 20130
rect 20690 20078 20692 20130
rect 20636 20076 20692 20078
rect 20300 19740 20356 19796
rect 20188 19180 20244 19236
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19404 18396 19460 18452
rect 19292 18172 19348 18228
rect 18844 17724 18900 17780
rect 19852 17948 19908 18004
rect 18732 17164 18788 17220
rect 18956 17164 19012 17220
rect 19068 17052 19124 17108
rect 19836 17274 19892 17276
rect 19068 16098 19124 16100
rect 19068 16046 19070 16098
rect 19070 16046 19122 16098
rect 19122 16046 19124 16098
rect 19068 16044 19124 16046
rect 19628 17164 19684 17220
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20188 16492 20244 16548
rect 20972 19068 21028 19124
rect 20748 19010 20804 19012
rect 20748 18958 20750 19010
rect 20750 18958 20802 19010
rect 20802 18958 20804 19010
rect 20748 18956 20804 18958
rect 20636 18450 20692 18452
rect 20636 18398 20638 18450
rect 20638 18398 20690 18450
rect 20690 18398 20692 18450
rect 20636 18396 20692 18398
rect 21196 18450 21252 18452
rect 21196 18398 21198 18450
rect 21198 18398 21250 18450
rect 21250 18398 21252 18450
rect 21196 18396 21252 18398
rect 21756 22370 21812 22372
rect 21756 22318 21758 22370
rect 21758 22318 21810 22370
rect 21810 22318 21812 22370
rect 21756 22316 21812 22318
rect 22876 22316 22932 22372
rect 21868 20802 21924 20804
rect 21868 20750 21870 20802
rect 21870 20750 21922 20802
rect 21922 20750 21924 20802
rect 21868 20748 21924 20750
rect 22092 20690 22148 20692
rect 22092 20638 22094 20690
rect 22094 20638 22146 20690
rect 22146 20638 22148 20690
rect 22092 20636 22148 20638
rect 22540 22092 22596 22148
rect 22316 19234 22372 19236
rect 22316 19182 22318 19234
rect 22318 19182 22370 19234
rect 22370 19182 22372 19234
rect 22316 19180 22372 19182
rect 21980 19122 22036 19124
rect 21980 19070 21982 19122
rect 21982 19070 22034 19122
rect 22034 19070 22036 19122
rect 21980 19068 22036 19070
rect 21532 17948 21588 18004
rect 20524 17666 20580 17668
rect 20524 17614 20526 17666
rect 20526 17614 20578 17666
rect 20578 17614 20580 17666
rect 20524 17612 20580 17614
rect 20300 16380 20356 16436
rect 20636 16268 20692 16324
rect 19964 16210 20020 16212
rect 19964 16158 19966 16210
rect 19966 16158 20018 16210
rect 20018 16158 20020 16210
rect 19964 16156 20020 16158
rect 19068 15708 19124 15764
rect 20076 16098 20132 16100
rect 20076 16046 20078 16098
rect 20078 16046 20130 16098
rect 20130 16046 20132 16098
rect 20076 16044 20132 16046
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 18172 14306 18228 14308
rect 18172 14254 18174 14306
rect 18174 14254 18226 14306
rect 18226 14254 18228 14306
rect 18172 14252 18228 14254
rect 17500 13970 17556 13972
rect 17500 13918 17502 13970
rect 17502 13918 17554 13970
rect 17554 13918 17556 13970
rect 17500 13916 17556 13918
rect 18060 13580 18116 13636
rect 18060 13132 18116 13188
rect 16716 12348 16772 12404
rect 17500 12402 17556 12404
rect 17500 12350 17502 12402
rect 17502 12350 17554 12402
rect 17554 12350 17556 12402
rect 17500 12348 17556 12350
rect 16828 12066 16884 12068
rect 16828 12014 16830 12066
rect 16830 12014 16882 12066
rect 16882 12014 16884 12066
rect 16828 12012 16884 12014
rect 17612 12012 17668 12068
rect 15372 10892 15428 10948
rect 15260 10834 15316 10836
rect 15260 10782 15262 10834
rect 15262 10782 15314 10834
rect 15314 10782 15316 10834
rect 15260 10780 15316 10782
rect 13804 10722 13860 10724
rect 13804 10670 13806 10722
rect 13806 10670 13858 10722
rect 13858 10670 13860 10722
rect 13804 10668 13860 10670
rect 15820 11340 15876 11396
rect 15820 10834 15876 10836
rect 15820 10782 15822 10834
rect 15822 10782 15874 10834
rect 15874 10782 15876 10834
rect 15820 10780 15876 10782
rect 16156 9884 16212 9940
rect 14364 9212 14420 9268
rect 13804 8876 13860 8932
rect 14140 8652 14196 8708
rect 15820 9266 15876 9268
rect 15820 9214 15822 9266
rect 15822 9214 15874 9266
rect 15874 9214 15876 9266
rect 15820 9212 15876 9214
rect 17500 9660 17556 9716
rect 15260 9042 15316 9044
rect 15260 8990 15262 9042
rect 15262 8990 15314 9042
rect 15314 8990 15316 9042
rect 15260 8988 15316 8990
rect 15596 8818 15652 8820
rect 15596 8766 15598 8818
rect 15598 8766 15650 8818
rect 15650 8766 15652 8818
rect 15596 8764 15652 8766
rect 14924 8652 14980 8708
rect 13692 8258 13748 8260
rect 13692 8206 13694 8258
rect 13694 8206 13746 8258
rect 13746 8206 13748 8258
rect 13692 8204 13748 8206
rect 13468 8092 13524 8148
rect 12124 8034 12180 8036
rect 12124 7982 12126 8034
rect 12126 7982 12178 8034
rect 12178 7982 12180 8034
rect 12124 7980 12180 7982
rect 12348 7980 12404 8036
rect 11228 6636 11284 6692
rect 12124 6860 12180 6916
rect 11788 6466 11844 6468
rect 11788 6414 11790 6466
rect 11790 6414 11842 6466
rect 11842 6414 11844 6466
rect 11788 6412 11844 6414
rect 8876 6076 8932 6132
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 12684 6748 12740 6804
rect 12572 6690 12628 6692
rect 12572 6638 12574 6690
rect 12574 6638 12626 6690
rect 12626 6638 12628 6690
rect 12572 6636 12628 6638
rect 12236 6412 12292 6468
rect 13132 6130 13188 6132
rect 13132 6078 13134 6130
rect 13134 6078 13186 6130
rect 13186 6078 13188 6130
rect 13132 6076 13188 6078
rect 12460 5628 12516 5684
rect 13468 6748 13524 6804
rect 14028 6748 14084 6804
rect 13916 6412 13972 6468
rect 13356 5628 13412 5684
rect 15820 8146 15876 8148
rect 15820 8094 15822 8146
rect 15822 8094 15874 8146
rect 15874 8094 15876 8146
rect 15820 8092 15876 8094
rect 16044 8876 16100 8932
rect 17052 8092 17108 8148
rect 15932 7756 15988 7812
rect 17388 7980 17444 8036
rect 16828 7474 16884 7476
rect 16828 7422 16830 7474
rect 16830 7422 16882 7474
rect 16882 7422 16884 7474
rect 16828 7420 16884 7422
rect 16716 7362 16772 7364
rect 16716 7310 16718 7362
rect 16718 7310 16770 7362
rect 16770 7310 16772 7362
rect 16716 7308 16772 7310
rect 16716 6860 16772 6916
rect 14364 5964 14420 6020
rect 12572 5234 12628 5236
rect 12572 5182 12574 5234
rect 12574 5182 12626 5234
rect 12626 5182 12628 5234
rect 12572 5180 12628 5182
rect 14252 5234 14308 5236
rect 14252 5182 14254 5234
rect 14254 5182 14306 5234
rect 14306 5182 14308 5234
rect 14252 5180 14308 5182
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 15148 5628 15204 5684
rect 14924 5180 14980 5236
rect 16492 6466 16548 6468
rect 16492 6414 16494 6466
rect 16494 6414 16546 6466
rect 16546 6414 16548 6466
rect 16492 6412 16548 6414
rect 15708 5180 15764 5236
rect 16380 5122 16436 5124
rect 16380 5070 16382 5122
rect 16382 5070 16434 5122
rect 16434 5070 16436 5122
rect 16380 5068 16436 5070
rect 16380 4732 16436 4788
rect 18844 14700 18900 14756
rect 19068 14588 19124 14644
rect 18508 12684 18564 12740
rect 18620 14306 18676 14308
rect 18620 14254 18622 14306
rect 18622 14254 18674 14306
rect 18674 14254 18676 14306
rect 18620 14252 18676 14254
rect 18396 12290 18452 12292
rect 18396 12238 18398 12290
rect 18398 12238 18450 12290
rect 18450 12238 18452 12290
rect 18396 12236 18452 12238
rect 18844 14306 18900 14308
rect 18844 14254 18846 14306
rect 18846 14254 18898 14306
rect 18898 14254 18900 14306
rect 18844 14252 18900 14254
rect 19404 15372 19460 15428
rect 18956 13692 19012 13748
rect 19292 13692 19348 13748
rect 19516 15260 19572 15316
rect 19628 15148 19684 15204
rect 19516 14700 19572 14756
rect 19404 13186 19460 13188
rect 19404 13134 19406 13186
rect 19406 13134 19458 13186
rect 19458 13134 19460 13186
rect 19404 13132 19460 13134
rect 19180 13020 19236 13076
rect 19068 11564 19124 11620
rect 18732 10108 18788 10164
rect 18396 9714 18452 9716
rect 18396 9662 18398 9714
rect 18398 9662 18450 9714
rect 18450 9662 18452 9714
rect 18396 9660 18452 9662
rect 18844 9938 18900 9940
rect 18844 9886 18846 9938
rect 18846 9886 18898 9938
rect 18898 9886 18900 9938
rect 18844 9884 18900 9886
rect 18620 9660 18676 9716
rect 17612 7868 17668 7924
rect 18732 8316 18788 8372
rect 19068 8876 19124 8932
rect 18956 8764 19012 8820
rect 18620 8034 18676 8036
rect 18620 7982 18622 8034
rect 18622 7982 18674 8034
rect 18674 7982 18676 8034
rect 18620 7980 18676 7982
rect 18508 7868 18564 7924
rect 19068 7532 19124 7588
rect 20076 14588 20132 14644
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20524 15874 20580 15876
rect 20524 15822 20526 15874
rect 20526 15822 20578 15874
rect 20578 15822 20580 15874
rect 20524 15820 20580 15822
rect 20860 15372 20916 15428
rect 20636 15148 20692 15204
rect 21196 17612 21252 17668
rect 21308 17554 21364 17556
rect 21308 17502 21310 17554
rect 21310 17502 21362 17554
rect 21362 17502 21364 17554
rect 21308 17500 21364 17502
rect 21308 16156 21364 16212
rect 21644 16940 21700 16996
rect 22428 18172 22484 18228
rect 22204 17554 22260 17556
rect 22204 17502 22206 17554
rect 22206 17502 22258 17554
rect 22258 17502 22260 17554
rect 22204 17500 22260 17502
rect 21756 16492 21812 16548
rect 21980 16492 22036 16548
rect 21868 16098 21924 16100
rect 21868 16046 21870 16098
rect 21870 16046 21922 16098
rect 21922 16046 21924 16098
rect 21868 16044 21924 16046
rect 21420 15372 21476 15428
rect 21532 15932 21588 15988
rect 22316 16770 22372 16772
rect 22316 16718 22318 16770
rect 22318 16718 22370 16770
rect 22370 16718 22372 16770
rect 22316 16716 22372 16718
rect 23996 23100 24052 23156
rect 25564 28642 25620 28644
rect 25564 28590 25566 28642
rect 25566 28590 25618 28642
rect 25618 28590 25620 28642
rect 25564 28588 25620 28590
rect 26012 28082 26068 28084
rect 26012 28030 26014 28082
rect 26014 28030 26066 28082
rect 26066 28030 26068 28082
rect 26012 28028 26068 28030
rect 25900 27970 25956 27972
rect 25900 27918 25902 27970
rect 25902 27918 25954 27970
rect 25954 27918 25956 27970
rect 25900 27916 25956 27918
rect 26012 26908 26068 26964
rect 26236 27244 26292 27300
rect 27020 29426 27076 29428
rect 27020 29374 27022 29426
rect 27022 29374 27074 29426
rect 27074 29374 27076 29426
rect 27020 29372 27076 29374
rect 26908 28588 26964 28644
rect 26572 27858 26628 27860
rect 26572 27806 26574 27858
rect 26574 27806 26626 27858
rect 26626 27806 26628 27858
rect 26572 27804 26628 27806
rect 26572 27020 26628 27076
rect 27020 26962 27076 26964
rect 27020 26910 27022 26962
rect 27022 26910 27074 26962
rect 27074 26910 27076 26962
rect 27020 26908 27076 26910
rect 27468 30044 27524 30100
rect 29932 30940 29988 30996
rect 29596 30156 29652 30212
rect 27804 29986 27860 29988
rect 27804 29934 27806 29986
rect 27806 29934 27858 29986
rect 27858 29934 27860 29986
rect 27804 29932 27860 29934
rect 27580 29708 27636 29764
rect 27916 29372 27972 29428
rect 27244 27916 27300 27972
rect 27804 28476 27860 28532
rect 27468 27692 27524 27748
rect 27356 27020 27412 27076
rect 25676 25506 25732 25508
rect 25676 25454 25678 25506
rect 25678 25454 25730 25506
rect 25730 25454 25732 25506
rect 25676 25452 25732 25454
rect 26348 25506 26404 25508
rect 26348 25454 26350 25506
rect 26350 25454 26402 25506
rect 26402 25454 26404 25506
rect 26348 25452 26404 25454
rect 26460 24610 26516 24612
rect 26460 24558 26462 24610
rect 26462 24558 26514 24610
rect 26514 24558 26516 24610
rect 26460 24556 26516 24558
rect 25452 23660 25508 23716
rect 23100 22146 23156 22148
rect 23100 22094 23102 22146
rect 23102 22094 23154 22146
rect 23154 22094 23156 22146
rect 23100 22092 23156 22094
rect 22764 20748 22820 20804
rect 22652 20690 22708 20692
rect 22652 20638 22654 20690
rect 22654 20638 22706 20690
rect 22706 20638 22708 20690
rect 22652 20636 22708 20638
rect 23212 20690 23268 20692
rect 23212 20638 23214 20690
rect 23214 20638 23266 20690
rect 23266 20638 23268 20690
rect 23212 20636 23268 20638
rect 26348 21756 26404 21812
rect 25900 20188 25956 20244
rect 27244 24834 27300 24836
rect 27244 24782 27246 24834
rect 27246 24782 27298 24834
rect 27298 24782 27300 24834
rect 27244 24780 27300 24782
rect 26908 24220 26964 24276
rect 27020 24556 27076 24612
rect 27132 22428 27188 22484
rect 27244 24220 27300 24276
rect 26908 22204 26964 22260
rect 26684 22092 26740 22148
rect 26796 21644 26852 21700
rect 26908 20690 26964 20692
rect 26908 20638 26910 20690
rect 26910 20638 26962 20690
rect 26962 20638 26964 20690
rect 26908 20636 26964 20638
rect 27468 21980 27524 22036
rect 26796 20188 26852 20244
rect 24220 19180 24276 19236
rect 23884 18284 23940 18340
rect 22428 16604 22484 16660
rect 22652 18172 22708 18228
rect 23436 18172 23492 18228
rect 22876 16940 22932 16996
rect 23996 16882 24052 16884
rect 23996 16830 23998 16882
rect 23998 16830 24050 16882
rect 24050 16830 24052 16882
rect 23996 16828 24052 16830
rect 22988 16716 23044 16772
rect 22316 15820 22372 15876
rect 22316 15372 22372 15428
rect 21532 15260 21588 15316
rect 19852 13634 19908 13636
rect 19852 13582 19854 13634
rect 19854 13582 19906 13634
rect 19906 13582 19908 13634
rect 19852 13580 19908 13582
rect 20300 13858 20356 13860
rect 20300 13806 20302 13858
rect 20302 13806 20354 13858
rect 20354 13806 20356 13858
rect 20300 13804 20356 13806
rect 20412 13746 20468 13748
rect 20412 13694 20414 13746
rect 20414 13694 20466 13746
rect 20466 13694 20468 13746
rect 20412 13692 20468 13694
rect 20860 13746 20916 13748
rect 20860 13694 20862 13746
rect 20862 13694 20914 13746
rect 20914 13694 20916 13746
rect 20860 13692 20916 13694
rect 21980 13916 22036 13972
rect 22204 14306 22260 14308
rect 22204 14254 22206 14306
rect 22206 14254 22258 14306
rect 22258 14254 22260 14306
rect 22204 14252 22260 14254
rect 22204 13692 22260 13748
rect 20076 13132 20132 13188
rect 20188 13074 20244 13076
rect 20188 13022 20190 13074
rect 20190 13022 20242 13074
rect 20242 13022 20244 13074
rect 20188 13020 20244 13022
rect 20636 13074 20692 13076
rect 20636 13022 20638 13074
rect 20638 13022 20690 13074
rect 20690 13022 20692 13074
rect 20636 13020 20692 13022
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19852 12290 19908 12292
rect 19852 12238 19854 12290
rect 19854 12238 19906 12290
rect 19906 12238 19908 12290
rect 19852 12236 19908 12238
rect 19628 11564 19684 11620
rect 21196 11564 21252 11620
rect 20748 11506 20804 11508
rect 20748 11454 20750 11506
rect 20750 11454 20802 11506
rect 20802 11454 20804 11506
rect 20748 11452 20804 11454
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 24220 16716 24276 16772
rect 25788 18508 25844 18564
rect 24556 17500 24612 17556
rect 23100 16268 23156 16324
rect 23100 16098 23156 16100
rect 23100 16046 23102 16098
rect 23102 16046 23154 16098
rect 23154 16046 23156 16098
rect 23100 16044 23156 16046
rect 22540 15596 22596 15652
rect 22876 15202 22932 15204
rect 22876 15150 22878 15202
rect 22878 15150 22930 15202
rect 22930 15150 22932 15202
rect 22876 15148 22932 15150
rect 22652 14530 22708 14532
rect 22652 14478 22654 14530
rect 22654 14478 22706 14530
rect 22706 14478 22708 14530
rect 22652 14476 22708 14478
rect 23884 16098 23940 16100
rect 23884 16046 23886 16098
rect 23886 16046 23938 16098
rect 23938 16046 23940 16098
rect 23884 16044 23940 16046
rect 23772 14588 23828 14644
rect 23660 14252 23716 14308
rect 23436 13916 23492 13972
rect 21756 12402 21812 12404
rect 21756 12350 21758 12402
rect 21758 12350 21810 12402
rect 21810 12350 21812 12402
rect 21756 12348 21812 12350
rect 21756 11618 21812 11620
rect 21756 11566 21758 11618
rect 21758 11566 21810 11618
rect 21810 11566 21812 11618
rect 21756 11564 21812 11566
rect 21532 11452 21588 11508
rect 21420 10668 21476 10724
rect 20972 10220 21028 10276
rect 19516 10108 19572 10164
rect 20636 10108 20692 10164
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19292 7980 19348 8036
rect 19740 8876 19796 8932
rect 19516 8204 19572 8260
rect 20636 9714 20692 9716
rect 20636 9662 20638 9714
rect 20638 9662 20690 9714
rect 20690 9662 20692 9714
rect 20636 9660 20692 9662
rect 21420 10220 21476 10276
rect 21868 9996 21924 10052
rect 22988 13132 23044 13188
rect 22876 12738 22932 12740
rect 22876 12686 22878 12738
rect 22878 12686 22930 12738
rect 22930 12686 22932 12738
rect 22876 12684 22932 12686
rect 22092 12348 22148 12404
rect 22428 11676 22484 11732
rect 22092 11618 22148 11620
rect 22092 11566 22094 11618
rect 22094 11566 22146 11618
rect 22146 11566 22148 11618
rect 22092 11564 22148 11566
rect 22988 12402 23044 12404
rect 22988 12350 22990 12402
rect 22990 12350 23042 12402
rect 23042 12350 23044 12402
rect 22988 12348 23044 12350
rect 23660 12402 23716 12404
rect 23660 12350 23662 12402
rect 23662 12350 23714 12402
rect 23714 12350 23716 12402
rect 23660 12348 23716 12350
rect 22764 11676 22820 11732
rect 22428 11394 22484 11396
rect 22428 11342 22430 11394
rect 22430 11342 22482 11394
rect 22482 11342 22484 11394
rect 22428 11340 22484 11342
rect 22764 11394 22820 11396
rect 22764 11342 22766 11394
rect 22766 11342 22818 11394
rect 22818 11342 22820 11394
rect 22764 11340 22820 11342
rect 22204 11170 22260 11172
rect 22204 11118 22206 11170
rect 22206 11118 22258 11170
rect 22258 11118 22260 11170
rect 22204 11116 22260 11118
rect 22204 10722 22260 10724
rect 22204 10670 22206 10722
rect 22206 10670 22258 10722
rect 22258 10670 22260 10722
rect 22204 10668 22260 10670
rect 22092 10108 22148 10164
rect 22428 9996 22484 10052
rect 20412 8764 20468 8820
rect 20300 8370 20356 8372
rect 20300 8318 20302 8370
rect 20302 8318 20354 8370
rect 20354 8318 20356 8370
rect 20300 8316 20356 8318
rect 21308 8540 21364 8596
rect 21420 8204 21476 8260
rect 21644 8204 21700 8260
rect 19516 7756 19572 7812
rect 19740 7980 19796 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20188 7868 20244 7924
rect 20748 7980 20804 8036
rect 20044 7812 20100 7814
rect 19292 7308 19348 7364
rect 18060 6636 18116 6692
rect 18396 6748 18452 6804
rect 17388 6412 17444 6468
rect 17724 6018 17780 6020
rect 17724 5966 17726 6018
rect 17726 5966 17778 6018
rect 17778 5966 17780 6018
rect 17724 5964 17780 5966
rect 19852 7308 19908 7364
rect 19964 7474 20020 7476
rect 19964 7422 19966 7474
rect 19966 7422 20018 7474
rect 20018 7422 20020 7474
rect 19964 7420 20020 7422
rect 19628 6748 19684 6804
rect 20300 6690 20356 6692
rect 20300 6638 20302 6690
rect 20302 6638 20354 6690
rect 20354 6638 20356 6690
rect 20300 6636 20356 6638
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 18844 6130 18900 6132
rect 18844 6078 18846 6130
rect 18846 6078 18898 6130
rect 18898 6078 18900 6130
rect 18844 6076 18900 6078
rect 16716 5068 16772 5124
rect 17388 5122 17444 5124
rect 17388 5070 17390 5122
rect 17390 5070 17442 5122
rect 17442 5070 17444 5122
rect 17388 5068 17444 5070
rect 17948 4956 18004 5012
rect 17388 4732 17444 4788
rect 20188 5964 20244 6020
rect 21532 8034 21588 8036
rect 21532 7982 21534 8034
rect 21534 7982 21586 8034
rect 21586 7982 21588 8034
rect 21532 7980 21588 7982
rect 24332 15932 24388 15988
rect 24220 15596 24276 15652
rect 24444 15148 24500 15204
rect 24444 14700 24500 14756
rect 26124 18844 26180 18900
rect 25900 18284 25956 18340
rect 26124 17612 26180 17668
rect 25676 16940 25732 16996
rect 24780 16882 24836 16884
rect 24780 16830 24782 16882
rect 24782 16830 24834 16882
rect 24834 16830 24836 16882
rect 24780 16828 24836 16830
rect 25340 16098 25396 16100
rect 25340 16046 25342 16098
rect 25342 16046 25394 16098
rect 25394 16046 25396 16098
rect 25340 16044 25396 16046
rect 25788 16098 25844 16100
rect 25788 16046 25790 16098
rect 25790 16046 25842 16098
rect 25842 16046 25844 16098
rect 25788 16044 25844 16046
rect 24892 15986 24948 15988
rect 24892 15934 24894 15986
rect 24894 15934 24946 15986
rect 24946 15934 24948 15986
rect 24892 15932 24948 15934
rect 25228 15426 25284 15428
rect 25228 15374 25230 15426
rect 25230 15374 25282 15426
rect 25282 15374 25284 15426
rect 25228 15372 25284 15374
rect 25452 15426 25508 15428
rect 25452 15374 25454 15426
rect 25454 15374 25506 15426
rect 25506 15374 25508 15426
rect 25452 15372 25508 15374
rect 24556 14476 24612 14532
rect 24780 13634 24836 13636
rect 24780 13582 24782 13634
rect 24782 13582 24834 13634
rect 24834 13582 24836 13634
rect 24780 13580 24836 13582
rect 25452 14642 25508 14644
rect 25452 14590 25454 14642
rect 25454 14590 25506 14642
rect 25506 14590 25508 14642
rect 25452 14588 25508 14590
rect 25340 14252 25396 14308
rect 25676 15036 25732 15092
rect 26124 17164 26180 17220
rect 26124 16940 26180 16996
rect 26460 17724 26516 17780
rect 27804 27298 27860 27300
rect 27804 27246 27806 27298
rect 27806 27246 27858 27298
rect 27858 27246 27860 27298
rect 27804 27244 27860 27246
rect 28028 29484 28084 29540
rect 29036 29708 29092 29764
rect 28588 29596 28644 29652
rect 28700 29538 28756 29540
rect 28700 29486 28702 29538
rect 28702 29486 28754 29538
rect 28754 29486 28756 29538
rect 28700 29484 28756 29486
rect 28252 28082 28308 28084
rect 28252 28030 28254 28082
rect 28254 28030 28306 28082
rect 28306 28030 28308 28082
rect 28252 28028 28308 28030
rect 28812 28700 28868 28756
rect 28700 28642 28756 28644
rect 28700 28590 28702 28642
rect 28702 28590 28754 28642
rect 28754 28590 28756 28642
rect 28700 28588 28756 28590
rect 28364 27970 28420 27972
rect 28364 27918 28366 27970
rect 28366 27918 28418 27970
rect 28418 27918 28420 27970
rect 28364 27916 28420 27918
rect 27804 24834 27860 24836
rect 27804 24782 27806 24834
rect 27806 24782 27858 24834
rect 27858 24782 27860 24834
rect 27804 24780 27860 24782
rect 27804 23548 27860 23604
rect 28588 25282 28644 25284
rect 28588 25230 28590 25282
rect 28590 25230 28642 25282
rect 28642 25230 28644 25282
rect 28588 25228 28644 25230
rect 28140 23714 28196 23716
rect 28140 23662 28142 23714
rect 28142 23662 28194 23714
rect 28194 23662 28196 23714
rect 28140 23660 28196 23662
rect 29260 29426 29316 29428
rect 29260 29374 29262 29426
rect 29262 29374 29314 29426
rect 29314 29374 29316 29426
rect 29260 29372 29316 29374
rect 29708 30044 29764 30100
rect 29708 29708 29764 29764
rect 31052 36316 31108 36372
rect 31164 34802 31220 34804
rect 31164 34750 31166 34802
rect 31166 34750 31218 34802
rect 31218 34750 31220 34802
rect 31164 34748 31220 34750
rect 31052 34242 31108 34244
rect 31052 34190 31054 34242
rect 31054 34190 31106 34242
rect 31106 34190 31108 34242
rect 31052 34188 31108 34190
rect 30604 33628 30660 33684
rect 32732 36370 32788 36372
rect 32732 36318 32734 36370
rect 32734 36318 32786 36370
rect 32786 36318 32788 36370
rect 32732 36316 32788 36318
rect 31836 35308 31892 35364
rect 32284 35026 32340 35028
rect 32284 34974 32286 35026
rect 32286 34974 32338 35026
rect 32338 34974 32340 35026
rect 32284 34972 32340 34974
rect 32396 34300 32452 34356
rect 32284 34242 32340 34244
rect 32284 34190 32286 34242
rect 32286 34190 32338 34242
rect 32338 34190 32340 34242
rect 32284 34188 32340 34190
rect 31948 34130 32004 34132
rect 31948 34078 31950 34130
rect 31950 34078 32002 34130
rect 32002 34078 32004 34130
rect 31948 34076 32004 34078
rect 32060 34018 32116 34020
rect 32060 33966 32062 34018
rect 32062 33966 32114 34018
rect 32114 33966 32116 34018
rect 32060 33964 32116 33966
rect 32508 35532 32564 35588
rect 32508 33628 32564 33684
rect 31836 32002 31892 32004
rect 31836 31950 31838 32002
rect 31838 31950 31890 32002
rect 31890 31950 31892 32002
rect 31836 31948 31892 31950
rect 31052 31890 31108 31892
rect 31052 31838 31054 31890
rect 31054 31838 31106 31890
rect 31106 31838 31108 31890
rect 31052 31836 31108 31838
rect 30716 30268 30772 30324
rect 30268 30156 30324 30212
rect 30604 30044 30660 30100
rect 31612 31388 31668 31444
rect 31612 30828 31668 30884
rect 31500 30770 31556 30772
rect 31500 30718 31502 30770
rect 31502 30718 31554 30770
rect 31554 30718 31556 30770
rect 31500 30716 31556 30718
rect 31276 30380 31332 30436
rect 30156 29372 30212 29428
rect 29596 28700 29652 28756
rect 29820 29036 29876 29092
rect 29708 28642 29764 28644
rect 29708 28590 29710 28642
rect 29710 28590 29762 28642
rect 29762 28590 29764 28642
rect 29708 28588 29764 28590
rect 30268 28812 30324 28868
rect 29820 28530 29876 28532
rect 29820 28478 29822 28530
rect 29822 28478 29874 28530
rect 29874 28478 29876 28530
rect 29820 28476 29876 28478
rect 29148 27970 29204 27972
rect 29148 27918 29150 27970
rect 29150 27918 29202 27970
rect 29202 27918 29204 27970
rect 29148 27916 29204 27918
rect 29596 27858 29652 27860
rect 29596 27806 29598 27858
rect 29598 27806 29650 27858
rect 29650 27806 29652 27858
rect 29596 27804 29652 27806
rect 29260 27746 29316 27748
rect 29260 27694 29262 27746
rect 29262 27694 29314 27746
rect 29314 27694 29316 27746
rect 29260 27692 29316 27694
rect 30828 29426 30884 29428
rect 30828 29374 30830 29426
rect 30830 29374 30882 29426
rect 30882 29374 30884 29426
rect 30828 29372 30884 29374
rect 30716 29036 30772 29092
rect 30716 28866 30772 28868
rect 30716 28814 30718 28866
rect 30718 28814 30770 28866
rect 30770 28814 30772 28866
rect 30716 28812 30772 28814
rect 31276 29484 31332 29540
rect 33852 41244 33908 41300
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 33068 40402 33124 40404
rect 33068 40350 33070 40402
rect 33070 40350 33122 40402
rect 33122 40350 33124 40402
rect 33068 40348 33124 40350
rect 33516 40402 33572 40404
rect 33516 40350 33518 40402
rect 33518 40350 33570 40402
rect 33570 40350 33572 40402
rect 33516 40348 33572 40350
rect 33740 40236 33796 40292
rect 33964 40124 34020 40180
rect 34412 40290 34468 40292
rect 34412 40238 34414 40290
rect 34414 40238 34466 40290
rect 34466 40238 34468 40290
rect 34412 40236 34468 40238
rect 34076 39788 34132 39844
rect 34524 40124 34580 40180
rect 33068 38834 33124 38836
rect 33068 38782 33070 38834
rect 33070 38782 33122 38834
rect 33122 38782 33124 38834
rect 33068 38780 33124 38782
rect 34860 39564 34916 39620
rect 34524 38668 34580 38724
rect 35084 40348 35140 40404
rect 35196 40124 35252 40180
rect 35868 40962 35924 40964
rect 35868 40910 35870 40962
rect 35870 40910 35922 40962
rect 35922 40910 35924 40962
rect 35868 40908 35924 40910
rect 36428 40348 36484 40404
rect 35644 40236 35700 40292
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35308 39788 35364 39844
rect 35980 40236 36036 40292
rect 33292 38050 33348 38052
rect 33292 37998 33294 38050
rect 33294 37998 33346 38050
rect 33346 37998 33348 38050
rect 33292 37996 33348 37998
rect 34076 38050 34132 38052
rect 34076 37998 34078 38050
rect 34078 37998 34130 38050
rect 34130 37998 34132 38050
rect 34076 37996 34132 37998
rect 34748 37996 34804 38052
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 36316 39058 36372 39060
rect 36316 39006 36318 39058
rect 36318 39006 36370 39058
rect 36370 39006 36372 39058
rect 36316 39004 36372 39006
rect 37548 40684 37604 40740
rect 36988 39618 37044 39620
rect 36988 39566 36990 39618
rect 36990 39566 37042 39618
rect 37042 39566 37044 39618
rect 36988 39564 37044 39566
rect 35980 38722 36036 38724
rect 35980 38670 35982 38722
rect 35982 38670 36034 38722
rect 36034 38670 36036 38722
rect 35980 38668 36036 38670
rect 38108 40684 38164 40740
rect 39340 41020 39396 41076
rect 39116 40626 39172 40628
rect 39116 40574 39118 40626
rect 39118 40574 39170 40626
rect 39170 40574 39172 40626
rect 39116 40572 39172 40574
rect 37324 38668 37380 38724
rect 37436 38780 37492 38836
rect 37884 40460 37940 40516
rect 39788 40236 39844 40292
rect 39004 39676 39060 39732
rect 38892 39004 38948 39060
rect 37548 38556 37604 38612
rect 35420 37996 35476 38052
rect 36988 38108 37044 38164
rect 33068 37212 33124 37268
rect 33964 37266 34020 37268
rect 33964 37214 33966 37266
rect 33966 37214 34018 37266
rect 34018 37214 34020 37266
rect 33964 37212 34020 37214
rect 35084 37212 35140 37268
rect 32956 35756 33012 35812
rect 34860 35756 34916 35812
rect 33180 34972 33236 35028
rect 33292 35308 33348 35364
rect 33628 34972 33684 35028
rect 34412 34636 34468 34692
rect 33516 34188 33572 34244
rect 33852 34018 33908 34020
rect 33852 33966 33854 34018
rect 33854 33966 33906 34018
rect 33906 33966 33908 34018
rect 33852 33964 33908 33966
rect 34524 33852 34580 33908
rect 33852 33068 33908 33124
rect 33180 31948 33236 32004
rect 34972 32450 35028 32452
rect 34972 32398 34974 32450
rect 34974 32398 35026 32450
rect 35026 32398 35028 32450
rect 34972 32396 35028 32398
rect 35868 37212 35924 37268
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35532 35810 35588 35812
rect 35532 35758 35534 35810
rect 35534 35758 35586 35810
rect 35586 35758 35588 35810
rect 35532 35756 35588 35758
rect 35420 35586 35476 35588
rect 35420 35534 35422 35586
rect 35422 35534 35474 35586
rect 35474 35534 35476 35586
rect 35420 35532 35476 35534
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35420 34972 35476 35028
rect 35308 34914 35364 34916
rect 35308 34862 35310 34914
rect 35310 34862 35362 34914
rect 35362 34862 35364 34914
rect 35308 34860 35364 34862
rect 35644 34972 35700 35028
rect 36764 37266 36820 37268
rect 36764 37214 36766 37266
rect 36766 37214 36818 37266
rect 36818 37214 36820 37266
rect 36764 37212 36820 37214
rect 38108 38556 38164 38612
rect 35980 35922 36036 35924
rect 35980 35870 35982 35922
rect 35982 35870 36034 35922
rect 36034 35870 36036 35922
rect 35980 35868 36036 35870
rect 37212 35868 37268 35924
rect 36764 35810 36820 35812
rect 36764 35758 36766 35810
rect 36766 35758 36818 35810
rect 36818 35758 36820 35810
rect 36764 35756 36820 35758
rect 36316 35698 36372 35700
rect 36316 35646 36318 35698
rect 36318 35646 36370 35698
rect 36370 35646 36372 35698
rect 36316 35644 36372 35646
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35420 33570 35476 33572
rect 35420 33518 35422 33570
rect 35422 33518 35474 33570
rect 35474 33518 35476 33570
rect 35420 33516 35476 33518
rect 35756 33516 35812 33572
rect 35532 33346 35588 33348
rect 35532 33294 35534 33346
rect 35534 33294 35586 33346
rect 35586 33294 35588 33346
rect 35532 33292 35588 33294
rect 35644 33180 35700 33236
rect 35196 32562 35252 32564
rect 35196 32510 35198 32562
rect 35198 32510 35250 32562
rect 35250 32510 35252 32562
rect 35196 32508 35252 32510
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 31724 29932 31780 29988
rect 33068 31106 33124 31108
rect 33068 31054 33070 31106
rect 33070 31054 33122 31106
rect 33122 31054 33124 31106
rect 33068 31052 33124 31054
rect 32620 30940 32676 30996
rect 31948 29820 32004 29876
rect 32508 29596 32564 29652
rect 31724 28812 31780 28868
rect 32396 29202 32452 29204
rect 32396 29150 32398 29202
rect 32398 29150 32450 29202
rect 32450 29150 32452 29202
rect 32396 29148 32452 29150
rect 31948 28588 32004 28644
rect 30268 28364 30324 28420
rect 30268 27916 30324 27972
rect 30380 27746 30436 27748
rect 30380 27694 30382 27746
rect 30382 27694 30434 27746
rect 30434 27694 30436 27746
rect 30380 27692 30436 27694
rect 30044 26348 30100 26404
rect 30828 26402 30884 26404
rect 30828 26350 30830 26402
rect 30830 26350 30882 26402
rect 30882 26350 30884 26402
rect 30828 26348 30884 26350
rect 31836 26012 31892 26068
rect 29260 25282 29316 25284
rect 29260 25230 29262 25282
rect 29262 25230 29314 25282
rect 29314 25230 29316 25282
rect 29260 25228 29316 25230
rect 32508 28364 32564 28420
rect 31948 25452 32004 25508
rect 31724 25228 31780 25284
rect 29484 23938 29540 23940
rect 29484 23886 29486 23938
rect 29486 23886 29538 23938
rect 29538 23886 29540 23938
rect 29484 23884 29540 23886
rect 28812 23212 28868 23268
rect 28924 23660 28980 23716
rect 28476 23154 28532 23156
rect 28476 23102 28478 23154
rect 28478 23102 28530 23154
rect 28530 23102 28532 23154
rect 28476 23100 28532 23102
rect 28140 22652 28196 22708
rect 27804 22204 27860 22260
rect 27916 22428 27972 22484
rect 27692 21532 27748 21588
rect 27804 21868 27860 21924
rect 28588 22258 28644 22260
rect 28588 22206 28590 22258
rect 28590 22206 28642 22258
rect 28642 22206 28644 22258
rect 28588 22204 28644 22206
rect 28812 23042 28868 23044
rect 28812 22990 28814 23042
rect 28814 22990 28866 23042
rect 28866 22990 28868 23042
rect 28812 22988 28868 22990
rect 28700 21868 28756 21924
rect 28140 21756 28196 21812
rect 28588 21698 28644 21700
rect 28588 21646 28590 21698
rect 28590 21646 28642 21698
rect 28642 21646 28644 21698
rect 28588 21644 28644 21646
rect 29036 22988 29092 23044
rect 29260 23548 29316 23604
rect 29148 22204 29204 22260
rect 29036 21980 29092 22036
rect 28588 21362 28644 21364
rect 28588 21310 28590 21362
rect 28590 21310 28642 21362
rect 28642 21310 28644 21362
rect 28588 21308 28644 21310
rect 27580 20412 27636 20468
rect 28476 20636 28532 20692
rect 27916 20130 27972 20132
rect 27916 20078 27918 20130
rect 27918 20078 27970 20130
rect 27970 20078 27972 20130
rect 27916 20076 27972 20078
rect 27580 19010 27636 19012
rect 27580 18958 27582 19010
rect 27582 18958 27634 19010
rect 27634 18958 27636 19010
rect 27580 18956 27636 18958
rect 27580 17836 27636 17892
rect 27916 19122 27972 19124
rect 27916 19070 27918 19122
rect 27918 19070 27970 19122
rect 27970 19070 27972 19122
rect 27916 19068 27972 19070
rect 27692 18396 27748 18452
rect 27804 18508 27860 18564
rect 26796 17778 26852 17780
rect 26796 17726 26798 17778
rect 26798 17726 26850 17778
rect 26850 17726 26852 17778
rect 26796 17724 26852 17726
rect 26796 17164 26852 17220
rect 26684 16156 26740 16212
rect 26348 15596 26404 15652
rect 26348 15426 26404 15428
rect 26348 15374 26350 15426
rect 26350 15374 26402 15426
rect 26402 15374 26404 15426
rect 26348 15372 26404 15374
rect 26236 15260 26292 15316
rect 26012 14700 26068 14756
rect 25788 14588 25844 14644
rect 25228 13580 25284 13636
rect 26124 14418 26180 14420
rect 26124 14366 26126 14418
rect 26126 14366 26178 14418
rect 26178 14366 26180 14418
rect 26124 14364 26180 14366
rect 26460 14700 26516 14756
rect 26796 16828 26852 16884
rect 26908 16716 26964 16772
rect 27356 17666 27412 17668
rect 27356 17614 27358 17666
rect 27358 17614 27410 17666
rect 27410 17614 27412 17666
rect 27356 17612 27412 17614
rect 27916 18172 27972 18228
rect 28252 20076 28308 20132
rect 28476 20412 28532 20468
rect 28700 19404 28756 19460
rect 28364 18562 28420 18564
rect 28364 18510 28366 18562
rect 28366 18510 28418 18562
rect 28418 18510 28420 18562
rect 28364 18508 28420 18510
rect 28252 18450 28308 18452
rect 28252 18398 28254 18450
rect 28254 18398 28306 18450
rect 28306 18398 28308 18450
rect 28252 18396 28308 18398
rect 28476 18172 28532 18228
rect 28252 17724 28308 17780
rect 27356 16828 27412 16884
rect 27020 16268 27076 16324
rect 26908 15708 26964 15764
rect 27580 16716 27636 16772
rect 26908 15372 26964 15428
rect 27132 15372 27188 15428
rect 26796 15036 26852 15092
rect 27020 15260 27076 15316
rect 27132 15148 27188 15204
rect 27692 16044 27748 16100
rect 27692 15372 27748 15428
rect 27020 14252 27076 14308
rect 27916 15260 27972 15316
rect 27804 15148 27860 15204
rect 28588 17388 28644 17444
rect 28476 16882 28532 16884
rect 28476 16830 28478 16882
rect 28478 16830 28530 16882
rect 28530 16830 28532 16882
rect 28476 16828 28532 16830
rect 28140 16268 28196 16324
rect 28140 15932 28196 15988
rect 28140 15484 28196 15540
rect 28476 15708 28532 15764
rect 28588 16268 28644 16324
rect 28924 18396 28980 18452
rect 28700 15820 28756 15876
rect 28812 15372 28868 15428
rect 28476 15314 28532 15316
rect 28476 15262 28478 15314
rect 28478 15262 28530 15314
rect 28530 15262 28532 15314
rect 28476 15260 28532 15262
rect 28364 14700 28420 14756
rect 28588 15148 28644 15204
rect 28252 14642 28308 14644
rect 28252 14590 28254 14642
rect 28254 14590 28306 14642
rect 28306 14590 28308 14642
rect 28252 14588 28308 14590
rect 27804 14530 27860 14532
rect 27804 14478 27806 14530
rect 27806 14478 27858 14530
rect 27858 14478 27860 14530
rect 27804 14476 27860 14478
rect 27132 13970 27188 13972
rect 27132 13918 27134 13970
rect 27134 13918 27186 13970
rect 27186 13918 27188 13970
rect 27132 13916 27188 13918
rect 26572 13692 26628 13748
rect 27132 13692 27188 13748
rect 26908 13580 26964 13636
rect 27244 12850 27300 12852
rect 27244 12798 27246 12850
rect 27246 12798 27298 12850
rect 27298 12798 27300 12850
rect 27244 12796 27300 12798
rect 27916 12178 27972 12180
rect 27916 12126 27918 12178
rect 27918 12126 27970 12178
rect 27970 12126 27972 12178
rect 27916 12124 27972 12126
rect 27692 11618 27748 11620
rect 27692 11566 27694 11618
rect 27694 11566 27746 11618
rect 27746 11566 27748 11618
rect 27692 11564 27748 11566
rect 23996 11340 24052 11396
rect 24556 11452 24612 11508
rect 23996 11116 24052 11172
rect 23212 10722 23268 10724
rect 23212 10670 23214 10722
rect 23214 10670 23266 10722
rect 23266 10670 23268 10722
rect 23212 10668 23268 10670
rect 22764 9660 22820 9716
rect 22988 9996 23044 10052
rect 25676 11506 25732 11508
rect 25676 11454 25678 11506
rect 25678 11454 25730 11506
rect 25730 11454 25732 11506
rect 25676 11452 25732 11454
rect 22652 8764 22708 8820
rect 22540 8652 22596 8708
rect 22764 8540 22820 8596
rect 23324 8652 23380 8708
rect 22876 8428 22932 8484
rect 21644 7868 21700 7924
rect 22092 7532 22148 7588
rect 22316 7980 22372 8036
rect 22540 7980 22596 8036
rect 22764 8034 22820 8036
rect 22764 7982 22766 8034
rect 22766 7982 22818 8034
rect 22818 7982 22820 8034
rect 22764 7980 22820 7982
rect 24332 9154 24388 9156
rect 24332 9102 24334 9154
rect 24334 9102 24386 9154
rect 24386 9102 24388 9154
rect 24332 9100 24388 9102
rect 26572 11282 26628 11284
rect 26572 11230 26574 11282
rect 26574 11230 26626 11282
rect 26626 11230 26628 11282
rect 26572 11228 26628 11230
rect 27356 11282 27412 11284
rect 27356 11230 27358 11282
rect 27358 11230 27410 11282
rect 27410 11230 27412 11282
rect 27356 11228 27412 11230
rect 27692 10610 27748 10612
rect 27692 10558 27694 10610
rect 27694 10558 27746 10610
rect 27746 10558 27748 10610
rect 27692 10556 27748 10558
rect 26908 9660 26964 9716
rect 25340 9100 25396 9156
rect 25788 9154 25844 9156
rect 25788 9102 25790 9154
rect 25790 9102 25842 9154
rect 25842 9102 25844 9154
rect 25788 9100 25844 9102
rect 24220 8818 24276 8820
rect 24220 8766 24222 8818
rect 24222 8766 24274 8818
rect 24274 8766 24276 8818
rect 24220 8764 24276 8766
rect 23772 8652 23828 8708
rect 23324 7980 23380 8036
rect 25116 8204 25172 8260
rect 22764 7756 22820 7812
rect 22316 7474 22372 7476
rect 22316 7422 22318 7474
rect 22318 7422 22370 7474
rect 22370 7422 22372 7474
rect 22316 7420 22372 7422
rect 24668 7698 24724 7700
rect 24668 7646 24670 7698
rect 24670 7646 24722 7698
rect 24722 7646 24724 7698
rect 24668 7644 24724 7646
rect 21420 6690 21476 6692
rect 21420 6638 21422 6690
rect 21422 6638 21474 6690
rect 21474 6638 21476 6690
rect 21420 6636 21476 6638
rect 24556 7586 24612 7588
rect 24556 7534 24558 7586
rect 24558 7534 24610 7586
rect 24610 7534 24612 7586
rect 24556 7532 24612 7534
rect 24892 7420 24948 7476
rect 24556 6748 24612 6804
rect 22764 6636 22820 6692
rect 22428 6524 22484 6580
rect 20860 5964 20916 6020
rect 18844 4956 18900 5012
rect 28364 13916 28420 13972
rect 29260 20690 29316 20692
rect 29260 20638 29262 20690
rect 29262 20638 29314 20690
rect 29314 20638 29316 20690
rect 29260 20636 29316 20638
rect 29148 20412 29204 20468
rect 31612 23378 31668 23380
rect 31612 23326 31614 23378
rect 31614 23326 31666 23378
rect 31666 23326 31668 23378
rect 31612 23324 31668 23326
rect 30380 23212 30436 23268
rect 30044 23100 30100 23156
rect 29484 22258 29540 22260
rect 29484 22206 29486 22258
rect 29486 22206 29538 22258
rect 29538 22206 29540 22258
rect 29484 22204 29540 22206
rect 31052 23266 31108 23268
rect 31052 23214 31054 23266
rect 31054 23214 31106 23266
rect 31106 23214 31108 23266
rect 31052 23212 31108 23214
rect 30604 23154 30660 23156
rect 30604 23102 30606 23154
rect 30606 23102 30658 23154
rect 30658 23102 30660 23154
rect 30604 23100 30660 23102
rect 31612 22988 31668 23044
rect 32284 23884 32340 23940
rect 32396 23324 32452 23380
rect 31724 23100 31780 23156
rect 30044 22204 30100 22260
rect 29484 20690 29540 20692
rect 29484 20638 29486 20690
rect 29486 20638 29538 20690
rect 29538 20638 29540 20690
rect 29484 20636 29540 20638
rect 29372 20300 29428 20356
rect 29260 20188 29316 20244
rect 29148 20076 29204 20132
rect 29596 20188 29652 20244
rect 29148 19234 29204 19236
rect 29148 19182 29150 19234
rect 29150 19182 29202 19234
rect 29202 19182 29204 19234
rect 29148 19180 29204 19182
rect 29820 20076 29876 20132
rect 32396 23154 32452 23156
rect 32396 23102 32398 23154
rect 32398 23102 32450 23154
rect 32450 23102 32452 23154
rect 32396 23100 32452 23102
rect 31836 21980 31892 22036
rect 31948 22428 32004 22484
rect 30828 21532 30884 21588
rect 30492 19964 30548 20020
rect 30044 19180 30100 19236
rect 30156 19740 30212 19796
rect 29708 18956 29764 19012
rect 30156 19068 30212 19124
rect 29596 18620 29652 18676
rect 29484 18284 29540 18340
rect 30604 18620 30660 18676
rect 30716 18338 30772 18340
rect 30716 18286 30718 18338
rect 30718 18286 30770 18338
rect 30770 18286 30772 18338
rect 30716 18284 30772 18286
rect 29932 18172 29988 18228
rect 29372 17442 29428 17444
rect 29372 17390 29374 17442
rect 29374 17390 29426 17442
rect 29426 17390 29428 17442
rect 29372 17388 29428 17390
rect 29148 16716 29204 16772
rect 29484 16770 29540 16772
rect 29484 16718 29486 16770
rect 29486 16718 29538 16770
rect 29538 16718 29540 16770
rect 29484 16716 29540 16718
rect 29148 16492 29204 16548
rect 29484 16098 29540 16100
rect 29484 16046 29486 16098
rect 29486 16046 29538 16098
rect 29538 16046 29540 16098
rect 29484 16044 29540 16046
rect 29372 15260 29428 15316
rect 28812 14588 28868 14644
rect 28812 13020 28868 13076
rect 28140 12796 28196 12852
rect 28588 12572 28644 12628
rect 29148 14530 29204 14532
rect 29148 14478 29150 14530
rect 29150 14478 29202 14530
rect 29202 14478 29204 14530
rect 29148 14476 29204 14478
rect 29708 16210 29764 16212
rect 29708 16158 29710 16210
rect 29710 16158 29762 16210
rect 29762 16158 29764 16210
rect 29708 16156 29764 16158
rect 29596 14140 29652 14196
rect 31724 21586 31780 21588
rect 31724 21534 31726 21586
rect 31726 21534 31778 21586
rect 31778 21534 31780 21586
rect 31724 21532 31780 21534
rect 32396 21532 32452 21588
rect 31052 19964 31108 20020
rect 31388 19906 31444 19908
rect 31388 19854 31390 19906
rect 31390 19854 31442 19906
rect 31442 19854 31444 19906
rect 31388 19852 31444 19854
rect 31164 19292 31220 19348
rect 31724 18284 31780 18340
rect 32060 20130 32116 20132
rect 32060 20078 32062 20130
rect 32062 20078 32114 20130
rect 32114 20078 32116 20130
rect 32060 20076 32116 20078
rect 32060 19346 32116 19348
rect 32060 19294 32062 19346
rect 32062 19294 32114 19346
rect 32114 19294 32116 19346
rect 32060 19292 32116 19294
rect 32508 20636 32564 20692
rect 32396 19906 32452 19908
rect 32396 19854 32398 19906
rect 32398 19854 32450 19906
rect 32450 19854 32452 19906
rect 32396 19852 32452 19854
rect 31164 17388 31220 17444
rect 30828 17106 30884 17108
rect 30828 17054 30830 17106
rect 30830 17054 30882 17106
rect 30882 17054 30884 17106
rect 30828 17052 30884 17054
rect 29932 16882 29988 16884
rect 29932 16830 29934 16882
rect 29934 16830 29986 16882
rect 29986 16830 29988 16882
rect 29932 16828 29988 16830
rect 30716 16828 30772 16884
rect 30604 16156 30660 16212
rect 30044 15986 30100 15988
rect 30044 15934 30046 15986
rect 30046 15934 30098 15986
rect 30098 15934 30100 15986
rect 30044 15932 30100 15934
rect 30380 15874 30436 15876
rect 30380 15822 30382 15874
rect 30382 15822 30434 15874
rect 30434 15822 30436 15874
rect 30380 15820 30436 15822
rect 30716 15708 30772 15764
rect 30828 16268 30884 16324
rect 30380 15426 30436 15428
rect 30380 15374 30382 15426
rect 30382 15374 30434 15426
rect 30434 15374 30436 15426
rect 30380 15372 30436 15374
rect 29820 13356 29876 13412
rect 30044 15260 30100 15316
rect 30268 14306 30324 14308
rect 30268 14254 30270 14306
rect 30270 14254 30322 14306
rect 30322 14254 30324 14306
rect 30268 14252 30324 14254
rect 30716 14476 30772 14532
rect 30044 13074 30100 13076
rect 30044 13022 30046 13074
rect 30046 13022 30098 13074
rect 30098 13022 30100 13074
rect 30044 13020 30100 13022
rect 28028 11340 28084 11396
rect 28812 12236 28868 12292
rect 28588 12178 28644 12180
rect 28588 12126 28590 12178
rect 28590 12126 28642 12178
rect 28642 12126 28644 12178
rect 28588 12124 28644 12126
rect 27804 9324 27860 9380
rect 25564 8258 25620 8260
rect 25564 8206 25566 8258
rect 25566 8206 25618 8258
rect 25618 8206 25620 8258
rect 25564 8204 25620 8206
rect 25228 7644 25284 7700
rect 25228 7474 25284 7476
rect 25228 7422 25230 7474
rect 25230 7422 25282 7474
rect 25282 7422 25284 7474
rect 25228 7420 25284 7422
rect 29820 11394 29876 11396
rect 29820 11342 29822 11394
rect 29822 11342 29874 11394
rect 29874 11342 29876 11394
rect 29820 11340 29876 11342
rect 29484 11282 29540 11284
rect 29484 11230 29486 11282
rect 29486 11230 29538 11282
rect 29538 11230 29540 11282
rect 29484 11228 29540 11230
rect 29036 9100 29092 9156
rect 31052 15596 31108 15652
rect 30940 15372 30996 15428
rect 31612 15874 31668 15876
rect 31612 15822 31614 15874
rect 31614 15822 31666 15874
rect 31666 15822 31668 15874
rect 31612 15820 31668 15822
rect 31388 15596 31444 15652
rect 31276 15484 31332 15540
rect 31388 15426 31444 15428
rect 31388 15374 31390 15426
rect 31390 15374 31442 15426
rect 31442 15374 31444 15426
rect 31388 15372 31444 15374
rect 32172 18450 32228 18452
rect 32172 18398 32174 18450
rect 32174 18398 32226 18450
rect 32226 18398 32228 18450
rect 32172 18396 32228 18398
rect 32508 18338 32564 18340
rect 32508 18286 32510 18338
rect 32510 18286 32562 18338
rect 32562 18286 32564 18338
rect 32508 18284 32564 18286
rect 33292 30994 33348 30996
rect 33292 30942 33294 30994
rect 33294 30942 33346 30994
rect 33346 30942 33348 30994
rect 33292 30940 33348 30942
rect 34076 30828 34132 30884
rect 33740 30434 33796 30436
rect 33740 30382 33742 30434
rect 33742 30382 33794 30434
rect 33794 30382 33796 30434
rect 33740 30380 33796 30382
rect 33404 30322 33460 30324
rect 33404 30270 33406 30322
rect 33406 30270 33458 30322
rect 33458 30270 33460 30322
rect 33404 30268 33460 30270
rect 33628 30268 33684 30324
rect 32732 29708 32788 29764
rect 33068 29538 33124 29540
rect 33068 29486 33070 29538
rect 33070 29486 33122 29538
rect 33122 29486 33124 29538
rect 33068 29484 33124 29486
rect 35980 34860 36036 34916
rect 36428 34860 36484 34916
rect 36988 34972 37044 35028
rect 36204 34636 36260 34692
rect 36092 34524 36148 34580
rect 36204 34412 36260 34468
rect 37100 34748 37156 34804
rect 38220 38108 38276 38164
rect 38444 38892 38500 38948
rect 39228 38834 39284 38836
rect 39228 38782 39230 38834
rect 39230 38782 39282 38834
rect 39282 38782 39284 38834
rect 39228 38780 39284 38782
rect 38780 38668 38836 38724
rect 39900 39116 39956 39172
rect 39788 39058 39844 39060
rect 39788 39006 39790 39058
rect 39790 39006 39842 39058
rect 39842 39006 39844 39058
rect 39788 39004 39844 39006
rect 39676 38946 39732 38948
rect 39676 38894 39678 38946
rect 39678 38894 39730 38946
rect 39730 38894 39732 38946
rect 39676 38892 39732 38894
rect 37660 37100 37716 37156
rect 38220 37266 38276 37268
rect 38220 37214 38222 37266
rect 38222 37214 38274 37266
rect 38274 37214 38276 37266
rect 38220 37212 38276 37214
rect 37660 35868 37716 35924
rect 37436 35698 37492 35700
rect 37436 35646 37438 35698
rect 37438 35646 37490 35698
rect 37490 35646 37492 35698
rect 37436 35644 37492 35646
rect 35868 33404 35924 33460
rect 36204 33964 36260 34020
rect 36316 33628 36372 33684
rect 35980 32674 36036 32676
rect 35980 32622 35982 32674
rect 35982 32622 36034 32674
rect 36034 32622 36036 32674
rect 35980 32620 36036 32622
rect 36204 33122 36260 33124
rect 36204 33070 36206 33122
rect 36206 33070 36258 33122
rect 36258 33070 36260 33122
rect 36204 33068 36260 33070
rect 36540 34130 36596 34132
rect 36540 34078 36542 34130
rect 36542 34078 36594 34130
rect 36594 34078 36596 34130
rect 36540 34076 36596 34078
rect 36652 33964 36708 34020
rect 36428 33516 36484 33572
rect 37324 34412 37380 34468
rect 37772 34636 37828 34692
rect 37324 33906 37380 33908
rect 37324 33854 37326 33906
rect 37326 33854 37378 33906
rect 37378 33854 37380 33906
rect 37324 33852 37380 33854
rect 37660 33628 37716 33684
rect 37436 33180 37492 33236
rect 36764 32674 36820 32676
rect 36764 32622 36766 32674
rect 36766 32622 36818 32674
rect 36818 32622 36820 32674
rect 36764 32620 36820 32622
rect 36316 32396 36372 32452
rect 35308 31836 35364 31892
rect 35308 30716 35364 30772
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35084 30268 35140 30324
rect 33628 29986 33684 29988
rect 33628 29934 33630 29986
rect 33630 29934 33682 29986
rect 33682 29934 33684 29986
rect 33628 29932 33684 29934
rect 34188 29650 34244 29652
rect 34188 29598 34190 29650
rect 34190 29598 34242 29650
rect 34242 29598 34244 29650
rect 34188 29596 34244 29598
rect 34748 29426 34804 29428
rect 34748 29374 34750 29426
rect 34750 29374 34802 29426
rect 34802 29374 34804 29426
rect 34748 29372 34804 29374
rect 37100 31948 37156 32004
rect 36876 30604 36932 30660
rect 37660 33404 37716 33460
rect 39116 38556 39172 38612
rect 39452 37266 39508 37268
rect 39452 37214 39454 37266
rect 39454 37214 39506 37266
rect 39506 37214 39508 37266
rect 39452 37212 39508 37214
rect 39676 37212 39732 37268
rect 39004 35698 39060 35700
rect 39004 35646 39006 35698
rect 39006 35646 39058 35698
rect 39058 35646 39060 35698
rect 39004 35644 39060 35646
rect 38108 34524 38164 34580
rect 38668 34412 38724 34468
rect 39228 34412 39284 34468
rect 39452 34300 39508 34356
rect 39340 34242 39396 34244
rect 39340 34190 39342 34242
rect 39342 34190 39394 34242
rect 39394 34190 39396 34242
rect 39340 34188 39396 34190
rect 38332 33852 38388 33908
rect 38668 34076 38724 34132
rect 38108 33292 38164 33348
rect 37884 32508 37940 32564
rect 38780 33234 38836 33236
rect 38780 33182 38782 33234
rect 38782 33182 38834 33234
rect 38834 33182 38836 33234
rect 38780 33180 38836 33182
rect 37212 31836 37268 31892
rect 36988 30828 37044 30884
rect 37436 30604 37492 30660
rect 36540 30044 36596 30100
rect 37100 30098 37156 30100
rect 37100 30046 37102 30098
rect 37102 30046 37154 30098
rect 37154 30046 37156 30098
rect 37100 30044 37156 30046
rect 35756 29372 35812 29428
rect 34300 29314 34356 29316
rect 34300 29262 34302 29314
rect 34302 29262 34354 29314
rect 34354 29262 34356 29314
rect 34300 29260 34356 29262
rect 38892 32508 38948 32564
rect 37996 31836 38052 31892
rect 38668 31836 38724 31892
rect 40012 38556 40068 38612
rect 40236 40514 40292 40516
rect 40236 40462 40238 40514
rect 40238 40462 40290 40514
rect 40290 40462 40292 40514
rect 40236 40460 40292 40462
rect 41804 42028 41860 42084
rect 40796 40460 40852 40516
rect 40908 40684 40964 40740
rect 40236 40178 40292 40180
rect 40236 40126 40238 40178
rect 40238 40126 40290 40178
rect 40290 40126 40292 40178
rect 40236 40124 40292 40126
rect 40460 39004 40516 39060
rect 40572 39676 40628 39732
rect 40124 38050 40180 38052
rect 40124 37998 40126 38050
rect 40126 37998 40178 38050
rect 40178 37998 40180 38050
rect 40124 37996 40180 37998
rect 40236 37826 40292 37828
rect 40236 37774 40238 37826
rect 40238 37774 40290 37826
rect 40290 37774 40292 37826
rect 40236 37772 40292 37774
rect 41244 39564 41300 39620
rect 40460 37938 40516 37940
rect 40460 37886 40462 37938
rect 40462 37886 40514 37938
rect 40514 37886 40516 37938
rect 40460 37884 40516 37886
rect 41020 39116 41076 39172
rect 40796 38892 40852 38948
rect 40908 38050 40964 38052
rect 40908 37998 40910 38050
rect 40910 37998 40962 38050
rect 40962 37998 40964 38050
rect 40908 37996 40964 37998
rect 40684 37772 40740 37828
rect 41356 40124 41412 40180
rect 43596 42082 43652 42084
rect 43596 42030 43598 42082
rect 43598 42030 43650 42082
rect 43650 42030 43652 42082
rect 43596 42028 43652 42030
rect 43036 41970 43092 41972
rect 43036 41918 43038 41970
rect 43038 41918 43090 41970
rect 43090 41918 43092 41970
rect 43036 41916 43092 41918
rect 42028 41074 42084 41076
rect 42028 41022 42030 41074
rect 42030 41022 42082 41074
rect 42082 41022 42084 41074
rect 42028 41020 42084 41022
rect 41916 40124 41972 40180
rect 43148 39676 43204 39732
rect 41916 38892 41972 38948
rect 44492 41916 44548 41972
rect 44044 40572 44100 40628
rect 43820 40290 43876 40292
rect 43820 40238 43822 40290
rect 43822 40238 43874 40290
rect 43874 40238 43876 40290
rect 43820 40236 43876 40238
rect 41804 37996 41860 38052
rect 42700 37996 42756 38052
rect 40796 37212 40852 37268
rect 40012 35084 40068 35140
rect 39676 33180 39732 33236
rect 39452 32620 39508 32676
rect 39564 31948 39620 32004
rect 38444 31554 38500 31556
rect 38444 31502 38446 31554
rect 38446 31502 38498 31554
rect 38498 31502 38500 31554
rect 38444 31500 38500 31502
rect 38668 30882 38724 30884
rect 38668 30830 38670 30882
rect 38670 30830 38722 30882
rect 38722 30830 38724 30882
rect 38668 30828 38724 30830
rect 39228 30994 39284 30996
rect 39228 30942 39230 30994
rect 39230 30942 39282 30994
rect 39282 30942 39284 30994
rect 39228 30940 39284 30942
rect 39340 31052 39396 31108
rect 39900 34188 39956 34244
rect 40012 34636 40068 34692
rect 40348 35308 40404 35364
rect 40460 34860 40516 34916
rect 41132 35644 41188 35700
rect 40348 34076 40404 34132
rect 39564 31724 39620 31780
rect 40124 32732 40180 32788
rect 41580 37266 41636 37268
rect 41580 37214 41582 37266
rect 41582 37214 41634 37266
rect 41634 37214 41636 37266
rect 41580 37212 41636 37214
rect 41356 35532 41412 35588
rect 41244 35308 41300 35364
rect 41804 34860 41860 34916
rect 41804 34354 41860 34356
rect 41804 34302 41806 34354
rect 41806 34302 41858 34354
rect 41858 34302 41860 34354
rect 41804 34300 41860 34302
rect 40908 34242 40964 34244
rect 40908 34190 40910 34242
rect 40910 34190 40962 34242
rect 40962 34190 40964 34242
rect 40908 34188 40964 34190
rect 41244 34242 41300 34244
rect 41244 34190 41246 34242
rect 41246 34190 41298 34242
rect 41298 34190 41300 34242
rect 41244 34188 41300 34190
rect 42140 34130 42196 34132
rect 42140 34078 42142 34130
rect 42142 34078 42194 34130
rect 42194 34078 42196 34130
rect 42140 34076 42196 34078
rect 42588 37826 42644 37828
rect 42588 37774 42590 37826
rect 42590 37774 42642 37826
rect 42642 37774 42644 37826
rect 42588 37772 42644 37774
rect 43596 38050 43652 38052
rect 43596 37998 43598 38050
rect 43598 37998 43650 38050
rect 43650 37998 43652 38050
rect 43596 37996 43652 37998
rect 43036 37938 43092 37940
rect 43036 37886 43038 37938
rect 43038 37886 43090 37938
rect 43090 37886 43092 37938
rect 43036 37884 43092 37886
rect 43932 39618 43988 39620
rect 43932 39566 43934 39618
rect 43934 39566 43986 39618
rect 43986 39566 43988 39618
rect 43932 39564 43988 39566
rect 44156 40124 44212 40180
rect 43484 37042 43540 37044
rect 43484 36990 43486 37042
rect 43486 36990 43538 37042
rect 43538 36990 43540 37042
rect 43484 36988 43540 36990
rect 43148 35532 43204 35588
rect 42588 34242 42644 34244
rect 42588 34190 42590 34242
rect 42590 34190 42642 34242
rect 42642 34190 42644 34242
rect 42588 34188 42644 34190
rect 43820 35698 43876 35700
rect 43820 35646 43822 35698
rect 43822 35646 43874 35698
rect 43874 35646 43876 35698
rect 43820 35644 43876 35646
rect 43932 36204 43988 36260
rect 43820 34018 43876 34020
rect 43820 33966 43822 34018
rect 43822 33966 43874 34018
rect 43874 33966 43876 34018
rect 43820 33964 43876 33966
rect 40012 32674 40068 32676
rect 40012 32622 40014 32674
rect 40014 32622 40066 32674
rect 40066 32622 40068 32674
rect 40012 32620 40068 32622
rect 40348 32786 40404 32788
rect 40348 32734 40350 32786
rect 40350 32734 40402 32786
rect 40402 32734 40404 32786
rect 40348 32732 40404 32734
rect 39676 31276 39732 31332
rect 40236 32284 40292 32340
rect 40572 33234 40628 33236
rect 40572 33182 40574 33234
rect 40574 33182 40626 33234
rect 40626 33182 40628 33234
rect 40572 33180 40628 33182
rect 41356 32732 41412 32788
rect 40460 32060 40516 32116
rect 41020 32562 41076 32564
rect 41020 32510 41022 32562
rect 41022 32510 41074 32562
rect 41074 32510 41076 32562
rect 41020 32508 41076 32510
rect 43148 33122 43204 33124
rect 43148 33070 43150 33122
rect 43150 33070 43202 33122
rect 43202 33070 43204 33122
rect 43148 33068 43204 33070
rect 42924 32786 42980 32788
rect 42924 32734 42926 32786
rect 42926 32734 42978 32786
rect 42978 32734 42980 32786
rect 42924 32732 42980 32734
rect 41132 32338 41188 32340
rect 41132 32286 41134 32338
rect 41134 32286 41186 32338
rect 41186 32286 41188 32338
rect 41132 32284 41188 32286
rect 40348 31778 40404 31780
rect 40348 31726 40350 31778
rect 40350 31726 40402 31778
rect 40402 31726 40404 31778
rect 40348 31724 40404 31726
rect 40124 31276 40180 31332
rect 39900 31106 39956 31108
rect 39900 31054 39902 31106
rect 39902 31054 39954 31106
rect 39954 31054 39956 31106
rect 39900 31052 39956 31054
rect 41020 31554 41076 31556
rect 41020 31502 41022 31554
rect 41022 31502 41074 31554
rect 41074 31502 41076 31554
rect 41020 31500 41076 31502
rect 40572 31052 40628 31108
rect 41020 30940 41076 30996
rect 39788 30828 39844 30884
rect 40908 30882 40964 30884
rect 40908 30830 40910 30882
rect 40910 30830 40962 30882
rect 40962 30830 40964 30882
rect 40908 30828 40964 30830
rect 39452 30268 39508 30324
rect 39116 30044 39172 30100
rect 37996 29932 38052 29988
rect 37996 29260 38052 29316
rect 38780 29986 38836 29988
rect 38780 29934 38782 29986
rect 38782 29934 38834 29986
rect 38834 29934 38836 29986
rect 38780 29932 38836 29934
rect 34748 29148 34804 29204
rect 33740 28642 33796 28644
rect 33740 28590 33742 28642
rect 33742 28590 33794 28642
rect 33794 28590 33796 28642
rect 33740 28588 33796 28590
rect 34300 28642 34356 28644
rect 34300 28590 34302 28642
rect 34302 28590 34354 28642
rect 34354 28590 34356 28642
rect 34300 28588 34356 28590
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 40012 29372 40068 29428
rect 40908 29426 40964 29428
rect 40908 29374 40910 29426
rect 40910 29374 40962 29426
rect 40962 29374 40964 29426
rect 40908 29372 40964 29374
rect 41244 30156 41300 30212
rect 41804 30828 41860 30884
rect 41916 30268 41972 30324
rect 42476 32562 42532 32564
rect 42476 32510 42478 32562
rect 42478 32510 42530 32562
rect 42530 32510 42532 32562
rect 42476 32508 42532 32510
rect 42028 30044 42084 30100
rect 42588 30210 42644 30212
rect 42588 30158 42590 30210
rect 42590 30158 42642 30210
rect 42642 30158 42644 30210
rect 42588 30156 42644 30158
rect 43596 32620 43652 32676
rect 43708 30994 43764 30996
rect 43708 30942 43710 30994
rect 43710 30942 43762 30994
rect 43762 30942 43764 30994
rect 43708 30940 43764 30942
rect 43148 30380 43204 30436
rect 42140 29372 42196 29428
rect 43484 30044 43540 30100
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35084 27186 35140 27188
rect 35084 27134 35086 27186
rect 35086 27134 35138 27186
rect 35138 27134 35140 27186
rect 35084 27132 35140 27134
rect 37100 27186 37156 27188
rect 37100 27134 37102 27186
rect 37102 27134 37154 27186
rect 37154 27134 37156 27186
rect 37100 27132 37156 27134
rect 34748 26962 34804 26964
rect 34748 26910 34750 26962
rect 34750 26910 34802 26962
rect 34802 26910 34804 26962
rect 34748 26908 34804 26910
rect 35644 26962 35700 26964
rect 35644 26910 35646 26962
rect 35646 26910 35698 26962
rect 35698 26910 35700 26962
rect 35644 26908 35700 26910
rect 34076 26178 34132 26180
rect 34076 26126 34078 26178
rect 34078 26126 34130 26178
rect 34130 26126 34132 26178
rect 34076 26124 34132 26126
rect 33068 24668 33124 24724
rect 33068 23324 33124 23380
rect 34636 25564 34692 25620
rect 33740 24610 33796 24612
rect 33740 24558 33742 24610
rect 33742 24558 33794 24610
rect 33794 24558 33796 24610
rect 33740 24556 33796 24558
rect 34188 23548 34244 23604
rect 33404 23212 33460 23268
rect 33964 23212 34020 23268
rect 33068 22482 33124 22484
rect 33068 22430 33070 22482
rect 33070 22430 33122 22482
rect 33122 22430 33124 22482
rect 33068 22428 33124 22430
rect 34076 22316 34132 22372
rect 34412 22652 34468 22708
rect 35084 26124 35140 26180
rect 34972 24668 35028 24724
rect 34524 22428 34580 22484
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35868 24892 35924 24948
rect 36092 24668 36148 24724
rect 36204 26908 36260 26964
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 23938 35252 23940
rect 35196 23886 35198 23938
rect 35198 23886 35250 23938
rect 35250 23886 35252 23938
rect 35196 23884 35252 23886
rect 37996 26348 38052 26404
rect 37884 26178 37940 26180
rect 37884 26126 37886 26178
rect 37886 26126 37938 26178
rect 37938 26126 37940 26178
rect 37884 26124 37940 26126
rect 35532 23714 35588 23716
rect 35532 23662 35534 23714
rect 35534 23662 35586 23714
rect 35586 23662 35588 23714
rect 35532 23660 35588 23662
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35644 22540 35700 22596
rect 35420 22370 35476 22372
rect 35420 22318 35422 22370
rect 35422 22318 35474 22370
rect 35474 22318 35476 22370
rect 35420 22316 35476 22318
rect 35644 22370 35700 22372
rect 35644 22318 35646 22370
rect 35646 22318 35698 22370
rect 35698 22318 35700 22370
rect 35644 22316 35700 22318
rect 34412 22258 34468 22260
rect 34412 22206 34414 22258
rect 34414 22206 34466 22258
rect 34466 22206 34468 22258
rect 34412 22204 34468 22206
rect 34188 21868 34244 21924
rect 35084 21980 35140 22036
rect 35196 22092 35252 22148
rect 34748 21644 34804 21700
rect 35196 21644 35252 21700
rect 35644 21644 35700 21700
rect 34188 20860 34244 20916
rect 34300 20972 34356 21028
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34188 20690 34244 20692
rect 34188 20638 34190 20690
rect 34190 20638 34242 20690
rect 34242 20638 34244 20690
rect 34188 20636 34244 20638
rect 32844 19964 32900 20020
rect 32620 18172 32676 18228
rect 32508 17442 32564 17444
rect 32508 17390 32510 17442
rect 32510 17390 32562 17442
rect 32562 17390 32564 17442
rect 32508 17388 32564 17390
rect 31948 16268 32004 16324
rect 31276 13916 31332 13972
rect 31276 13746 31332 13748
rect 31276 13694 31278 13746
rect 31278 13694 31330 13746
rect 31330 13694 31332 13746
rect 31276 13692 31332 13694
rect 30940 12290 30996 12292
rect 30940 12238 30942 12290
rect 30942 12238 30994 12290
rect 30994 12238 30996 12290
rect 30940 12236 30996 12238
rect 31500 13858 31556 13860
rect 31500 13806 31502 13858
rect 31502 13806 31554 13858
rect 31554 13806 31556 13858
rect 31500 13804 31556 13806
rect 32060 15090 32116 15092
rect 32060 15038 32062 15090
rect 32062 15038 32114 15090
rect 32114 15038 32116 15090
rect 32060 15036 32116 15038
rect 31836 13916 31892 13972
rect 32060 13858 32116 13860
rect 32060 13806 32062 13858
rect 32062 13806 32114 13858
rect 32114 13806 32116 13858
rect 32060 13804 32116 13806
rect 32620 13804 32676 13860
rect 31724 13692 31780 13748
rect 31948 13692 32004 13748
rect 31500 12738 31556 12740
rect 31500 12686 31502 12738
rect 31502 12686 31554 12738
rect 31554 12686 31556 12738
rect 31500 12684 31556 12686
rect 30268 11564 30324 11620
rect 29148 10556 29204 10612
rect 29932 10444 29988 10500
rect 31052 10722 31108 10724
rect 31052 10670 31054 10722
rect 31054 10670 31106 10722
rect 31106 10670 31108 10722
rect 31052 10668 31108 10670
rect 30492 9996 30548 10052
rect 28476 8876 28532 8932
rect 25788 8092 25844 8148
rect 28812 7868 28868 7924
rect 25900 6748 25956 6804
rect 24332 6466 24388 6468
rect 24332 6414 24334 6466
rect 24334 6414 24386 6466
rect 24386 6414 24388 6466
rect 24332 6412 24388 6414
rect 22764 6076 22820 6132
rect 23772 6130 23828 6132
rect 23772 6078 23774 6130
rect 23774 6078 23826 6130
rect 23826 6078 23828 6130
rect 23772 6076 23828 6078
rect 22428 5964 22484 6020
rect 21644 5234 21700 5236
rect 21644 5182 21646 5234
rect 21646 5182 21698 5234
rect 21698 5182 21700 5234
rect 21644 5180 21700 5182
rect 20300 4898 20356 4900
rect 20300 4846 20302 4898
rect 20302 4846 20354 4898
rect 20354 4846 20356 4898
rect 20300 4844 20356 4846
rect 21084 4844 21140 4900
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19292 4396 19348 4452
rect 19852 4396 19908 4452
rect 19516 4060 19572 4116
rect 12684 3500 12740 3556
rect 14028 3554 14084 3556
rect 14028 3502 14030 3554
rect 14030 3502 14082 3554
rect 14082 3502 14084 3554
rect 14028 3500 14084 3502
rect 19516 3500 19572 3556
rect 22204 5122 22260 5124
rect 22204 5070 22206 5122
rect 22206 5070 22258 5122
rect 22258 5070 22260 5122
rect 22204 5068 22260 5070
rect 21644 4284 21700 4340
rect 22316 4338 22372 4340
rect 22316 4286 22318 4338
rect 22318 4286 22370 4338
rect 22370 4286 22372 4338
rect 22316 4284 22372 4286
rect 21420 4226 21476 4228
rect 21420 4174 21422 4226
rect 21422 4174 21474 4226
rect 21474 4174 21476 4226
rect 21420 4172 21476 4174
rect 25228 6018 25284 6020
rect 25228 5966 25230 6018
rect 25230 5966 25282 6018
rect 25282 5966 25284 6018
rect 25228 5964 25284 5966
rect 24332 5852 24388 5908
rect 23212 4898 23268 4900
rect 23212 4846 23214 4898
rect 23214 4846 23266 4898
rect 23266 4846 23268 4898
rect 23212 4844 23268 4846
rect 24444 5068 24500 5124
rect 26908 6412 26964 6468
rect 28140 6466 28196 6468
rect 28140 6414 28142 6466
rect 28142 6414 28194 6466
rect 28194 6414 28196 6466
rect 28140 6412 28196 6414
rect 30604 9548 30660 9604
rect 29820 8930 29876 8932
rect 29820 8878 29822 8930
rect 29822 8878 29874 8930
rect 29874 8878 29876 8930
rect 29820 8876 29876 8878
rect 29260 8370 29316 8372
rect 29260 8318 29262 8370
rect 29262 8318 29314 8370
rect 29314 8318 29316 8370
rect 29260 8316 29316 8318
rect 30940 10498 30996 10500
rect 30940 10446 30942 10498
rect 30942 10446 30994 10498
rect 30994 10446 30996 10498
rect 30940 10444 30996 10446
rect 33404 20076 33460 20132
rect 33404 19404 33460 19460
rect 33292 19234 33348 19236
rect 33292 19182 33294 19234
rect 33294 19182 33346 19234
rect 33346 19182 33348 19234
rect 33292 19180 33348 19182
rect 33068 18450 33124 18452
rect 33068 18398 33070 18450
rect 33070 18398 33122 18450
rect 33122 18398 33124 18450
rect 33068 18396 33124 18398
rect 33628 18396 33684 18452
rect 33068 17500 33124 17556
rect 33404 17388 33460 17444
rect 33068 16268 33124 16324
rect 33964 20018 34020 20020
rect 33964 19966 33966 20018
rect 33966 19966 34018 20018
rect 34018 19966 34020 20018
rect 33964 19964 34020 19966
rect 34076 18284 34132 18340
rect 34972 20636 35028 20692
rect 35196 20690 35252 20692
rect 35196 20638 35198 20690
rect 35198 20638 35250 20690
rect 35250 20638 35252 20690
rect 35196 20636 35252 20638
rect 35420 20578 35476 20580
rect 35420 20526 35422 20578
rect 35422 20526 35474 20578
rect 35474 20526 35476 20578
rect 35420 20524 35476 20526
rect 35196 20076 35252 20132
rect 35420 20018 35476 20020
rect 35420 19966 35422 20018
rect 35422 19966 35474 20018
rect 35474 19966 35476 20018
rect 35420 19964 35476 19966
rect 34972 19906 35028 19908
rect 34972 19854 34974 19906
rect 34974 19854 35026 19906
rect 35026 19854 35028 19906
rect 34972 19852 35028 19854
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34748 19180 34804 19236
rect 35644 19068 35700 19124
rect 34636 18450 34692 18452
rect 34636 18398 34638 18450
rect 34638 18398 34690 18450
rect 34690 18398 34692 18450
rect 34636 18396 34692 18398
rect 35308 18450 35364 18452
rect 35308 18398 35310 18450
rect 35310 18398 35362 18450
rect 35362 18398 35364 18450
rect 35308 18396 35364 18398
rect 34300 18284 34356 18340
rect 33852 17724 33908 17780
rect 34300 17554 34356 17556
rect 34300 17502 34302 17554
rect 34302 17502 34354 17554
rect 34354 17502 34356 17554
rect 34300 17500 34356 17502
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35084 17500 35140 17556
rect 35532 16828 35588 16884
rect 34300 16716 34356 16772
rect 36204 23548 36260 23604
rect 37212 24892 37268 24948
rect 37884 25228 37940 25284
rect 38892 26348 38948 26404
rect 41804 27692 41860 27748
rect 38444 25228 38500 25284
rect 38332 24668 38388 24724
rect 36988 23548 37044 23604
rect 35980 23324 36036 23380
rect 35868 23100 35924 23156
rect 36092 23212 36148 23268
rect 36540 23266 36596 23268
rect 36540 23214 36542 23266
rect 36542 23214 36594 23266
rect 36594 23214 36596 23266
rect 36540 23212 36596 23214
rect 36092 22652 36148 22708
rect 35980 22316 36036 22372
rect 35868 21756 35924 21812
rect 36764 23154 36820 23156
rect 36764 23102 36766 23154
rect 36766 23102 36818 23154
rect 36818 23102 36820 23154
rect 36764 23100 36820 23102
rect 36988 23324 37044 23380
rect 37884 23266 37940 23268
rect 37884 23214 37886 23266
rect 37886 23214 37938 23266
rect 37938 23214 37940 23266
rect 37884 23212 37940 23214
rect 36428 21868 36484 21924
rect 37772 23154 37828 23156
rect 37772 23102 37774 23154
rect 37774 23102 37826 23154
rect 37826 23102 37828 23154
rect 37772 23100 37828 23102
rect 36540 21698 36596 21700
rect 36540 21646 36542 21698
rect 36542 21646 36594 21698
rect 36594 21646 36596 21698
rect 36540 21644 36596 21646
rect 35868 21026 35924 21028
rect 35868 20974 35870 21026
rect 35870 20974 35922 21026
rect 35922 20974 35924 21026
rect 35868 20972 35924 20974
rect 35980 20188 36036 20244
rect 36652 21586 36708 21588
rect 36652 21534 36654 21586
rect 36654 21534 36706 21586
rect 36706 21534 36708 21586
rect 36652 21532 36708 21534
rect 36540 21420 36596 21476
rect 35868 17612 35924 17668
rect 35756 16716 35812 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 32956 15708 33012 15764
rect 34300 15820 34356 15876
rect 35532 15708 35588 15764
rect 34076 15036 34132 15092
rect 33068 13916 33124 13972
rect 33404 13858 33460 13860
rect 33404 13806 33406 13858
rect 33406 13806 33458 13858
rect 33458 13806 33460 13858
rect 33404 13804 33460 13806
rect 32956 13692 33012 13748
rect 33180 13468 33236 13524
rect 32844 12908 32900 12964
rect 32396 12066 32452 12068
rect 32396 12014 32398 12066
rect 32398 12014 32450 12066
rect 32450 12014 32452 12066
rect 32396 12012 32452 12014
rect 33516 12908 33572 12964
rect 32956 11564 33012 11620
rect 32844 11452 32900 11508
rect 32620 11228 32676 11284
rect 32284 10780 32340 10836
rect 31724 10722 31780 10724
rect 31724 10670 31726 10722
rect 31726 10670 31778 10722
rect 31778 10670 31780 10722
rect 31724 10668 31780 10670
rect 31388 9548 31444 9604
rect 30940 9154 30996 9156
rect 30940 9102 30942 9154
rect 30942 9102 30994 9154
rect 30994 9102 30996 9154
rect 30940 9100 30996 9102
rect 30044 8316 30100 8372
rect 30380 7644 30436 7700
rect 28588 6802 28644 6804
rect 28588 6750 28590 6802
rect 28590 6750 28642 6802
rect 28642 6750 28644 6802
rect 28588 6748 28644 6750
rect 31052 8034 31108 8036
rect 31052 7982 31054 8034
rect 31054 7982 31106 8034
rect 31106 7982 31108 8034
rect 31052 7980 31108 7982
rect 31724 9100 31780 9156
rect 32508 9602 32564 9604
rect 32508 9550 32510 9602
rect 32510 9550 32562 9602
rect 32562 9550 32564 9602
rect 32508 9548 32564 9550
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34188 13858 34244 13860
rect 34188 13806 34190 13858
rect 34190 13806 34242 13858
rect 34242 13806 34244 13858
rect 34188 13804 34244 13806
rect 35084 13916 35140 13972
rect 36428 20188 36484 20244
rect 36540 20018 36596 20020
rect 36540 19966 36542 20018
rect 36542 19966 36594 20018
rect 36594 19966 36596 20018
rect 36540 19964 36596 19966
rect 36428 19068 36484 19124
rect 36540 18450 36596 18452
rect 36540 18398 36542 18450
rect 36542 18398 36594 18450
rect 36594 18398 36596 18450
rect 36540 18396 36596 18398
rect 36204 18172 36260 18228
rect 36316 17500 36372 17556
rect 36876 22652 36932 22708
rect 37100 22540 37156 22596
rect 37884 22316 37940 22372
rect 38892 23436 38948 23492
rect 37212 22258 37268 22260
rect 37212 22206 37214 22258
rect 37214 22206 37266 22258
rect 37266 22206 37268 22258
rect 37212 22204 37268 22206
rect 37324 22146 37380 22148
rect 37324 22094 37326 22146
rect 37326 22094 37378 22146
rect 37378 22094 37380 22146
rect 37324 22092 37380 22094
rect 38556 22594 38612 22596
rect 38556 22542 38558 22594
rect 38558 22542 38610 22594
rect 38610 22542 38612 22594
rect 38556 22540 38612 22542
rect 38556 21756 38612 21812
rect 37548 20972 37604 21028
rect 38108 21532 38164 21588
rect 37100 20914 37156 20916
rect 37100 20862 37102 20914
rect 37102 20862 37154 20914
rect 37154 20862 37156 20914
rect 37100 20860 37156 20862
rect 37212 20690 37268 20692
rect 37212 20638 37214 20690
rect 37214 20638 37266 20690
rect 37266 20638 37268 20690
rect 37212 20636 37268 20638
rect 37100 20578 37156 20580
rect 37100 20526 37102 20578
rect 37102 20526 37154 20578
rect 37154 20526 37156 20578
rect 37100 20524 37156 20526
rect 36876 19964 36932 20020
rect 37100 19964 37156 20020
rect 37100 18172 37156 18228
rect 37436 20076 37492 20132
rect 39116 20860 39172 20916
rect 39452 24668 39508 24724
rect 39788 23436 39844 23492
rect 39900 23212 39956 23268
rect 39452 22370 39508 22372
rect 39452 22318 39454 22370
rect 39454 22318 39506 22370
rect 39506 22318 39508 22370
rect 39452 22316 39508 22318
rect 39788 21810 39844 21812
rect 39788 21758 39790 21810
rect 39790 21758 39842 21810
rect 39842 21758 39844 21810
rect 39788 21756 39844 21758
rect 38108 19964 38164 20020
rect 37660 19852 37716 19908
rect 37660 19068 37716 19124
rect 37212 18284 37268 18340
rect 37548 17778 37604 17780
rect 37548 17726 37550 17778
rect 37550 17726 37602 17778
rect 37602 17726 37604 17778
rect 37548 17724 37604 17726
rect 38892 17666 38948 17668
rect 38892 17614 38894 17666
rect 38894 17614 38946 17666
rect 38946 17614 38948 17666
rect 38892 17612 38948 17614
rect 36988 17554 37044 17556
rect 36988 17502 36990 17554
rect 36990 17502 37042 17554
rect 37042 17502 37044 17554
rect 36988 17500 37044 17502
rect 38892 17052 38948 17108
rect 36540 16716 36596 16772
rect 40684 23100 40740 23156
rect 40348 23042 40404 23044
rect 40348 22990 40350 23042
rect 40350 22990 40402 23042
rect 40402 22990 40404 23042
rect 40348 22988 40404 22990
rect 40684 22428 40740 22484
rect 39116 20076 39172 20132
rect 39676 20018 39732 20020
rect 39676 19966 39678 20018
rect 39678 19966 39730 20018
rect 39730 19966 39732 20018
rect 39676 19964 39732 19966
rect 40012 20130 40068 20132
rect 40012 20078 40014 20130
rect 40014 20078 40066 20130
rect 40066 20078 40068 20130
rect 40012 20076 40068 20078
rect 40348 20130 40404 20132
rect 40348 20078 40350 20130
rect 40350 20078 40402 20130
rect 40402 20078 40404 20130
rect 40348 20076 40404 20078
rect 40236 19292 40292 19348
rect 40684 19234 40740 19236
rect 40684 19182 40686 19234
rect 40686 19182 40738 19234
rect 40738 19182 40740 19234
rect 40684 19180 40740 19182
rect 40236 19122 40292 19124
rect 40236 19070 40238 19122
rect 40238 19070 40290 19122
rect 40290 19070 40292 19122
rect 40236 19068 40292 19070
rect 43148 27746 43204 27748
rect 43148 27694 43150 27746
rect 43150 27694 43202 27746
rect 43202 27694 43204 27746
rect 43148 27692 43204 27694
rect 43596 27746 43652 27748
rect 43596 27694 43598 27746
rect 43598 27694 43650 27746
rect 43650 27694 43652 27746
rect 43596 27692 43652 27694
rect 43148 26908 43204 26964
rect 44492 36204 44548 36260
rect 44492 33964 44548 34020
rect 44156 27692 44212 27748
rect 44268 26908 44324 26964
rect 43820 26012 43876 26068
rect 41468 25618 41524 25620
rect 41468 25566 41470 25618
rect 41470 25566 41522 25618
rect 41522 25566 41524 25618
rect 41468 25564 41524 25566
rect 44044 25564 44100 25620
rect 41468 24722 41524 24724
rect 41468 24670 41470 24722
rect 41470 24670 41522 24722
rect 41522 24670 41524 24722
rect 41468 24668 41524 24670
rect 41580 23154 41636 23156
rect 41580 23102 41582 23154
rect 41582 23102 41634 23154
rect 41634 23102 41636 23154
rect 41580 23100 41636 23102
rect 41020 21308 41076 21364
rect 41692 23042 41748 23044
rect 41692 22990 41694 23042
rect 41694 22990 41746 23042
rect 41746 22990 41748 23042
rect 41692 22988 41748 22990
rect 42812 23154 42868 23156
rect 42812 23102 42814 23154
rect 42814 23102 42866 23154
rect 42866 23102 42868 23154
rect 42812 23100 42868 23102
rect 42364 22482 42420 22484
rect 42364 22430 42366 22482
rect 42366 22430 42418 22482
rect 42418 22430 42420 22482
rect 42364 22428 42420 22430
rect 41468 20914 41524 20916
rect 41468 20862 41470 20914
rect 41470 20862 41522 20914
rect 41522 20862 41524 20914
rect 41468 20860 41524 20862
rect 41132 20578 41188 20580
rect 41132 20526 41134 20578
rect 41134 20526 41186 20578
rect 41186 20526 41188 20578
rect 41132 20524 41188 20526
rect 40908 20130 40964 20132
rect 40908 20078 40910 20130
rect 40910 20078 40962 20130
rect 40962 20078 40964 20130
rect 40908 20076 40964 20078
rect 42252 21362 42308 21364
rect 42252 21310 42254 21362
rect 42254 21310 42306 21362
rect 42306 21310 42308 21362
rect 42252 21308 42308 21310
rect 43372 21308 43428 21364
rect 43260 20578 43316 20580
rect 43260 20526 43262 20578
rect 43262 20526 43314 20578
rect 43314 20526 43316 20578
rect 43260 20524 43316 20526
rect 42028 19964 42084 20020
rect 40796 18844 40852 18900
rect 41244 19180 41300 19236
rect 40124 18338 40180 18340
rect 40124 18286 40126 18338
rect 40126 18286 40178 18338
rect 40178 18286 40180 18338
rect 40124 18284 40180 18286
rect 40684 18284 40740 18340
rect 36540 15148 36596 15204
rect 35420 13522 35476 13524
rect 35420 13470 35422 13522
rect 35422 13470 35474 13522
rect 35474 13470 35476 13522
rect 35420 13468 35476 13470
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 34524 13132 34580 13188
rect 39228 15202 39284 15204
rect 39228 15150 39230 15202
rect 39230 15150 39282 15202
rect 39282 15150 39284 15202
rect 39228 15148 39284 15150
rect 39116 13970 39172 13972
rect 39116 13918 39118 13970
rect 39118 13918 39170 13970
rect 39170 13918 39172 13970
rect 39116 13916 39172 13918
rect 36652 13244 36708 13300
rect 37436 13244 37492 13300
rect 36988 13186 37044 13188
rect 36988 13134 36990 13186
rect 36990 13134 37042 13186
rect 37042 13134 37044 13186
rect 36988 13132 37044 13134
rect 36428 12796 36484 12852
rect 33964 12460 34020 12516
rect 33852 12066 33908 12068
rect 33852 12014 33854 12066
rect 33854 12014 33906 12066
rect 33906 12014 33908 12066
rect 33852 12012 33908 12014
rect 33852 11506 33908 11508
rect 33852 11454 33854 11506
rect 33854 11454 33906 11506
rect 33906 11454 33908 11506
rect 33852 11452 33908 11454
rect 33516 11228 33572 11284
rect 36540 12460 36596 12516
rect 34076 12348 34132 12404
rect 36316 12348 36372 12404
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 36092 11788 36148 11844
rect 35980 11506 36036 11508
rect 35980 11454 35982 11506
rect 35982 11454 36034 11506
rect 36034 11454 36036 11506
rect 35980 11452 36036 11454
rect 35532 11340 35588 11396
rect 31388 7196 31444 7252
rect 31948 7644 32004 7700
rect 31948 7196 32004 7252
rect 32396 7698 32452 7700
rect 32396 7646 32398 7698
rect 32398 7646 32450 7698
rect 32450 7646 32452 7698
rect 32396 7644 32452 7646
rect 33292 7698 33348 7700
rect 33292 7646 33294 7698
rect 33294 7646 33346 7698
rect 33346 7646 33348 7698
rect 33292 7644 33348 7646
rect 32620 7586 32676 7588
rect 32620 7534 32622 7586
rect 32622 7534 32674 7586
rect 32674 7534 32676 7586
rect 32620 7532 32676 7534
rect 32956 7308 33012 7364
rect 29148 6412 29204 6468
rect 32396 6636 32452 6692
rect 32620 6412 32676 6468
rect 32620 6130 32676 6132
rect 32620 6078 32622 6130
rect 32622 6078 32674 6130
rect 32674 6078 32676 6130
rect 32620 6076 32676 6078
rect 34524 9996 34580 10052
rect 34860 10780 34916 10836
rect 35308 10722 35364 10724
rect 35308 10670 35310 10722
rect 35310 10670 35362 10722
rect 35362 10670 35364 10722
rect 35308 10668 35364 10670
rect 36764 13020 36820 13076
rect 37100 12850 37156 12852
rect 37100 12798 37102 12850
rect 37102 12798 37154 12850
rect 37154 12798 37156 12850
rect 37100 12796 37156 12798
rect 36764 11340 36820 11396
rect 36316 10892 36372 10948
rect 34748 10444 34804 10500
rect 35084 10610 35140 10612
rect 35084 10558 35086 10610
rect 35086 10558 35138 10610
rect 35138 10558 35140 10610
rect 35084 10556 35140 10558
rect 35532 10332 35588 10388
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34524 9436 34580 9492
rect 35084 9266 35140 9268
rect 35084 9214 35086 9266
rect 35086 9214 35138 9266
rect 35138 9214 35140 9266
rect 35084 9212 35140 9214
rect 35980 9772 36036 9828
rect 36316 9996 36372 10052
rect 34300 9100 34356 9156
rect 34188 8988 34244 9044
rect 34076 7980 34132 8036
rect 33516 7586 33572 7588
rect 33516 7534 33518 7586
rect 33518 7534 33570 7586
rect 33570 7534 33572 7586
rect 33516 7532 33572 7534
rect 34076 7420 34132 7476
rect 35868 9100 35924 9156
rect 35756 8764 35812 8820
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 34748 7980 34804 8036
rect 36316 8652 36372 8708
rect 36540 10668 36596 10724
rect 37548 13074 37604 13076
rect 37548 13022 37550 13074
rect 37550 13022 37602 13074
rect 37602 13022 37604 13074
rect 37548 13020 37604 13022
rect 38220 13020 38276 13076
rect 38780 12402 38836 12404
rect 38780 12350 38782 12402
rect 38782 12350 38834 12402
rect 38834 12350 38836 12402
rect 38780 12348 38836 12350
rect 38892 12684 38948 12740
rect 36988 10610 37044 10612
rect 36988 10558 36990 10610
rect 36990 10558 37042 10610
rect 37042 10558 37044 10610
rect 36988 10556 37044 10558
rect 37772 11394 37828 11396
rect 37772 11342 37774 11394
rect 37774 11342 37826 11394
rect 37826 11342 37828 11394
rect 37772 11340 37828 11342
rect 38220 11618 38276 11620
rect 38220 11566 38222 11618
rect 38222 11566 38274 11618
rect 38274 11566 38276 11618
rect 38220 11564 38276 11566
rect 38108 11506 38164 11508
rect 38108 11454 38110 11506
rect 38110 11454 38162 11506
rect 38162 11454 38164 11506
rect 38108 11452 38164 11454
rect 37548 10780 37604 10836
rect 38556 11564 38612 11620
rect 38332 11340 38388 11396
rect 37436 10722 37492 10724
rect 37436 10670 37438 10722
rect 37438 10670 37490 10722
rect 37490 10670 37492 10722
rect 37436 10668 37492 10670
rect 36652 9042 36708 9044
rect 36652 8990 36654 9042
rect 36654 8990 36706 9042
rect 36706 8990 36708 9042
rect 36652 8988 36708 8990
rect 37212 9212 37268 9268
rect 37212 8876 37268 8932
rect 36988 8764 37044 8820
rect 34860 7868 34916 7924
rect 33964 7362 34020 7364
rect 33964 7310 33966 7362
rect 33966 7310 34018 7362
rect 34018 7310 34020 7362
rect 33964 7308 34020 7310
rect 33292 6690 33348 6692
rect 33292 6638 33294 6690
rect 33294 6638 33346 6690
rect 33346 6638 33348 6690
rect 33292 6636 33348 6638
rect 33180 6524 33236 6580
rect 33292 6130 33348 6132
rect 33292 6078 33294 6130
rect 33294 6078 33346 6130
rect 33346 6078 33348 6130
rect 33292 6076 33348 6078
rect 28028 5906 28084 5908
rect 28028 5854 28030 5906
rect 28030 5854 28082 5906
rect 28082 5854 28084 5906
rect 28028 5852 28084 5854
rect 25228 4844 25284 4900
rect 24332 4396 24388 4452
rect 22988 4226 23044 4228
rect 22988 4174 22990 4226
rect 22990 4174 23042 4226
rect 23042 4174 23044 4226
rect 22988 4172 23044 4174
rect 24668 4338 24724 4340
rect 24668 4286 24670 4338
rect 24670 4286 24722 4338
rect 24722 4286 24724 4338
rect 24668 4284 24724 4286
rect 25452 4338 25508 4340
rect 25452 4286 25454 4338
rect 25454 4286 25506 4338
rect 25506 4286 25508 4338
rect 25452 4284 25508 4286
rect 28140 4226 28196 4228
rect 28140 4174 28142 4226
rect 28142 4174 28194 4226
rect 28194 4174 28196 4226
rect 28140 4172 28196 4174
rect 28588 4172 28644 4228
rect 23772 4060 23828 4116
rect 29484 5852 29540 5908
rect 31612 6018 31668 6020
rect 31612 5966 31614 6018
rect 31614 5966 31666 6018
rect 31666 5966 31668 6018
rect 31612 5964 31668 5966
rect 34300 6748 34356 6804
rect 34076 6578 34132 6580
rect 34076 6526 34078 6578
rect 34078 6526 34130 6578
rect 34130 6526 34132 6578
rect 34076 6524 34132 6526
rect 34188 6130 34244 6132
rect 34188 6078 34190 6130
rect 34190 6078 34242 6130
rect 34242 6078 34244 6130
rect 34188 6076 34244 6078
rect 34412 6300 34468 6356
rect 33068 5628 33124 5684
rect 30604 5180 30660 5236
rect 30044 5122 30100 5124
rect 30044 5070 30046 5122
rect 30046 5070 30098 5122
rect 30098 5070 30100 5122
rect 30044 5068 30100 5070
rect 31052 5068 31108 5124
rect 33628 4898 33684 4900
rect 33628 4846 33630 4898
rect 33630 4846 33682 4898
rect 33682 4846 33684 4898
rect 33628 4844 33684 4846
rect 34972 7474 35028 7476
rect 34972 7422 34974 7474
rect 34974 7422 35026 7474
rect 35026 7422 35028 7474
rect 34972 7420 35028 7422
rect 34860 6300 34916 6356
rect 35308 8204 35364 8260
rect 35868 8258 35924 8260
rect 35868 8206 35870 8258
rect 35870 8206 35922 8258
rect 35922 8206 35924 8258
rect 35868 8204 35924 8206
rect 35644 7756 35700 7812
rect 35756 7868 35812 7924
rect 35868 7698 35924 7700
rect 35868 7646 35870 7698
rect 35870 7646 35922 7698
rect 35922 7646 35924 7698
rect 35868 7644 35924 7646
rect 36876 8652 36932 8708
rect 35308 7196 35364 7252
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 6636 35252 6692
rect 36428 7196 36484 7252
rect 36204 6802 36260 6804
rect 36204 6750 36206 6802
rect 36206 6750 36258 6802
rect 36258 6750 36260 6802
rect 36204 6748 36260 6750
rect 36092 6412 36148 6468
rect 35532 6076 35588 6132
rect 34748 5628 34804 5684
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35980 5122 36036 5124
rect 35980 5070 35982 5122
rect 35982 5070 36034 5122
rect 36034 5070 36036 5122
rect 35980 5068 36036 5070
rect 36988 6690 37044 6692
rect 36988 6638 36990 6690
rect 36990 6638 37042 6690
rect 37042 6638 37044 6690
rect 36988 6636 37044 6638
rect 37100 5740 37156 5796
rect 38444 11452 38500 11508
rect 37772 8988 37828 9044
rect 38332 10556 38388 10612
rect 38220 10332 38276 10388
rect 38108 9826 38164 9828
rect 38108 9774 38110 9826
rect 38110 9774 38162 9826
rect 38162 9774 38164 9826
rect 38108 9772 38164 9774
rect 38668 9938 38724 9940
rect 38668 9886 38670 9938
rect 38670 9886 38722 9938
rect 38722 9886 38724 9938
rect 38668 9884 38724 9886
rect 38444 9436 38500 9492
rect 38556 9042 38612 9044
rect 38556 8990 38558 9042
rect 38558 8990 38610 9042
rect 38610 8990 38612 9042
rect 38556 8988 38612 8990
rect 37996 8876 38052 8932
rect 37436 7756 37492 7812
rect 38668 8204 38724 8260
rect 38892 8316 38948 8372
rect 39004 7756 39060 7812
rect 37772 6636 37828 6692
rect 37436 6300 37492 6356
rect 37996 5794 38052 5796
rect 37996 5742 37998 5794
rect 37998 5742 38050 5794
rect 38050 5742 38052 5794
rect 37996 5740 38052 5742
rect 29484 4226 29540 4228
rect 29484 4174 29486 4226
rect 29486 4174 29538 4226
rect 29538 4174 29540 4226
rect 29484 4172 29540 4174
rect 29932 4226 29988 4228
rect 29932 4174 29934 4226
rect 29934 4174 29986 4226
rect 29986 4174 29988 4226
rect 29932 4172 29988 4174
rect 30492 4226 30548 4228
rect 30492 4174 30494 4226
rect 30494 4174 30546 4226
rect 30546 4174 30548 4226
rect 30492 4172 30548 4174
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35196 3666 35252 3668
rect 35196 3614 35198 3666
rect 35198 3614 35250 3666
rect 35250 3614 35252 3666
rect 35196 3612 35252 3614
rect 37772 3612 37828 3668
rect 38668 5906 38724 5908
rect 38668 5854 38670 5906
rect 38670 5854 38722 5906
rect 38722 5854 38724 5906
rect 38668 5852 38724 5854
rect 38668 5180 38724 5236
rect 39228 11394 39284 11396
rect 39228 11342 39230 11394
rect 39230 11342 39282 11394
rect 39282 11342 39284 11394
rect 39228 11340 39284 11342
rect 39452 8930 39508 8932
rect 39452 8878 39454 8930
rect 39454 8878 39506 8930
rect 39506 8878 39508 8930
rect 39452 8876 39508 8878
rect 40348 17106 40404 17108
rect 40348 17054 40350 17106
rect 40350 17054 40402 17106
rect 40402 17054 40404 17106
rect 40348 17052 40404 17054
rect 40012 16098 40068 16100
rect 40012 16046 40014 16098
rect 40014 16046 40066 16098
rect 40066 16046 40068 16098
rect 40012 16044 40068 16046
rect 42812 20018 42868 20020
rect 42812 19966 42814 20018
rect 42814 19966 42866 20018
rect 42866 19966 42868 20018
rect 42812 19964 42868 19966
rect 42252 19292 42308 19348
rect 41244 18060 41300 18116
rect 42140 18284 42196 18340
rect 39788 15484 39844 15540
rect 40908 15538 40964 15540
rect 40908 15486 40910 15538
rect 40910 15486 40962 15538
rect 40962 15486 40964 15538
rect 40908 15484 40964 15486
rect 40236 15372 40292 15428
rect 41132 15372 41188 15428
rect 39900 15260 39956 15316
rect 40796 15260 40852 15316
rect 39676 15148 39732 15204
rect 42028 16044 42084 16100
rect 44156 22876 44212 22932
rect 43820 20130 43876 20132
rect 43820 20078 43822 20130
rect 43822 20078 43874 20130
rect 43874 20078 43876 20130
rect 43820 20076 43876 20078
rect 43708 19404 43764 19460
rect 44268 19516 44324 19572
rect 44044 19346 44100 19348
rect 44044 19294 44046 19346
rect 44046 19294 44098 19346
rect 44098 19294 44100 19346
rect 44044 19292 44100 19294
rect 43596 16882 43652 16884
rect 43596 16830 43598 16882
rect 43598 16830 43650 16882
rect 43650 16830 43652 16882
rect 43596 16828 43652 16830
rect 43820 16268 43876 16324
rect 43932 18060 43988 18116
rect 44156 16882 44212 16884
rect 44156 16830 44158 16882
rect 44158 16830 44210 16882
rect 44210 16830 44212 16882
rect 44156 16828 44212 16830
rect 43484 15314 43540 15316
rect 43484 15262 43486 15314
rect 43486 15262 43538 15314
rect 43538 15262 43540 15314
rect 43484 15260 43540 15262
rect 41244 14530 41300 14532
rect 41244 14478 41246 14530
rect 41246 14478 41298 14530
rect 41298 14478 41300 14530
rect 41244 14476 41300 14478
rect 41244 14252 41300 14308
rect 39788 13916 39844 13972
rect 40348 13746 40404 13748
rect 40348 13694 40350 13746
rect 40350 13694 40402 13746
rect 40402 13694 40404 13746
rect 40348 13692 40404 13694
rect 41244 13746 41300 13748
rect 41244 13694 41246 13746
rect 41246 13694 41298 13746
rect 41298 13694 41300 13746
rect 41244 13692 41300 13694
rect 39676 13020 39732 13076
rect 41804 13634 41860 13636
rect 41804 13582 41806 13634
rect 41806 13582 41858 13634
rect 41858 13582 41860 13634
rect 41804 13580 41860 13582
rect 42028 14530 42084 14532
rect 42028 14478 42030 14530
rect 42030 14478 42082 14530
rect 42082 14478 42084 14530
rect 42028 14476 42084 14478
rect 42700 14252 42756 14308
rect 42364 13580 42420 13636
rect 43148 13634 43204 13636
rect 43148 13582 43150 13634
rect 43150 13582 43202 13634
rect 43202 13582 43204 13634
rect 43148 13580 43204 13582
rect 41692 12738 41748 12740
rect 41692 12686 41694 12738
rect 41694 12686 41746 12738
rect 41746 12686 41748 12738
rect 41692 12684 41748 12686
rect 41804 12236 41860 12292
rect 39564 6636 39620 6692
rect 39788 10220 39844 10276
rect 40684 9826 40740 9828
rect 40684 9774 40686 9826
rect 40686 9774 40738 9826
rect 40738 9774 40740 9826
rect 40684 9772 40740 9774
rect 41804 10220 41860 10276
rect 42364 9772 42420 9828
rect 43260 12290 43316 12292
rect 43260 12238 43262 12290
rect 43262 12238 43314 12290
rect 43314 12238 43316 12290
rect 43260 12236 43316 12238
rect 44156 12850 44212 12852
rect 44156 12798 44158 12850
rect 44158 12798 44210 12850
rect 44210 12798 44212 12850
rect 44156 12796 44212 12798
rect 43708 12572 43764 12628
rect 44044 10220 44100 10276
rect 41020 9100 41076 9156
rect 42028 9100 42084 9156
rect 40684 8988 40740 9044
rect 41020 8428 41076 8484
rect 42028 8428 42084 8484
rect 39900 7698 39956 7700
rect 39900 7646 39902 7698
rect 39902 7646 39954 7698
rect 39954 7646 39956 7698
rect 39900 7644 39956 7646
rect 41804 8034 41860 8036
rect 41804 7982 41806 8034
rect 41806 7982 41858 8034
rect 41858 7982 41860 8034
rect 41804 7980 41860 7982
rect 40908 7756 40964 7812
rect 40460 7250 40516 7252
rect 40460 7198 40462 7250
rect 40462 7198 40514 7250
rect 40514 7198 40516 7250
rect 40460 7196 40516 7198
rect 42140 8876 42196 8932
rect 42812 8428 42868 8484
rect 42252 8204 42308 8260
rect 41020 7196 41076 7252
rect 40348 6300 40404 6356
rect 41468 6130 41524 6132
rect 41468 6078 41470 6130
rect 41470 6078 41522 6130
rect 41522 6078 41524 6130
rect 41468 6076 41524 6078
rect 42140 6076 42196 6132
rect 40908 5906 40964 5908
rect 40908 5854 40910 5906
rect 40910 5854 40962 5906
rect 40962 5854 40964 5906
rect 40908 5852 40964 5854
rect 41468 5852 41524 5908
rect 43372 9436 43428 9492
rect 44156 9436 44212 9492
rect 43708 9324 43764 9380
rect 44604 27692 44660 27748
rect 44604 26236 44660 26292
rect 43148 8258 43204 8260
rect 43148 8206 43150 8258
rect 43150 8206 43202 8258
rect 43202 8206 43204 8258
rect 43148 8204 43204 8206
rect 43372 8316 43428 8372
rect 43036 7980 43092 8036
rect 43596 7644 43652 7700
rect 43820 6636 43876 6692
rect 43596 6130 43652 6132
rect 43596 6078 43598 6130
rect 43598 6078 43650 6130
rect 43650 6078 43652 6130
rect 43596 6076 43652 6078
rect 42924 6018 42980 6020
rect 42924 5966 42926 6018
rect 42926 5966 42978 6018
rect 42978 5966 42980 6018
rect 42924 5964 42980 5966
rect 43932 5964 43988 6020
rect 44156 6076 44212 6132
rect 41692 5628 41748 5684
rect 39116 4172 39172 4228
rect 41580 5068 41636 5124
rect 42476 4898 42532 4900
rect 42476 4846 42478 4898
rect 42478 4846 42530 4898
rect 42530 4846 42532 4898
rect 42476 4844 42532 4846
rect 41020 4226 41076 4228
rect 41020 4174 41022 4226
rect 41022 4174 41074 4226
rect 41074 4174 41076 4226
rect 41020 4172 41076 4174
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 44156 2716 44212 2772
<< metal3 >>
rect 45200 43092 46000 43120
rect 41906 43036 41916 43092
rect 41972 43036 46000 43092
rect 45200 43008 46000 43036
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 32834 42028 32844 42084
rect 32900 42028 32910 42084
rect 34066 42028 34076 42084
rect 34132 42028 36316 42084
rect 36372 42028 36382 42084
rect 40338 42028 40348 42084
rect 40404 42028 41804 42084
rect 41860 42028 43596 42084
rect 43652 42028 43662 42084
rect 32844 41972 32900 42028
rect 31602 41916 31612 41972
rect 31668 41916 32900 41972
rect 43026 41916 43036 41972
rect 43092 41916 44492 41972
rect 44548 41916 44558 41972
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 32498 41244 32508 41300
rect 32564 41244 33852 41300
rect 33908 41244 33918 41300
rect 29922 41132 29932 41188
rect 29988 41132 31276 41188
rect 31332 41132 31342 41188
rect 39330 41020 39340 41076
rect 39396 41020 42028 41076
rect 42084 41020 42094 41076
rect 35830 40908 35868 40964
rect 35924 40908 35934 40964
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 37538 40684 37548 40740
rect 37604 40684 38108 40740
rect 38164 40684 40908 40740
rect 40964 40684 40974 40740
rect 39106 40572 39116 40628
rect 39172 40572 44044 40628
rect 44100 40572 44110 40628
rect 26898 40460 26908 40516
rect 26964 40460 27244 40516
rect 27300 40460 29260 40516
rect 29316 40460 31612 40516
rect 31668 40460 31678 40516
rect 37874 40460 37884 40516
rect 37940 40460 40236 40516
rect 40292 40460 40796 40516
rect 40852 40460 40862 40516
rect 28578 40348 28588 40404
rect 28644 40348 29708 40404
rect 29764 40348 30268 40404
rect 30324 40348 30334 40404
rect 31266 40348 31276 40404
rect 31332 40348 33068 40404
rect 33124 40348 33134 40404
rect 33506 40348 33516 40404
rect 33572 40348 35084 40404
rect 35140 40348 36428 40404
rect 36484 40348 36494 40404
rect 27682 40236 27692 40292
rect 27748 40236 30156 40292
rect 30212 40236 30222 40292
rect 33730 40236 33740 40292
rect 33796 40236 34412 40292
rect 34468 40236 35644 40292
rect 35700 40236 35710 40292
rect 35858 40236 35868 40292
rect 35924 40236 35980 40292
rect 36036 40236 36046 40292
rect 39778 40236 39788 40292
rect 39844 40236 43820 40292
rect 43876 40236 43886 40292
rect 33954 40124 33964 40180
rect 34020 40124 34524 40180
rect 34580 40124 35196 40180
rect 35252 40124 35262 40180
rect 40226 40124 40236 40180
rect 40292 40124 41356 40180
rect 41412 40124 41422 40180
rect 41906 40124 41916 40180
rect 41972 40124 44156 40180
rect 44212 40124 44222 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 34066 39788 34076 39844
rect 34132 39788 35308 39844
rect 35364 39788 35374 39844
rect 45200 39732 46000 39760
rect 26786 39676 26796 39732
rect 26852 39676 29932 39732
rect 29988 39676 29998 39732
rect 30370 39676 30380 39732
rect 30436 39676 32060 39732
rect 32116 39676 32126 39732
rect 38994 39676 39004 39732
rect 39060 39676 40572 39732
rect 40628 39676 40638 39732
rect 43138 39676 43148 39732
rect 43204 39676 46000 39732
rect 45200 39648 46000 39676
rect 26674 39564 26684 39620
rect 26740 39564 28364 39620
rect 28420 39564 30044 39620
rect 30100 39564 30110 39620
rect 31826 39564 31836 39620
rect 31892 39564 32508 39620
rect 32564 39564 32574 39620
rect 34850 39564 34860 39620
rect 34916 39564 36988 39620
rect 37044 39564 37054 39620
rect 41234 39564 41244 39620
rect 41300 39564 43932 39620
rect 43988 39564 43998 39620
rect 28018 39340 28028 39396
rect 28084 39340 29036 39396
rect 29092 39340 29102 39396
rect 30146 39228 30156 39284
rect 30212 39228 31276 39284
rect 31332 39228 31342 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 39890 39116 39900 39172
rect 39956 39116 41020 39172
rect 41076 39116 41086 39172
rect 29810 39004 29820 39060
rect 29876 39004 30380 39060
rect 30436 39004 30446 39060
rect 36278 39004 36316 39060
rect 36372 39004 36382 39060
rect 38882 39004 38892 39060
rect 38948 39004 39788 39060
rect 39844 39004 40460 39060
rect 40516 39004 40526 39060
rect 29698 38892 29708 38948
rect 29764 38892 30492 38948
rect 30548 38892 30558 38948
rect 38434 38892 38444 38948
rect 38500 38892 39676 38948
rect 39732 38892 39742 38948
rect 40786 38892 40796 38948
rect 40852 38892 41916 38948
rect 41972 38892 41982 38948
rect 29474 38780 29484 38836
rect 29540 38780 30044 38836
rect 30100 38780 30604 38836
rect 30660 38780 30670 38836
rect 32610 38780 32620 38836
rect 32676 38780 33068 38836
rect 33124 38780 33134 38836
rect 37426 38780 37436 38836
rect 37492 38780 39228 38836
rect 39284 38780 39294 38836
rect 29026 38668 29036 38724
rect 29092 38668 29820 38724
rect 29876 38668 29886 38724
rect 31602 38668 31612 38724
rect 31668 38668 32284 38724
rect 32340 38668 32350 38724
rect 34514 38668 34524 38724
rect 34580 38668 35980 38724
rect 36036 38668 36046 38724
rect 37314 38668 37324 38724
rect 37380 38668 38780 38724
rect 38836 38668 40068 38724
rect 40012 38612 40068 38668
rect 27010 38556 27020 38612
rect 27076 38556 30268 38612
rect 30324 38556 30334 38612
rect 37538 38556 37548 38612
rect 37604 38556 38108 38612
rect 38164 38556 39116 38612
rect 39172 38556 39182 38612
rect 40002 38556 40012 38612
rect 40068 38556 40078 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 27906 38108 27916 38164
rect 27972 38108 29260 38164
rect 29316 38108 29326 38164
rect 30818 38108 30828 38164
rect 30884 38108 36988 38164
rect 37044 38108 38220 38164
rect 38276 38108 38286 38164
rect 33282 37996 33292 38052
rect 33348 37996 34076 38052
rect 34132 37996 34748 38052
rect 34804 37996 35420 38052
rect 35476 37996 35486 38052
rect 40114 37996 40124 38052
rect 40180 37996 40908 38052
rect 40964 37996 40974 38052
rect 41794 37996 41804 38052
rect 41860 37996 42700 38052
rect 42756 37996 43596 38052
rect 43652 37996 43662 38052
rect 40450 37884 40460 37940
rect 40516 37884 43036 37940
rect 43092 37884 43102 37940
rect 40226 37772 40236 37828
rect 40292 37772 40684 37828
rect 40740 37772 42588 37828
rect 42644 37772 42654 37828
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 33058 37212 33068 37268
rect 33124 37212 33964 37268
rect 34020 37212 35084 37268
rect 35140 37212 35150 37268
rect 35858 37212 35868 37268
rect 35924 37212 36764 37268
rect 36820 37212 36830 37268
rect 38210 37212 38220 37268
rect 38276 37212 39452 37268
rect 39508 37212 39518 37268
rect 39666 37212 39676 37268
rect 39732 37212 40796 37268
rect 40852 37212 41580 37268
rect 41636 37212 41646 37268
rect 35084 37156 35140 37212
rect 35084 37100 37660 37156
rect 37716 37100 37726 37156
rect 43474 36988 43484 37044
rect 43540 36988 43708 37044
rect 43652 36932 43708 36988
rect 43652 36876 45332 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 45276 36596 45332 36876
rect 45052 36540 45332 36596
rect 26450 36428 26460 36484
rect 26516 36428 27132 36484
rect 27188 36428 27198 36484
rect 45052 36372 45108 36540
rect 45200 36372 46000 36400
rect 9426 36316 9436 36372
rect 9492 36316 10444 36372
rect 10500 36316 10510 36372
rect 26226 36316 26236 36372
rect 26292 36316 27468 36372
rect 27524 36316 27534 36372
rect 31042 36316 31052 36372
rect 31108 36316 32732 36372
rect 32788 36316 32798 36372
rect 45052 36316 46000 36372
rect 45200 36288 46000 36316
rect 26002 36204 26012 36260
rect 26068 36204 27916 36260
rect 27972 36204 27982 36260
rect 43922 36204 43932 36260
rect 43988 36204 44492 36260
rect 44548 36204 44558 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 24210 35980 24220 36036
rect 24276 35980 26124 36036
rect 26180 35980 27356 36036
rect 27412 35980 27422 36036
rect 17938 35868 17948 35924
rect 18004 35868 19404 35924
rect 19460 35868 19470 35924
rect 24658 35868 24668 35924
rect 24724 35868 26908 35924
rect 26964 35868 26974 35924
rect 35970 35868 35980 35924
rect 36036 35868 37212 35924
rect 37268 35868 37660 35924
rect 37716 35868 37726 35924
rect 16146 35756 16156 35812
rect 16212 35756 16716 35812
rect 16772 35756 18620 35812
rect 18676 35756 18686 35812
rect 23538 35756 23548 35812
rect 23604 35756 26460 35812
rect 26516 35756 26526 35812
rect 30370 35756 30380 35812
rect 30436 35756 32956 35812
rect 33012 35756 33022 35812
rect 34850 35756 34860 35812
rect 34916 35756 35532 35812
rect 35588 35756 36764 35812
rect 36820 35756 36830 35812
rect 10770 35644 10780 35700
rect 10836 35644 20188 35700
rect 23762 35644 23772 35700
rect 23828 35644 24444 35700
rect 24500 35644 25452 35700
rect 25508 35644 26348 35700
rect 26404 35644 26414 35700
rect 36306 35644 36316 35700
rect 36372 35644 37436 35700
rect 37492 35644 37502 35700
rect 38994 35644 39004 35700
rect 39060 35644 41132 35700
rect 41188 35644 41198 35700
rect 43652 35644 43820 35700
rect 43876 35644 43886 35700
rect 20132 35476 20188 35644
rect 24322 35532 24332 35588
rect 24388 35532 28700 35588
rect 28756 35532 28766 35588
rect 32498 35532 32508 35588
rect 32564 35532 35420 35588
rect 35476 35532 35486 35588
rect 41346 35532 41356 35588
rect 41412 35532 43148 35588
rect 43204 35532 43214 35588
rect 20132 35420 21084 35476
rect 21140 35420 21150 35476
rect 23090 35420 23100 35476
rect 23156 35420 25228 35476
rect 25284 35420 26236 35476
rect 26292 35420 26302 35476
rect 31892 35420 33348 35476
rect 31826 35308 31836 35364
rect 31892 35308 31948 35420
rect 33292 35364 33348 35420
rect 43652 35364 43708 35644
rect 33282 35308 33292 35364
rect 33348 35308 33358 35364
rect 40338 35308 40348 35364
rect 40404 35308 41244 35364
rect 41300 35308 43708 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 15810 35196 15820 35252
rect 15876 35196 17500 35252
rect 17556 35196 18284 35252
rect 18340 35196 18350 35252
rect 24434 35196 24444 35252
rect 24500 35196 24892 35252
rect 24948 35196 27804 35252
rect 27860 35196 27870 35252
rect 40002 35084 40012 35140
rect 40068 35084 40078 35140
rect 7298 34972 7308 35028
rect 7364 34972 9324 35028
rect 9380 34972 9390 35028
rect 26114 34972 26124 35028
rect 26180 34972 29708 35028
rect 29764 34972 29774 35028
rect 32274 34972 32284 35028
rect 32340 34972 33180 35028
rect 33236 34972 33246 35028
rect 33618 34972 33628 35028
rect 33684 34972 35420 35028
rect 35476 34972 35486 35028
rect 35634 34972 35644 35028
rect 35700 34972 36988 35028
rect 37044 34972 37054 35028
rect 14578 34860 14588 34916
rect 14644 34860 16828 34916
rect 16884 34860 16894 34916
rect 27682 34860 27692 34916
rect 27748 34860 29372 34916
rect 29428 34860 29438 34916
rect 35298 34860 35308 34916
rect 35364 34860 35980 34916
rect 36036 34860 36428 34916
rect 36484 34860 36494 34916
rect 15922 34748 15932 34804
rect 15988 34748 17388 34804
rect 17444 34748 17454 34804
rect 18274 34748 18284 34804
rect 18340 34748 18732 34804
rect 18788 34748 20412 34804
rect 20468 34748 20478 34804
rect 24546 34748 24556 34804
rect 24612 34748 26460 34804
rect 26516 34748 26526 34804
rect 28130 34748 28140 34804
rect 28196 34748 28700 34804
rect 28756 34748 29932 34804
rect 29988 34748 29998 34804
rect 31154 34748 31164 34804
rect 31220 34748 37100 34804
rect 37156 34748 37166 34804
rect 40012 34692 40068 35084
rect 40450 34860 40460 34916
rect 40516 34860 41804 34916
rect 41860 34860 41870 34916
rect 17938 34636 17948 34692
rect 18004 34636 19964 34692
rect 20020 34636 20972 34692
rect 21028 34636 21038 34692
rect 26226 34636 26236 34692
rect 26292 34636 27244 34692
rect 27300 34636 28364 34692
rect 28420 34636 28430 34692
rect 34402 34636 34412 34692
rect 34468 34636 36204 34692
rect 36260 34636 37772 34692
rect 37828 34636 37838 34692
rect 40002 34636 40012 34692
rect 40068 34636 40078 34692
rect 36082 34524 36092 34580
rect 36148 34524 38108 34580
rect 38164 34524 38174 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 36194 34412 36204 34468
rect 36260 34412 37324 34468
rect 37380 34412 38668 34468
rect 38724 34412 39228 34468
rect 39284 34412 39294 34468
rect 11442 34300 11452 34356
rect 11508 34300 18844 34356
rect 18900 34300 18910 34356
rect 21074 34300 21084 34356
rect 21140 34300 22092 34356
rect 22148 34300 22158 34356
rect 26450 34300 26460 34356
rect 26516 34300 28588 34356
rect 28644 34300 29148 34356
rect 29204 34300 29214 34356
rect 32386 34300 32396 34356
rect 32452 34300 39452 34356
rect 39508 34300 41804 34356
rect 41860 34300 41870 34356
rect 24098 34188 24108 34244
rect 24164 34188 25788 34244
rect 25844 34188 25854 34244
rect 27458 34188 27468 34244
rect 27524 34188 31052 34244
rect 31108 34188 31118 34244
rect 32274 34188 32284 34244
rect 32340 34188 33516 34244
rect 33572 34188 39340 34244
rect 39396 34188 39406 34244
rect 39890 34188 39900 34244
rect 39956 34188 40908 34244
rect 40964 34188 40974 34244
rect 41234 34188 41244 34244
rect 41300 34188 42588 34244
rect 42644 34188 42654 34244
rect 41244 34132 41300 34188
rect 12674 34076 12684 34132
rect 12740 34076 13468 34132
rect 13524 34076 16492 34132
rect 16548 34076 17276 34132
rect 17332 34076 17342 34132
rect 17714 34076 17724 34132
rect 17780 34076 18620 34132
rect 18676 34076 21980 34132
rect 22036 34076 22046 34132
rect 24770 34076 24780 34132
rect 24836 34076 28252 34132
rect 28308 34076 28318 34132
rect 28914 34076 28924 34132
rect 28980 34076 31948 34132
rect 32004 34076 32014 34132
rect 34076 34076 36540 34132
rect 36596 34076 36606 34132
rect 38658 34076 38668 34132
rect 38724 34076 40348 34132
rect 40404 34076 41300 34132
rect 42130 34076 42140 34132
rect 42196 34076 43708 34132
rect 17276 34020 17332 34076
rect 17276 33964 18172 34020
rect 18228 33964 18238 34020
rect 25554 33964 25564 34020
rect 25620 33964 26796 34020
rect 26852 33964 26862 34020
rect 32050 33964 32060 34020
rect 32116 33964 33852 34020
rect 33908 33964 33918 34020
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 34076 33684 34132 34076
rect 43652 34020 43708 34076
rect 36194 33964 36204 34020
rect 36260 33964 36652 34020
rect 36708 33964 36718 34020
rect 43652 33964 43820 34020
rect 43876 33964 44492 34020
rect 44548 33964 44558 34020
rect 34514 33852 34524 33908
rect 34580 33852 37324 33908
rect 37380 33852 38332 33908
rect 38388 33852 38398 33908
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 28018 33628 28028 33684
rect 28084 33628 30604 33684
rect 30660 33628 30670 33684
rect 32498 33628 32508 33684
rect 32564 33628 34132 33684
rect 36306 33628 36316 33684
rect 36372 33628 37660 33684
rect 37716 33628 37726 33684
rect 25330 33516 25340 33572
rect 25396 33516 25788 33572
rect 25844 33516 25854 33572
rect 35410 33516 35420 33572
rect 35476 33516 35756 33572
rect 35812 33516 36428 33572
rect 36484 33516 36494 33572
rect 6962 33404 6972 33460
rect 7028 33404 7756 33460
rect 7812 33404 8876 33460
rect 8932 33404 8942 33460
rect 35858 33404 35868 33460
rect 35924 33404 37660 33460
rect 37716 33404 37726 33460
rect 17378 33292 17388 33348
rect 17444 33292 17948 33348
rect 18004 33292 18620 33348
rect 18676 33292 20524 33348
rect 20580 33292 20590 33348
rect 24210 33292 24220 33348
rect 24276 33292 25788 33348
rect 25844 33292 25854 33348
rect 35522 33292 35532 33348
rect 35588 33292 38108 33348
rect 38164 33292 38174 33348
rect 7298 33180 7308 33236
rect 7364 33180 10108 33236
rect 10164 33180 10892 33236
rect 10948 33180 10958 33236
rect 22194 33180 22204 33236
rect 22260 33180 25900 33236
rect 25956 33180 26236 33236
rect 26292 33180 26302 33236
rect 30146 33180 30156 33236
rect 30212 33180 35644 33236
rect 35700 33180 35710 33236
rect 37426 33180 37436 33236
rect 37492 33180 38780 33236
rect 38836 33180 39676 33236
rect 39732 33180 40572 33236
rect 40628 33180 40638 33236
rect 24994 33068 25004 33124
rect 25060 33068 25676 33124
rect 25732 33068 27132 33124
rect 27188 33068 27198 33124
rect 33842 33068 33852 33124
rect 33908 33068 36204 33124
rect 36260 33068 36270 33124
rect 43138 33068 43148 33124
rect 43204 33068 43708 33124
rect 43652 33012 43708 33068
rect 45200 33012 46000 33040
rect 24658 32956 24668 33012
rect 24724 32956 26908 33012
rect 26964 32956 26974 33012
rect 43652 32956 46000 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 45200 32928 46000 32956
rect 24658 32732 24668 32788
rect 24724 32732 25564 32788
rect 25620 32732 26796 32788
rect 26852 32732 26862 32788
rect 40114 32732 40124 32788
rect 40180 32732 40348 32788
rect 40404 32732 40414 32788
rect 41346 32732 41356 32788
rect 41412 32732 42924 32788
rect 42980 32732 42990 32788
rect 40348 32676 40404 32732
rect 7970 32620 7980 32676
rect 8036 32620 9548 32676
rect 9604 32620 9614 32676
rect 14914 32620 14924 32676
rect 14980 32620 15596 32676
rect 15652 32620 16156 32676
rect 16212 32620 17500 32676
rect 17556 32620 17566 32676
rect 24322 32620 24332 32676
rect 24388 32620 26684 32676
rect 26740 32620 26750 32676
rect 28690 32620 28700 32676
rect 28756 32620 29036 32676
rect 29092 32620 29102 32676
rect 35970 32620 35980 32676
rect 36036 32620 36764 32676
rect 36820 32620 36830 32676
rect 39442 32620 39452 32676
rect 39508 32620 40012 32676
rect 40068 32620 40078 32676
rect 40348 32620 43596 32676
rect 43652 32620 43662 32676
rect 13122 32508 13132 32564
rect 13188 32508 14588 32564
rect 14644 32508 14654 32564
rect 22978 32508 22988 32564
rect 23044 32508 25340 32564
rect 25396 32508 27020 32564
rect 27076 32508 27086 32564
rect 35186 32508 35196 32564
rect 35252 32508 37884 32564
rect 37940 32508 38892 32564
rect 38948 32508 38958 32564
rect 41010 32508 41020 32564
rect 41076 32508 42476 32564
rect 42532 32508 42542 32564
rect 20132 32396 20860 32452
rect 20916 32396 20926 32452
rect 26002 32396 26012 32452
rect 26068 32396 27916 32452
rect 27972 32396 27982 32452
rect 34962 32396 34972 32452
rect 35028 32396 36316 32452
rect 36372 32396 36382 32452
rect 20132 32340 20188 32396
rect 11554 32284 11564 32340
rect 11620 32284 17164 32340
rect 17220 32284 20188 32340
rect 40226 32284 40236 32340
rect 40292 32284 41132 32340
rect 41188 32284 41198 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 40348 32060 40460 32116
rect 40516 32060 40526 32116
rect 31826 31948 31836 32004
rect 31892 31948 33180 32004
rect 33236 31948 33246 32004
rect 37090 31948 37100 32004
rect 37156 31948 39564 32004
rect 39620 31948 39630 32004
rect 40348 31892 40404 32060
rect 6066 31836 6076 31892
rect 6132 31836 7980 31892
rect 8036 31836 8046 31892
rect 15026 31836 15036 31892
rect 15092 31836 16268 31892
rect 16324 31836 16334 31892
rect 29698 31836 29708 31892
rect 29764 31836 31052 31892
rect 31108 31836 31118 31892
rect 35298 31836 35308 31892
rect 35364 31836 37212 31892
rect 37268 31836 37278 31892
rect 37986 31836 37996 31892
rect 38052 31836 38668 31892
rect 38724 31836 40404 31892
rect 39554 31724 39564 31780
rect 39620 31724 40348 31780
rect 40404 31724 40414 31780
rect 25890 31612 25900 31668
rect 25956 31612 27244 31668
rect 27300 31612 27804 31668
rect 27860 31612 27870 31668
rect 17826 31500 17836 31556
rect 17892 31500 18284 31556
rect 18340 31500 26068 31556
rect 26226 31500 26236 31556
rect 26292 31500 27132 31556
rect 27188 31500 27198 31556
rect 38434 31500 38444 31556
rect 38500 31500 41020 31556
rect 41076 31500 41086 31556
rect 26012 31444 26068 31500
rect 26012 31388 27020 31444
rect 27076 31388 27916 31444
rect 27972 31388 31612 31444
rect 31668 31388 31678 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 39666 31276 39676 31332
rect 39732 31276 40124 31332
rect 40180 31276 40190 31332
rect 26002 31052 26012 31108
rect 26068 31052 33068 31108
rect 33124 31052 33134 31108
rect 39330 31052 39340 31108
rect 39396 31052 39900 31108
rect 39956 31052 40572 31108
rect 40628 31052 40638 31108
rect 16706 30940 16716 30996
rect 16772 30940 18396 30996
rect 18452 30940 18462 30996
rect 19842 30940 19852 30996
rect 19908 30940 20748 30996
rect 20804 30940 20814 30996
rect 29922 30940 29932 30996
rect 29988 30940 32620 30996
rect 32676 30940 33292 30996
rect 33348 30940 33358 30996
rect 39218 30940 39228 30996
rect 39284 30940 40404 30996
rect 41010 30940 41020 30996
rect 41076 30940 43708 30996
rect 43764 30940 43774 30996
rect 40348 30884 40404 30940
rect 21410 30828 21420 30884
rect 21476 30828 22204 30884
rect 22260 30828 22764 30884
rect 22820 30828 22830 30884
rect 31602 30828 31612 30884
rect 31668 30828 34076 30884
rect 34132 30828 34142 30884
rect 36978 30828 36988 30884
rect 37044 30828 38668 30884
rect 38724 30828 39788 30884
rect 39844 30828 39854 30884
rect 40348 30828 40908 30884
rect 40964 30828 41804 30884
rect 41860 30828 41870 30884
rect 18610 30716 18620 30772
rect 18676 30716 20412 30772
rect 20468 30716 20478 30772
rect 31490 30716 31500 30772
rect 31556 30716 35308 30772
rect 35364 30716 35374 30772
rect 36866 30604 36876 30660
rect 36932 30604 37436 30660
rect 37492 30604 37502 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 31266 30380 31276 30436
rect 31332 30380 33740 30436
rect 33796 30380 33806 30436
rect 43138 30380 43148 30436
rect 43204 30380 43708 30436
rect 15138 30268 15148 30324
rect 15204 30268 15932 30324
rect 15988 30268 17052 30324
rect 17108 30268 17118 30324
rect 30706 30268 30716 30324
rect 30772 30268 33404 30324
rect 33460 30268 33470 30324
rect 33618 30268 33628 30324
rect 33684 30268 35084 30324
rect 35140 30268 35150 30324
rect 39442 30268 39452 30324
rect 39508 30268 41916 30324
rect 41972 30268 41982 30324
rect 43652 30212 43708 30380
rect 17826 30156 17836 30212
rect 17892 30156 20972 30212
rect 21028 30156 21038 30212
rect 29586 30156 29596 30212
rect 29652 30156 30268 30212
rect 30324 30156 30334 30212
rect 41234 30156 41244 30212
rect 41300 30156 42588 30212
rect 42644 30156 42654 30212
rect 43652 30156 45332 30212
rect 21634 30044 21644 30100
rect 21700 30044 27468 30100
rect 27524 30044 29708 30100
rect 29764 30044 30604 30100
rect 30660 30044 30670 30100
rect 36530 30044 36540 30100
rect 36596 30044 37100 30100
rect 37156 30044 37166 30100
rect 39106 30044 39116 30100
rect 39172 30044 42028 30100
rect 42084 30044 43484 30100
rect 43540 30044 43550 30100
rect 26450 29932 26460 29988
rect 26516 29932 27804 29988
rect 27860 29932 27870 29988
rect 30604 29876 30660 30044
rect 31714 29932 31724 29988
rect 31780 29932 33628 29988
rect 33684 29932 33694 29988
rect 37986 29932 37996 29988
rect 38052 29932 38780 29988
rect 38836 29932 38846 29988
rect 45276 29876 45332 30156
rect 30604 29820 31948 29876
rect 32004 29820 32014 29876
rect 45052 29820 45332 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 24770 29708 24780 29764
rect 24836 29708 25228 29764
rect 25284 29708 25676 29764
rect 25732 29708 25742 29764
rect 26226 29708 26236 29764
rect 26292 29708 27132 29764
rect 27188 29708 27580 29764
rect 27636 29708 27646 29764
rect 29026 29708 29036 29764
rect 29092 29708 29708 29764
rect 29764 29708 32732 29764
rect 32788 29708 32798 29764
rect 45052 29652 45108 29820
rect 45200 29652 46000 29680
rect 11442 29596 11452 29652
rect 11508 29596 13244 29652
rect 13300 29596 13310 29652
rect 24546 29596 24556 29652
rect 24612 29596 25340 29652
rect 25396 29596 25406 29652
rect 26338 29596 26348 29652
rect 26404 29596 28588 29652
rect 28644 29596 28654 29652
rect 32498 29596 32508 29652
rect 32564 29596 34188 29652
rect 34244 29596 34254 29652
rect 45052 29596 46000 29652
rect 45200 29568 46000 29596
rect 16258 29484 16268 29540
rect 16324 29484 17500 29540
rect 17556 29484 18284 29540
rect 18340 29484 18350 29540
rect 26674 29484 26684 29540
rect 26740 29484 28028 29540
rect 28084 29484 28700 29540
rect 28756 29484 28766 29540
rect 31266 29484 31276 29540
rect 31332 29484 33068 29540
rect 33124 29484 33134 29540
rect 8866 29372 8876 29428
rect 8932 29372 9548 29428
rect 9604 29372 10780 29428
rect 10836 29372 10846 29428
rect 17826 29372 17836 29428
rect 17892 29372 18396 29428
rect 18452 29372 21308 29428
rect 21364 29372 21374 29428
rect 24658 29372 24668 29428
rect 24724 29372 27020 29428
rect 27076 29372 27086 29428
rect 27906 29372 27916 29428
rect 27972 29372 29260 29428
rect 29316 29372 29326 29428
rect 30146 29372 30156 29428
rect 30212 29372 30828 29428
rect 30884 29372 30894 29428
rect 34738 29372 34748 29428
rect 34804 29372 35756 29428
rect 35812 29372 40012 29428
rect 40068 29372 40908 29428
rect 40964 29372 42140 29428
rect 42196 29372 42206 29428
rect 13010 29260 13020 29316
rect 13076 29260 13916 29316
rect 13972 29260 13982 29316
rect 16818 29260 16828 29316
rect 16884 29260 19180 29316
rect 19236 29260 19246 29316
rect 34290 29260 34300 29316
rect 34356 29260 37996 29316
rect 38052 29260 38062 29316
rect 32386 29148 32396 29204
rect 32452 29148 34748 29204
rect 34804 29148 34814 29204
rect 29810 29036 29820 29092
rect 29876 29036 30716 29092
rect 30772 29036 30782 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 30258 28812 30268 28868
rect 30324 28812 30334 28868
rect 30706 28812 30716 28868
rect 30772 28812 31724 28868
rect 31780 28812 31790 28868
rect 6066 28700 6076 28756
rect 6132 28700 8316 28756
rect 8372 28700 8382 28756
rect 28802 28700 28812 28756
rect 28868 28700 29596 28756
rect 29652 28700 29662 28756
rect 30268 28644 30324 28812
rect 7634 28588 7644 28644
rect 7700 28588 8876 28644
rect 8932 28588 8942 28644
rect 20626 28588 20636 28644
rect 20692 28588 21308 28644
rect 21364 28588 21374 28644
rect 25106 28588 25116 28644
rect 25172 28588 25564 28644
rect 25620 28588 25630 28644
rect 26898 28588 26908 28644
rect 26964 28588 28700 28644
rect 28756 28588 29708 28644
rect 29764 28588 30324 28644
rect 31938 28588 31948 28644
rect 32004 28588 33740 28644
rect 33796 28588 34300 28644
rect 34356 28588 34366 28644
rect 14018 28476 14028 28532
rect 14084 28476 16044 28532
rect 16100 28476 16110 28532
rect 27794 28476 27804 28532
rect 27860 28476 29820 28532
rect 29876 28476 29886 28532
rect 30258 28364 30268 28420
rect 30324 28364 32508 28420
rect 32564 28364 32574 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 26002 28028 26012 28084
rect 26068 28028 28252 28084
rect 28308 28028 28318 28084
rect 11106 27916 11116 27972
rect 11172 27916 12236 27972
rect 12292 27916 12302 27972
rect 13794 27916 13804 27972
rect 13860 27916 17388 27972
rect 17444 27916 17454 27972
rect 25890 27916 25900 27972
rect 25956 27916 27244 27972
rect 27300 27916 28364 27972
rect 28420 27916 28430 27972
rect 29138 27916 29148 27972
rect 29204 27916 30268 27972
rect 30324 27916 30334 27972
rect 19170 27804 19180 27860
rect 19236 27804 20188 27860
rect 20244 27804 20254 27860
rect 24434 27804 24444 27860
rect 24500 27804 26572 27860
rect 26628 27804 26638 27860
rect 29138 27804 29148 27860
rect 29204 27804 29596 27860
rect 29652 27804 29662 27860
rect 11554 27692 11564 27748
rect 11620 27692 12460 27748
rect 12516 27692 12526 27748
rect 20290 27692 20300 27748
rect 20356 27692 20860 27748
rect 20916 27692 21980 27748
rect 22036 27692 22046 27748
rect 23986 27692 23996 27748
rect 24052 27692 27468 27748
rect 27524 27692 27534 27748
rect 29250 27692 29260 27748
rect 29316 27692 30380 27748
rect 30436 27692 30446 27748
rect 41794 27692 41804 27748
rect 41860 27692 43148 27748
rect 43204 27692 43214 27748
rect 43586 27692 43596 27748
rect 43652 27692 44156 27748
rect 44212 27692 44604 27748
rect 44660 27692 44670 27748
rect 10770 27580 10780 27636
rect 10836 27580 11900 27636
rect 11956 27580 11966 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 8530 27244 8540 27300
rect 8596 27244 9212 27300
rect 9268 27244 20188 27300
rect 26226 27244 26236 27300
rect 26292 27244 27804 27300
rect 27860 27244 27870 27300
rect 20132 27188 20188 27244
rect 8978 27132 8988 27188
rect 9044 27132 10108 27188
rect 10164 27132 11228 27188
rect 11284 27132 11294 27188
rect 20132 27132 35084 27188
rect 35140 27132 37100 27188
rect 37156 27132 37166 27188
rect 8754 27020 8764 27076
rect 8820 27020 9660 27076
rect 9716 27020 11004 27076
rect 11060 27020 11070 27076
rect 26562 27020 26572 27076
rect 26628 27020 27356 27076
rect 27412 27020 27422 27076
rect 10210 26908 10220 26964
rect 10276 26908 12236 26964
rect 12292 26908 12302 26964
rect 15698 26908 15708 26964
rect 15764 26908 16716 26964
rect 16772 26908 16782 26964
rect 18274 26908 18284 26964
rect 18340 26908 18956 26964
rect 19012 26908 19022 26964
rect 26002 26908 26012 26964
rect 26068 26908 27020 26964
rect 27076 26908 27086 26964
rect 34738 26908 34748 26964
rect 34804 26908 35644 26964
rect 35700 26908 36204 26964
rect 36260 26908 36270 26964
rect 43138 26908 43148 26964
rect 43204 26908 44268 26964
rect 44324 26908 44334 26964
rect 20402 26796 20412 26852
rect 20468 26796 21308 26852
rect 21364 26796 21374 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 12338 26572 12348 26628
rect 12404 26572 13468 26628
rect 13524 26572 13534 26628
rect 13122 26460 13132 26516
rect 13188 26460 13916 26516
rect 13972 26460 13982 26516
rect 10546 26348 10556 26404
rect 10612 26348 14140 26404
rect 14196 26348 14206 26404
rect 22530 26348 22540 26404
rect 22596 26348 23548 26404
rect 23604 26348 23614 26404
rect 30034 26348 30044 26404
rect 30100 26348 30828 26404
rect 30884 26348 30894 26404
rect 37986 26348 37996 26404
rect 38052 26348 38892 26404
rect 38948 26348 38958 26404
rect 45200 26292 46000 26320
rect 16818 26236 16828 26292
rect 16884 26236 18732 26292
rect 18788 26236 19628 26292
rect 19684 26236 19694 26292
rect 21298 26236 21308 26292
rect 21364 26236 23996 26292
rect 24052 26236 24062 26292
rect 44594 26236 44604 26292
rect 44660 26236 46000 26292
rect 45200 26208 46000 26236
rect 19842 26124 19852 26180
rect 19908 26124 20412 26180
rect 20468 26124 20478 26180
rect 34066 26124 34076 26180
rect 34132 26124 35084 26180
rect 35140 26124 37884 26180
rect 37940 26124 37950 26180
rect 9762 26012 9772 26068
rect 9828 26012 12348 26068
rect 12404 26012 12414 26068
rect 16706 26012 16716 26068
rect 16772 26012 17388 26068
rect 17444 26012 17454 26068
rect 31826 26012 31836 26068
rect 31892 26012 43820 26068
rect 43876 26012 43886 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 16258 25676 16268 25732
rect 16324 25676 17500 25732
rect 17556 25676 19740 25732
rect 19796 25676 19806 25732
rect 23986 25676 23996 25732
rect 24052 25676 25116 25732
rect 25172 25676 25182 25732
rect 21410 25564 21420 25620
rect 21476 25564 22428 25620
rect 22484 25564 22494 25620
rect 34626 25564 34636 25620
rect 34692 25564 41468 25620
rect 41524 25564 44044 25620
rect 44100 25564 44110 25620
rect 25666 25452 25676 25508
rect 25732 25452 26348 25508
rect 26404 25452 31948 25508
rect 32004 25452 32014 25508
rect 18610 25340 18620 25396
rect 18676 25340 19292 25396
rect 19348 25340 19964 25396
rect 20020 25340 20030 25396
rect 6962 25228 6972 25284
rect 7028 25228 7756 25284
rect 7812 25228 7822 25284
rect 10322 25228 10332 25284
rect 10388 25228 11676 25284
rect 11732 25228 12796 25284
rect 12852 25228 12862 25284
rect 16034 25228 16044 25284
rect 16100 25228 19628 25284
rect 19684 25228 19694 25284
rect 28578 25228 28588 25284
rect 28644 25228 29260 25284
rect 29316 25228 31724 25284
rect 31780 25228 31790 25284
rect 37874 25228 37884 25284
rect 37940 25228 38444 25284
rect 38500 25228 38510 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 9874 24892 9884 24948
rect 9940 24892 10892 24948
rect 10948 24892 10958 24948
rect 20290 24892 20300 24948
rect 20356 24892 21980 24948
rect 22036 24892 22046 24948
rect 35858 24892 35868 24948
rect 35924 24892 37212 24948
rect 37268 24892 37278 24948
rect 17938 24780 17948 24836
rect 18004 24780 19068 24836
rect 19124 24780 19134 24836
rect 22530 24780 22540 24836
rect 22596 24780 23660 24836
rect 23716 24780 24108 24836
rect 24164 24780 24174 24836
rect 27234 24780 27244 24836
rect 27300 24780 27804 24836
rect 27860 24780 27870 24836
rect 18050 24668 18060 24724
rect 18116 24668 18844 24724
rect 18900 24668 18910 24724
rect 33058 24668 33068 24724
rect 33124 24668 34972 24724
rect 35028 24668 36092 24724
rect 36148 24668 38332 24724
rect 38388 24668 38398 24724
rect 39442 24668 39452 24724
rect 39508 24668 41468 24724
rect 41524 24668 41534 24724
rect 26450 24556 26460 24612
rect 26516 24556 27020 24612
rect 27076 24556 33740 24612
rect 33796 24556 33806 24612
rect 15810 24444 15820 24500
rect 15876 24444 18284 24500
rect 18340 24444 18350 24500
rect 19170 24444 19180 24500
rect 19236 24444 19628 24500
rect 19684 24444 22428 24500
rect 22484 24444 23772 24500
rect 23828 24444 23838 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 26898 24220 26908 24276
rect 26964 24220 27244 24276
rect 27300 24220 27310 24276
rect 7186 24108 7196 24164
rect 7252 24108 8428 24164
rect 18498 24108 18508 24164
rect 18564 24108 19740 24164
rect 19796 24108 19806 24164
rect 8372 23940 8428 24108
rect 8372 23884 8540 23940
rect 8596 23884 8606 23940
rect 29474 23884 29484 23940
rect 29540 23884 32284 23940
rect 32340 23884 35196 23940
rect 35252 23884 35262 23940
rect 7858 23772 7868 23828
rect 7924 23772 9548 23828
rect 9604 23772 9614 23828
rect 19058 23660 19068 23716
rect 19124 23660 19852 23716
rect 19908 23660 20300 23716
rect 20356 23660 25452 23716
rect 25508 23660 28140 23716
rect 28196 23660 28924 23716
rect 28980 23660 28990 23716
rect 35522 23660 35532 23716
rect 35588 23660 35644 23716
rect 35700 23660 35710 23716
rect 27794 23548 27804 23604
rect 27860 23548 29260 23604
rect 29316 23548 29326 23604
rect 34178 23548 34188 23604
rect 34244 23548 36204 23604
rect 36260 23548 36988 23604
rect 37044 23548 37054 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 29036 23436 38892 23492
rect 38948 23436 39788 23492
rect 39844 23436 39854 23492
rect 12786 23324 12796 23380
rect 12852 23324 13580 23380
rect 13636 23324 13646 23380
rect 21186 23212 21196 23268
rect 21252 23212 28812 23268
rect 28868 23212 28878 23268
rect 29036 23156 29092 23436
rect 31602 23324 31612 23380
rect 31668 23324 32396 23380
rect 32452 23324 32462 23380
rect 33058 23324 33068 23380
rect 33124 23324 35644 23380
rect 35700 23324 35710 23380
rect 35970 23324 35980 23380
rect 36036 23324 36988 23380
rect 37044 23324 38668 23380
rect 35644 23268 35700 23324
rect 38612 23268 38668 23324
rect 30370 23212 30380 23268
rect 30436 23212 30884 23268
rect 31042 23212 31052 23268
rect 31108 23212 33404 23268
rect 33460 23212 33964 23268
rect 34020 23212 34030 23268
rect 35644 23212 36092 23268
rect 36148 23212 36158 23268
rect 36530 23212 36540 23268
rect 36596 23212 37884 23268
rect 37940 23212 37950 23268
rect 38612 23212 39900 23268
rect 39956 23212 39966 23268
rect 30828 23156 30884 23212
rect 6402 23100 6412 23156
rect 6468 23100 7756 23156
rect 7812 23100 7822 23156
rect 23986 23100 23996 23156
rect 24052 23100 28476 23156
rect 28532 23100 28542 23156
rect 28812 23100 29092 23156
rect 30034 23100 30044 23156
rect 30100 23100 30604 23156
rect 30660 23100 30670 23156
rect 30828 23100 31724 23156
rect 31780 23100 32396 23156
rect 32452 23100 32462 23156
rect 35858 23100 35868 23156
rect 35924 23100 36764 23156
rect 36820 23100 36830 23156
rect 37762 23100 37772 23156
rect 37828 23100 40684 23156
rect 40740 23100 40750 23156
rect 41570 23100 41580 23156
rect 41636 23100 42812 23156
rect 42868 23100 42878 23156
rect 28812 23044 28868 23100
rect 6066 22988 6076 23044
rect 6132 22988 7196 23044
rect 7252 22988 7262 23044
rect 9202 22988 9212 23044
rect 9268 22988 10892 23044
rect 10948 22988 10958 23044
rect 14578 22988 14588 23044
rect 14644 22988 17836 23044
rect 17892 22988 19292 23044
rect 19348 22988 19358 23044
rect 28802 22988 28812 23044
rect 28868 22988 28878 23044
rect 29026 22988 29036 23044
rect 29092 22988 31612 23044
rect 31668 22988 31678 23044
rect 40338 22988 40348 23044
rect 40404 22988 41692 23044
rect 41748 22988 41758 23044
rect 45200 22932 46000 22960
rect 44146 22876 44156 22932
rect 44212 22876 46000 22932
rect 45200 22848 46000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 11890 22652 11900 22708
rect 11956 22652 12684 22708
rect 12740 22652 12750 22708
rect 28130 22652 28140 22708
rect 28196 22652 34412 22708
rect 34468 22652 34478 22708
rect 36082 22652 36092 22708
rect 36148 22652 36876 22708
rect 36932 22652 36942 22708
rect 10434 22540 10444 22596
rect 10500 22540 13692 22596
rect 13748 22540 13758 22596
rect 6514 22428 6524 22484
rect 6580 22428 18508 22484
rect 18564 22428 18574 22484
rect 27122 22428 27132 22484
rect 27188 22428 27916 22484
rect 27972 22428 27982 22484
rect 4834 22316 4844 22372
rect 4900 22316 5516 22372
rect 5572 22316 5582 22372
rect 7410 22316 7420 22372
rect 7476 22316 10444 22372
rect 10500 22316 10510 22372
rect 11330 22316 11340 22372
rect 11396 22316 12348 22372
rect 12404 22316 12414 22372
rect 12562 22316 12572 22372
rect 12628 22316 21756 22372
rect 21812 22316 22876 22372
rect 22932 22316 22942 22372
rect 12786 22204 12796 22260
rect 12852 22204 15260 22260
rect 15316 22204 15820 22260
rect 15876 22204 15886 22260
rect 23100 22204 26908 22260
rect 26964 22204 27804 22260
rect 27860 22204 27870 22260
rect 23100 22148 23156 22204
rect 28140 22148 28196 22652
rect 35634 22540 35644 22596
rect 35700 22540 37100 22596
rect 37156 22540 38556 22596
rect 38612 22540 38622 22596
rect 31938 22428 31948 22484
rect 32004 22428 33068 22484
rect 33124 22428 33134 22484
rect 34486 22428 34524 22484
rect 34580 22428 34590 22484
rect 40674 22428 40684 22484
rect 40740 22428 42364 22484
rect 42420 22428 42430 22484
rect 34066 22316 34076 22372
rect 34132 22316 35420 22372
rect 35476 22316 35486 22372
rect 35634 22316 35644 22372
rect 35700 22316 35980 22372
rect 36036 22316 36046 22372
rect 37874 22316 37884 22372
rect 37940 22316 39452 22372
rect 39508 22316 39518 22372
rect 28578 22204 28588 22260
rect 28644 22204 29148 22260
rect 29204 22204 29484 22260
rect 29540 22204 30044 22260
rect 30100 22204 30110 22260
rect 34402 22204 34412 22260
rect 34468 22204 37212 22260
rect 37268 22204 37278 22260
rect 10882 22092 10892 22148
rect 10948 22092 13244 22148
rect 13300 22092 13310 22148
rect 19170 22092 19180 22148
rect 19236 22092 20300 22148
rect 20356 22092 20366 22148
rect 22530 22092 22540 22148
rect 22596 22092 23100 22148
rect 23156 22092 23166 22148
rect 26674 22092 26684 22148
rect 26740 22092 28196 22148
rect 35186 22092 35196 22148
rect 35252 22092 37324 22148
rect 37380 22092 37390 22148
rect 27458 21980 27468 22036
rect 27524 21980 29036 22036
rect 29092 21980 29102 22036
rect 31826 21980 31836 22036
rect 31892 21980 35084 22036
rect 35140 21980 35150 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 9202 21868 9212 21924
rect 9268 21868 10668 21924
rect 10724 21868 10734 21924
rect 19030 21868 19068 21924
rect 19124 21868 19134 21924
rect 19618 21868 19628 21924
rect 19684 21868 19694 21924
rect 27794 21868 27804 21924
rect 27860 21868 28700 21924
rect 28756 21868 28766 21924
rect 34178 21868 34188 21924
rect 34244 21868 36428 21924
rect 36484 21868 36494 21924
rect 11554 21756 11564 21812
rect 11620 21756 12460 21812
rect 12516 21756 12526 21812
rect 13682 21756 13692 21812
rect 13748 21756 15484 21812
rect 15540 21756 16492 21812
rect 16548 21756 16558 21812
rect 19628 21700 19684 21868
rect 26338 21756 26348 21812
rect 26404 21756 28140 21812
rect 28196 21756 35868 21812
rect 35924 21756 35934 21812
rect 38546 21756 38556 21812
rect 38612 21756 39788 21812
rect 39844 21756 39854 21812
rect 5282 21644 5292 21700
rect 5348 21644 6636 21700
rect 6692 21644 6702 21700
rect 11666 21644 11676 21700
rect 11732 21644 14476 21700
rect 14532 21644 14542 21700
rect 14690 21644 14700 21700
rect 14756 21644 15932 21700
rect 15988 21644 17724 21700
rect 17780 21644 17790 21700
rect 19058 21644 19068 21700
rect 19124 21644 19684 21700
rect 26786 21644 26796 21700
rect 26852 21644 28588 21700
rect 28644 21644 28654 21700
rect 34738 21644 34748 21700
rect 34804 21644 35196 21700
rect 35252 21644 35262 21700
rect 35634 21644 35644 21700
rect 35700 21644 36540 21700
rect 36596 21644 36606 21700
rect 4386 21532 4396 21588
rect 4452 21532 7756 21588
rect 7812 21532 11788 21588
rect 11844 21532 13916 21588
rect 13972 21532 13982 21588
rect 16370 21532 16380 21588
rect 16436 21532 18732 21588
rect 18788 21532 18798 21588
rect 19394 21532 19404 21588
rect 19460 21532 21532 21588
rect 21588 21532 21598 21588
rect 27682 21532 27692 21588
rect 27748 21532 30828 21588
rect 30884 21532 31724 21588
rect 31780 21532 32396 21588
rect 32452 21532 32462 21588
rect 36642 21532 36652 21588
rect 36708 21532 38108 21588
rect 38164 21532 38174 21588
rect 12338 21420 12348 21476
rect 12404 21420 14364 21476
rect 14420 21420 14430 21476
rect 16706 21420 16716 21476
rect 16772 21420 17500 21476
rect 17556 21420 17566 21476
rect 18162 21420 18172 21476
rect 18228 21420 19964 21476
rect 20020 21420 20030 21476
rect 26852 21420 36540 21476
rect 36596 21420 36606 21476
rect 10882 21308 10892 21364
rect 10948 21308 12012 21364
rect 12068 21308 14140 21364
rect 14196 21308 14206 21364
rect 17266 21308 17276 21364
rect 17332 21308 18620 21364
rect 18676 21308 19292 21364
rect 19348 21308 19740 21364
rect 19796 21308 19806 21364
rect 20178 21308 20188 21364
rect 20244 21308 20524 21364
rect 20580 21308 20590 21364
rect 26852 21252 26908 21420
rect 28578 21308 28588 21364
rect 28644 21308 41020 21364
rect 41076 21308 41086 21364
rect 42242 21308 42252 21364
rect 42308 21308 43372 21364
rect 43428 21308 43438 21364
rect 18946 21196 18956 21252
rect 19012 21196 26908 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 12562 21084 12572 21140
rect 12628 21084 13804 21140
rect 13860 21084 13870 21140
rect 17938 20972 17948 21028
rect 18004 20972 19180 21028
rect 19236 20972 19246 21028
rect 34290 20972 34300 21028
rect 34356 20972 35868 21028
rect 35924 20972 37548 21028
rect 37604 20972 37614 21028
rect 11554 20860 11564 20916
rect 11620 20860 12460 20916
rect 12516 20860 12526 20916
rect 34178 20860 34188 20916
rect 34244 20860 37100 20916
rect 37156 20860 37166 20916
rect 39106 20860 39116 20916
rect 39172 20860 41468 20916
rect 41524 20860 41534 20916
rect 12226 20748 12236 20804
rect 12292 20748 14028 20804
rect 14084 20748 21868 20804
rect 21924 20748 22764 20804
rect 22820 20748 22830 20804
rect 34514 20748 34524 20804
rect 34580 20748 35252 20804
rect 35196 20692 35252 20748
rect 12898 20636 12908 20692
rect 12964 20636 13468 20692
rect 13524 20636 13534 20692
rect 17378 20636 17388 20692
rect 17444 20636 18172 20692
rect 18228 20636 18238 20692
rect 20066 20636 20076 20692
rect 20132 20636 22092 20692
rect 22148 20636 22158 20692
rect 22642 20636 22652 20692
rect 22708 20636 23212 20692
rect 23268 20636 26908 20692
rect 26964 20636 26974 20692
rect 28466 20636 28476 20692
rect 28532 20636 29260 20692
rect 29316 20636 29326 20692
rect 29474 20636 29484 20692
rect 29540 20636 32508 20692
rect 32564 20636 34188 20692
rect 34244 20636 34972 20692
rect 35028 20636 35038 20692
rect 35158 20636 35196 20692
rect 35252 20636 37212 20692
rect 37268 20636 37278 20692
rect 10434 20524 10444 20580
rect 10500 20524 14252 20580
rect 14308 20524 14318 20580
rect 26852 20468 26908 20636
rect 35410 20524 35420 20580
rect 35476 20524 37100 20580
rect 37156 20524 37166 20580
rect 41122 20524 41132 20580
rect 41188 20524 43260 20580
rect 43316 20524 43326 20580
rect 26852 20412 27580 20468
rect 27636 20412 28476 20468
rect 28532 20412 29148 20468
rect 29204 20412 29214 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 29334 20300 29372 20356
rect 29428 20300 29438 20356
rect 14466 20188 14476 20244
rect 14532 20188 15372 20244
rect 15428 20188 15438 20244
rect 19954 20188 19964 20244
rect 20020 20188 20412 20244
rect 20468 20188 20478 20244
rect 25890 20188 25900 20244
rect 25956 20188 26796 20244
rect 26852 20188 26862 20244
rect 29250 20188 29260 20244
rect 29316 20188 29596 20244
rect 29652 20188 29662 20244
rect 35970 20188 35980 20244
rect 36036 20188 36428 20244
rect 36484 20188 36494 20244
rect 4386 20076 4396 20132
rect 4452 20076 5628 20132
rect 5684 20076 5694 20132
rect 8418 20076 8428 20132
rect 8484 20076 11340 20132
rect 11396 20076 11406 20132
rect 12674 20076 12684 20132
rect 12740 20076 13916 20132
rect 13972 20076 13982 20132
rect 19618 20076 19628 20132
rect 19684 20076 20636 20132
rect 20692 20076 20702 20132
rect 27906 20076 27916 20132
rect 27972 20076 28252 20132
rect 28308 20076 29148 20132
rect 29204 20076 29820 20132
rect 29876 20076 29886 20132
rect 32050 20076 32060 20132
rect 32116 20076 33404 20132
rect 33460 20076 33470 20132
rect 34188 20076 35196 20132
rect 35252 20076 37436 20132
rect 37492 20076 37502 20132
rect 39106 20076 39116 20132
rect 39172 20076 40012 20132
rect 40068 20076 40078 20132
rect 40338 20076 40348 20132
rect 40404 20076 40908 20132
rect 40964 20076 40974 20132
rect 43652 20076 43820 20132
rect 43876 20076 43886 20132
rect 4946 19964 4956 20020
rect 5012 19964 11844 20020
rect 12002 19964 12012 20020
rect 12068 19964 14588 20020
rect 14644 19964 14654 20020
rect 17602 19964 17612 20020
rect 17668 19964 18284 20020
rect 18340 19964 18350 20020
rect 30482 19964 30492 20020
rect 30548 19964 31052 20020
rect 31108 19964 32676 20020
rect 32834 19964 32844 20020
rect 32900 19964 33964 20020
rect 34020 19964 34030 20020
rect 11788 19908 11844 19964
rect 32620 19908 32676 19964
rect 34188 19908 34244 20076
rect 35410 19964 35420 20020
rect 35476 19964 36540 20020
rect 36596 19964 36876 20020
rect 36932 19964 36942 20020
rect 37090 19964 37100 20020
rect 37156 19964 38108 20020
rect 38164 19964 39676 20020
rect 39732 19964 39742 20020
rect 42018 19964 42028 20020
rect 42084 19964 42812 20020
rect 42868 19964 42878 20020
rect 2594 19852 2604 19908
rect 2660 19852 4284 19908
rect 4340 19852 11116 19908
rect 11172 19852 11182 19908
rect 11788 19852 13580 19908
rect 13636 19852 13646 19908
rect 14130 19852 14140 19908
rect 14196 19852 15260 19908
rect 15316 19852 15326 19908
rect 31378 19852 31388 19908
rect 31444 19852 32396 19908
rect 32452 19852 32462 19908
rect 32620 19852 34244 19908
rect 34962 19852 34972 19908
rect 35028 19852 37660 19908
rect 37716 19852 37726 19908
rect 13580 19684 13636 19852
rect 43652 19796 43708 20076
rect 13794 19740 13804 19796
rect 13860 19740 19180 19796
rect 19236 19740 20300 19796
rect 20356 19740 20366 19796
rect 30146 19740 30156 19796
rect 30212 19740 43708 19796
rect 13580 19628 14700 19684
rect 14756 19628 14766 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 45200 19572 46000 19600
rect 13122 19516 13132 19572
rect 13188 19516 14812 19572
rect 14868 19516 14878 19572
rect 44258 19516 44268 19572
rect 44324 19516 46000 19572
rect 45200 19488 46000 19516
rect 28690 19404 28700 19460
rect 28756 19404 29204 19460
rect 33394 19404 33404 19460
rect 33460 19404 43708 19460
rect 43764 19404 43774 19460
rect 4946 19292 4956 19348
rect 5012 19292 6076 19348
rect 6132 19292 6524 19348
rect 6580 19292 6590 19348
rect 29148 19236 29204 19404
rect 31154 19292 31164 19348
rect 31220 19292 32060 19348
rect 32116 19292 32126 19348
rect 40226 19292 40236 19348
rect 40292 19292 42252 19348
rect 42308 19292 42318 19348
rect 43652 19292 44044 19348
rect 44100 19292 44110 19348
rect 3266 19180 3276 19236
rect 3332 19180 4844 19236
rect 4900 19180 4910 19236
rect 5058 19180 5068 19236
rect 5124 19180 5964 19236
rect 6020 19180 6030 19236
rect 10994 19180 11004 19236
rect 11060 19180 11900 19236
rect 11956 19180 11966 19236
rect 17042 19180 17052 19236
rect 17108 19180 20188 19236
rect 20244 19180 20254 19236
rect 22306 19180 22316 19236
rect 22372 19180 24220 19236
rect 24276 19180 24286 19236
rect 29138 19180 29148 19236
rect 29204 19180 30044 19236
rect 30100 19180 33292 19236
rect 33348 19180 33358 19236
rect 34738 19180 34748 19236
rect 34804 19180 40684 19236
rect 40740 19180 41244 19236
rect 41300 19180 41310 19236
rect 43652 19124 43708 19292
rect 2034 19068 2044 19124
rect 2100 19068 3164 19124
rect 3220 19068 3230 19124
rect 4610 19068 4620 19124
rect 4676 19068 6636 19124
rect 6692 19068 6702 19124
rect 12114 19068 12124 19124
rect 12180 19068 14140 19124
rect 14196 19068 14206 19124
rect 20962 19068 20972 19124
rect 21028 19068 21980 19124
rect 22036 19068 22046 19124
rect 27906 19068 27916 19124
rect 27972 19068 30156 19124
rect 30212 19068 30222 19124
rect 35634 19068 35644 19124
rect 35700 19068 36428 19124
rect 36484 19068 36494 19124
rect 37650 19068 37660 19124
rect 37716 19068 40236 19124
rect 40292 19068 43708 19124
rect 11106 18956 11116 19012
rect 11172 18956 12348 19012
rect 12404 18956 12414 19012
rect 18498 18956 18508 19012
rect 18564 18956 20748 19012
rect 20804 18956 20814 19012
rect 27570 18956 27580 19012
rect 27636 18956 29708 19012
rect 29764 18956 29774 19012
rect 26114 18844 26124 18900
rect 26180 18844 40796 18900
rect 40852 18844 40862 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 2370 18620 2380 18676
rect 2436 18620 5628 18676
rect 5684 18620 5694 18676
rect 12562 18620 12572 18676
rect 12628 18620 14028 18676
rect 14084 18620 14094 18676
rect 15362 18620 15372 18676
rect 15428 18620 15820 18676
rect 15876 18620 15886 18676
rect 29586 18620 29596 18676
rect 29652 18620 30604 18676
rect 30660 18620 30670 18676
rect 8866 18508 8876 18564
rect 8932 18508 9772 18564
rect 9828 18508 10668 18564
rect 10724 18508 10734 18564
rect 12786 18508 12796 18564
rect 12852 18508 13692 18564
rect 13748 18508 13758 18564
rect 15026 18508 15036 18564
rect 15092 18508 15596 18564
rect 15652 18508 16940 18564
rect 16996 18508 17612 18564
rect 17668 18508 18284 18564
rect 18340 18508 18350 18564
rect 25778 18508 25788 18564
rect 25844 18508 27804 18564
rect 27860 18508 28364 18564
rect 28420 18508 28430 18564
rect 25788 18452 25844 18508
rect 7186 18396 7196 18452
rect 7252 18396 8540 18452
rect 8596 18396 8606 18452
rect 10882 18396 10892 18452
rect 10948 18396 12460 18452
rect 12516 18396 12526 18452
rect 16258 18396 16268 18452
rect 16324 18396 17276 18452
rect 17332 18396 17342 18452
rect 18610 18396 18620 18452
rect 18676 18396 19404 18452
rect 19460 18396 20636 18452
rect 20692 18396 20702 18452
rect 21186 18396 21196 18452
rect 21252 18396 25844 18452
rect 27682 18396 27692 18452
rect 27748 18396 28252 18452
rect 28308 18396 28318 18452
rect 28914 18396 28924 18452
rect 28980 18396 32172 18452
rect 32228 18396 33068 18452
rect 33124 18396 33134 18452
rect 33618 18396 33628 18452
rect 33684 18396 34636 18452
rect 34692 18396 34702 18452
rect 35298 18396 35308 18452
rect 35364 18396 36540 18452
rect 36596 18396 36606 18452
rect 10546 18284 10556 18340
rect 10612 18284 11900 18340
rect 11956 18284 11966 18340
rect 23874 18284 23884 18340
rect 23940 18284 25900 18340
rect 25956 18284 25966 18340
rect 29474 18284 29484 18340
rect 29540 18284 30716 18340
rect 30772 18284 31724 18340
rect 31780 18284 31790 18340
rect 32498 18284 32508 18340
rect 32564 18284 34076 18340
rect 34132 18284 34142 18340
rect 34290 18284 34300 18340
rect 34356 18284 37212 18340
rect 37268 18284 37278 18340
rect 40114 18284 40124 18340
rect 40180 18284 40684 18340
rect 40740 18284 42140 18340
rect 42196 18284 42206 18340
rect 13794 18172 13804 18228
rect 13860 18172 14812 18228
rect 14868 18172 14878 18228
rect 19282 18172 19292 18228
rect 19348 18172 22428 18228
rect 22484 18172 22652 18228
rect 22708 18172 23436 18228
rect 23492 18172 27916 18228
rect 27972 18172 28476 18228
rect 28532 18172 29932 18228
rect 29988 18172 29998 18228
rect 32610 18172 32620 18228
rect 32676 18172 36204 18228
rect 36260 18172 37100 18228
rect 37156 18172 37166 18228
rect 41234 18060 41244 18116
rect 41300 18060 43932 18116
rect 43988 18060 43998 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 19842 17948 19852 18004
rect 19908 17948 21532 18004
rect 21588 17948 21598 18004
rect 14466 17836 14476 17892
rect 14532 17836 16660 17892
rect 18386 17836 18396 17892
rect 18452 17836 27580 17892
rect 27636 17836 27646 17892
rect 5170 17724 5180 17780
rect 5236 17724 5964 17780
rect 6020 17724 9660 17780
rect 9716 17724 9726 17780
rect 11666 17724 11676 17780
rect 11732 17724 13804 17780
rect 13860 17724 13870 17780
rect 14914 17724 14924 17780
rect 14980 17724 15596 17780
rect 15652 17724 15662 17780
rect 16604 17668 16660 17836
rect 18834 17724 18844 17780
rect 18900 17724 18910 17780
rect 26450 17724 26460 17780
rect 26516 17724 26796 17780
rect 26852 17724 28252 17780
rect 28308 17724 28318 17780
rect 33842 17724 33852 17780
rect 33908 17724 37548 17780
rect 37604 17724 38668 17780
rect 14018 17612 14028 17668
rect 14084 17612 16268 17668
rect 16324 17612 16334 17668
rect 16594 17612 16604 17668
rect 16660 17612 16670 17668
rect 6514 17500 6524 17556
rect 6580 17500 7644 17556
rect 7700 17500 7710 17556
rect 18844 17332 18900 17724
rect 38612 17668 38668 17724
rect 20514 17612 20524 17668
rect 20580 17612 21196 17668
rect 21252 17612 21262 17668
rect 26114 17612 26124 17668
rect 26180 17612 27356 17668
rect 27412 17612 27422 17668
rect 33068 17612 35868 17668
rect 35924 17612 35934 17668
rect 38612 17612 38892 17668
rect 38948 17612 38958 17668
rect 33068 17556 33124 17612
rect 21298 17500 21308 17556
rect 21364 17500 22204 17556
rect 22260 17500 22270 17556
rect 24546 17500 24556 17556
rect 24612 17500 33068 17556
rect 33124 17500 33134 17556
rect 34290 17500 34300 17556
rect 34356 17500 35084 17556
rect 35140 17500 35150 17556
rect 36306 17500 36316 17556
rect 36372 17500 36988 17556
rect 37044 17500 37054 17556
rect 28578 17388 28588 17444
rect 28644 17388 29372 17444
rect 29428 17388 29438 17444
rect 31154 17388 31164 17444
rect 31220 17388 32508 17444
rect 32564 17388 33404 17444
rect 33460 17388 33470 17444
rect 18844 17276 19012 17332
rect 18956 17220 19012 17276
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 15092 17164 18732 17220
rect 18788 17164 18798 17220
rect 18946 17164 18956 17220
rect 19012 17164 19628 17220
rect 19684 17164 19694 17220
rect 26114 17164 26124 17220
rect 26180 17164 26796 17220
rect 26852 17164 26862 17220
rect 15092 17108 15148 17164
rect 6066 17052 6076 17108
rect 6132 17052 8204 17108
rect 8260 17052 8270 17108
rect 8978 17052 8988 17108
rect 9044 17052 15148 17108
rect 17826 17052 17836 17108
rect 17892 17052 19068 17108
rect 19124 17052 30828 17108
rect 30884 17052 30894 17108
rect 38882 17052 38892 17108
rect 38948 17052 40348 17108
rect 40404 17052 40414 17108
rect 7186 16940 7196 16996
rect 7252 16940 8316 16996
rect 8372 16940 11900 16996
rect 11956 16940 11966 16996
rect 21634 16940 21644 16996
rect 21700 16940 22876 16996
rect 22932 16940 22942 16996
rect 25666 16940 25676 16996
rect 25732 16940 26124 16996
rect 26180 16940 26190 16996
rect 5282 16828 5292 16884
rect 5348 16828 7084 16884
rect 7140 16828 9324 16884
rect 9380 16828 9492 16884
rect 11778 16828 11788 16884
rect 11844 16828 12460 16884
rect 12516 16828 12526 16884
rect 23986 16828 23996 16884
rect 24052 16828 24062 16884
rect 24770 16828 24780 16884
rect 24836 16828 26796 16884
rect 26852 16828 26862 16884
rect 27346 16828 27356 16884
rect 27412 16828 28476 16884
rect 28532 16828 28542 16884
rect 29922 16828 29932 16884
rect 29988 16828 30716 16884
rect 30772 16828 30782 16884
rect 34300 16828 35532 16884
rect 35588 16828 35598 16884
rect 43586 16828 43596 16884
rect 43652 16828 44156 16884
rect 44212 16828 45332 16884
rect 9436 16772 9492 16828
rect 23996 16772 24052 16828
rect 34300 16772 34356 16828
rect 9436 16716 10332 16772
rect 10388 16716 10398 16772
rect 10658 16716 10668 16772
rect 10724 16716 13132 16772
rect 13188 16716 13198 16772
rect 14578 16716 14588 16772
rect 14644 16716 16828 16772
rect 16884 16716 16894 16772
rect 22306 16716 22316 16772
rect 22372 16716 22988 16772
rect 23044 16716 23054 16772
rect 23996 16716 24220 16772
rect 24276 16716 26908 16772
rect 26964 16716 27580 16772
rect 27636 16716 27646 16772
rect 29138 16716 29148 16772
rect 29204 16716 29484 16772
rect 29540 16716 29550 16772
rect 34290 16716 34300 16772
rect 34356 16716 34366 16772
rect 35746 16716 35756 16772
rect 35812 16716 36540 16772
rect 36596 16716 36606 16772
rect 10434 16604 10444 16660
rect 10500 16604 11340 16660
rect 11396 16604 11406 16660
rect 14242 16604 14252 16660
rect 14308 16604 22428 16660
rect 22484 16604 22494 16660
rect 45276 16548 45332 16828
rect 20178 16492 20188 16548
rect 20244 16492 21756 16548
rect 21812 16492 21822 16548
rect 21970 16492 21980 16548
rect 22036 16492 29148 16548
rect 29204 16492 29214 16548
rect 45052 16492 45332 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 21980 16436 22036 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 16594 16380 16604 16436
rect 16660 16380 17276 16436
rect 17332 16380 20300 16436
rect 20356 16380 22036 16436
rect 15922 16268 15932 16324
rect 15988 16268 17500 16324
rect 17556 16268 17566 16324
rect 20626 16268 20636 16324
rect 20692 16268 23100 16324
rect 23156 16268 27020 16324
rect 27076 16268 27086 16324
rect 28130 16268 28140 16324
rect 28196 16268 28588 16324
rect 28644 16268 28654 16324
rect 30818 16268 30828 16324
rect 30884 16268 31948 16324
rect 32004 16268 33068 16324
rect 33124 16268 43820 16324
rect 43876 16268 43886 16324
rect 45052 16212 45108 16492
rect 45200 16212 46000 16240
rect 11218 16156 11228 16212
rect 11284 16156 12124 16212
rect 12180 16156 12190 16212
rect 12450 16156 12460 16212
rect 12516 16156 14252 16212
rect 14308 16156 14318 16212
rect 19954 16156 19964 16212
rect 20020 16156 21308 16212
rect 21364 16156 21374 16212
rect 26674 16156 26684 16212
rect 26740 16156 29708 16212
rect 29764 16156 30604 16212
rect 30660 16156 30670 16212
rect 45052 16156 46000 16212
rect 45200 16128 46000 16156
rect 10546 16044 10556 16100
rect 10612 16044 15148 16100
rect 15204 16044 19068 16100
rect 19124 16044 19134 16100
rect 20066 16044 20076 16100
rect 20132 16044 21868 16100
rect 21924 16044 21934 16100
rect 23090 16044 23100 16100
rect 23156 16044 23884 16100
rect 23940 16044 25340 16100
rect 25396 16044 25406 16100
rect 25778 16044 25788 16100
rect 25844 16044 27524 16100
rect 27682 16044 27692 16100
rect 27748 16044 29484 16100
rect 29540 16044 29550 16100
rect 40002 16044 40012 16100
rect 40068 16044 42028 16100
rect 42084 16044 42094 16100
rect 23100 15988 23156 16044
rect 27468 15988 27524 16044
rect 9538 15932 9548 15988
rect 9604 15932 10220 15988
rect 10276 15932 11900 15988
rect 11956 15932 11966 15988
rect 14130 15932 14140 15988
rect 14196 15932 14812 15988
rect 14868 15932 14878 15988
rect 21522 15932 21532 15988
rect 21588 15932 23156 15988
rect 24322 15932 24332 15988
rect 24388 15932 24892 15988
rect 24948 15932 26908 15988
rect 27468 15932 28140 15988
rect 28196 15932 28206 15988
rect 30034 15932 30044 15988
rect 30100 15932 30110 15988
rect 26852 15876 26908 15932
rect 30044 15876 30100 15932
rect 8754 15820 8764 15876
rect 8820 15820 9436 15876
rect 9492 15820 10108 15876
rect 10164 15820 10174 15876
rect 12226 15820 12236 15876
rect 12292 15820 13804 15876
rect 13860 15820 13870 15876
rect 20514 15820 20524 15876
rect 20580 15820 22316 15876
rect 22372 15820 22382 15876
rect 26852 15820 28700 15876
rect 28756 15820 30100 15876
rect 30370 15820 30380 15876
rect 30436 15820 31612 15876
rect 31668 15820 34300 15876
rect 34356 15820 34366 15876
rect 19030 15708 19068 15764
rect 19124 15708 19134 15764
rect 26898 15708 26908 15764
rect 26964 15708 28476 15764
rect 28532 15708 28542 15764
rect 30706 15708 30716 15764
rect 30772 15708 32956 15764
rect 33012 15708 35532 15764
rect 35588 15708 35598 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 22530 15596 22540 15652
rect 22596 15596 24220 15652
rect 24276 15596 26348 15652
rect 26404 15596 26414 15652
rect 26852 15596 31052 15652
rect 31108 15596 31388 15652
rect 31444 15596 31454 15652
rect 26852 15540 26908 15596
rect 11106 15484 11116 15540
rect 11172 15484 13132 15540
rect 13188 15484 13198 15540
rect 14130 15484 14140 15540
rect 14196 15484 14588 15540
rect 14644 15484 16604 15540
rect 16660 15484 16670 15540
rect 17714 15484 17724 15540
rect 17780 15484 26908 15540
rect 28130 15484 28140 15540
rect 28196 15484 31276 15540
rect 31332 15484 31342 15540
rect 39778 15484 39788 15540
rect 39844 15484 40908 15540
rect 40964 15484 40974 15540
rect 8978 15372 8988 15428
rect 9044 15372 12236 15428
rect 12292 15372 13356 15428
rect 13412 15372 13422 15428
rect 18498 15372 18508 15428
rect 18564 15372 19404 15428
rect 19460 15372 19470 15428
rect 20850 15372 20860 15428
rect 20916 15372 21420 15428
rect 21476 15372 21486 15428
rect 22306 15372 22316 15428
rect 22372 15372 25228 15428
rect 25284 15372 25294 15428
rect 25442 15372 25452 15428
rect 25508 15372 26348 15428
rect 26404 15372 26908 15428
rect 26964 15372 26974 15428
rect 27122 15372 27132 15428
rect 27188 15372 27692 15428
rect 27748 15372 27758 15428
rect 28802 15372 28812 15428
rect 28868 15372 30380 15428
rect 30436 15372 30446 15428
rect 30930 15372 30940 15428
rect 30996 15372 31388 15428
rect 31444 15372 31454 15428
rect 40226 15372 40236 15428
rect 40292 15372 41132 15428
rect 41188 15372 41198 15428
rect 8418 15260 8428 15316
rect 8484 15260 13468 15316
rect 13524 15260 13534 15316
rect 19506 15260 19516 15316
rect 19572 15260 21532 15316
rect 21588 15260 21598 15316
rect 26226 15260 26236 15316
rect 26292 15260 26908 15316
rect 27010 15260 27020 15316
rect 27076 15260 27916 15316
rect 27972 15260 28476 15316
rect 28532 15260 28542 15316
rect 29334 15260 29372 15316
rect 29428 15260 30044 15316
rect 30100 15260 30110 15316
rect 39890 15260 39900 15316
rect 39956 15260 40796 15316
rect 40852 15260 43484 15316
rect 43540 15260 43550 15316
rect 26852 15204 26908 15260
rect 10322 15148 10332 15204
rect 10388 15148 13244 15204
rect 13300 15148 13310 15204
rect 19618 15148 19628 15204
rect 19684 15148 20636 15204
rect 20692 15148 20702 15204
rect 22866 15148 22876 15204
rect 22932 15148 24444 15204
rect 24500 15148 24510 15204
rect 26852 15148 27132 15204
rect 27188 15148 27198 15204
rect 27794 15148 27804 15204
rect 27860 15148 28588 15204
rect 28644 15148 28654 15204
rect 36530 15148 36540 15204
rect 36596 15148 39228 15204
rect 39284 15148 39676 15204
rect 39732 15148 39742 15204
rect 25666 15036 25676 15092
rect 25732 15036 26796 15092
rect 26852 15036 26862 15092
rect 32050 15036 32060 15092
rect 32116 15036 34076 15092
rect 34132 15036 34142 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 18834 14700 18844 14756
rect 18900 14700 19516 14756
rect 19572 14700 19582 14756
rect 24434 14700 24444 14756
rect 24500 14700 26012 14756
rect 26068 14700 26078 14756
rect 26450 14700 26460 14756
rect 26516 14700 28364 14756
rect 28420 14700 28430 14756
rect 19058 14588 19068 14644
rect 19124 14588 20076 14644
rect 20132 14588 23772 14644
rect 23828 14588 23838 14644
rect 25442 14588 25452 14644
rect 25508 14588 25788 14644
rect 25844 14588 25854 14644
rect 28242 14588 28252 14644
rect 28308 14588 28812 14644
rect 28868 14588 28878 14644
rect 22642 14476 22652 14532
rect 22708 14476 24556 14532
rect 24612 14476 24622 14532
rect 25340 14476 26908 14532
rect 27794 14476 27804 14532
rect 27860 14476 27870 14532
rect 29110 14476 29148 14532
rect 29204 14476 30716 14532
rect 30772 14476 30782 14532
rect 41234 14476 41244 14532
rect 41300 14476 42028 14532
rect 42084 14476 42094 14532
rect 25340 14308 25396 14476
rect 26852 14420 26908 14476
rect 27804 14420 27860 14476
rect 26114 14364 26124 14420
rect 26180 14364 26190 14420
rect 26852 14364 27860 14420
rect 26124 14308 26180 14364
rect 12786 14252 12796 14308
rect 12852 14252 14812 14308
rect 14868 14252 14878 14308
rect 15698 14252 15708 14308
rect 15764 14252 17164 14308
rect 17220 14252 17230 14308
rect 18162 14252 18172 14308
rect 18228 14252 18620 14308
rect 18676 14252 18686 14308
rect 18806 14252 18844 14308
rect 18900 14252 18910 14308
rect 22194 14252 22204 14308
rect 22260 14252 23660 14308
rect 23716 14252 25340 14308
rect 25396 14252 25406 14308
rect 26124 14252 27020 14308
rect 27076 14252 27086 14308
rect 30258 14252 30268 14308
rect 30324 14252 41244 14308
rect 41300 14252 42700 14308
rect 42756 14252 42766 14308
rect 15932 14084 15988 14252
rect 20188 14140 29596 14196
rect 29652 14140 29662 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 15922 14028 15932 14084
rect 15988 14028 15998 14084
rect 20188 13972 20244 14140
rect 17490 13916 17500 13972
rect 17556 13916 20244 13972
rect 21970 13916 21980 13972
rect 22036 13916 23436 13972
rect 23492 13916 27132 13972
rect 27188 13916 28364 13972
rect 28420 13916 28430 13972
rect 31266 13916 31276 13972
rect 31332 13916 31836 13972
rect 31892 13916 33068 13972
rect 33124 13916 35084 13972
rect 35140 13916 35150 13972
rect 39106 13916 39116 13972
rect 39172 13916 39788 13972
rect 39844 13916 39854 13972
rect 15362 13804 15372 13860
rect 15428 13804 16492 13860
rect 16548 13804 20300 13860
rect 20356 13804 20366 13860
rect 31490 13804 31500 13860
rect 31556 13804 32060 13860
rect 32116 13804 32452 13860
rect 32610 13804 32620 13860
rect 32676 13804 33404 13860
rect 33460 13804 34188 13860
rect 34244 13804 34254 13860
rect 32396 13748 32452 13804
rect 9090 13692 9100 13748
rect 9156 13692 9884 13748
rect 9940 13692 10892 13748
rect 10948 13692 10958 13748
rect 13346 13692 13356 13748
rect 13412 13692 18788 13748
rect 18946 13692 18956 13748
rect 19012 13692 19292 13748
rect 19348 13692 20412 13748
rect 20468 13692 20478 13748
rect 20850 13692 20860 13748
rect 20916 13692 22204 13748
rect 22260 13692 22270 13748
rect 26562 13692 26572 13748
rect 26628 13692 27132 13748
rect 27188 13692 27198 13748
rect 31266 13692 31276 13748
rect 31332 13692 31724 13748
rect 31780 13692 31948 13748
rect 32004 13692 32014 13748
rect 32396 13692 32956 13748
rect 33012 13692 33022 13748
rect 40338 13692 40348 13748
rect 40404 13692 41244 13748
rect 41300 13692 41310 13748
rect 13580 13636 13636 13692
rect 18732 13636 18788 13692
rect 13570 13580 13580 13636
rect 13636 13580 13646 13636
rect 13794 13580 13804 13636
rect 13860 13580 15148 13636
rect 15204 13580 15214 13636
rect 15474 13580 15484 13636
rect 15540 13580 18060 13636
rect 18116 13580 18126 13636
rect 18732 13580 19628 13636
rect 19684 13580 19852 13636
rect 19908 13580 19918 13636
rect 24770 13580 24780 13636
rect 24836 13580 25228 13636
rect 25284 13580 26908 13636
rect 26964 13580 26974 13636
rect 41794 13580 41804 13636
rect 41860 13580 42364 13636
rect 42420 13580 43148 13636
rect 43204 13580 43214 13636
rect 12338 13468 12348 13524
rect 12404 13468 13356 13524
rect 13412 13468 14140 13524
rect 14196 13468 14206 13524
rect 14354 13468 14364 13524
rect 14420 13468 15596 13524
rect 15652 13468 15662 13524
rect 33170 13468 33180 13524
rect 33236 13468 35420 13524
rect 35476 13468 35486 13524
rect 26852 13356 29820 13412
rect 29876 13356 29886 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 26852 13188 26908 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 36642 13244 36652 13300
rect 36708 13244 37436 13300
rect 37492 13244 37502 13300
rect 18050 13132 18060 13188
rect 18116 13132 19404 13188
rect 19460 13132 19470 13188
rect 20066 13132 20076 13188
rect 20132 13132 22988 13188
rect 23044 13132 26908 13188
rect 34514 13132 34524 13188
rect 34580 13132 36988 13188
rect 37044 13132 37054 13188
rect 19170 13020 19180 13076
rect 19236 13020 20188 13076
rect 20244 13020 20636 13076
rect 20692 13020 20702 13076
rect 28802 13020 28812 13076
rect 28868 13020 30044 13076
rect 30100 13020 30110 13076
rect 36754 13020 36764 13076
rect 36820 13020 37548 13076
rect 37604 13020 38220 13076
rect 38276 13020 39676 13076
rect 39732 13020 39742 13076
rect 32834 12908 32844 12964
rect 32900 12908 33516 12964
rect 33572 12908 33582 12964
rect 45200 12852 46000 12880
rect 11666 12796 11676 12852
rect 11732 12796 12460 12852
rect 12516 12796 12526 12852
rect 27234 12796 27244 12852
rect 27300 12796 28140 12852
rect 28196 12796 28206 12852
rect 36418 12796 36428 12852
rect 36484 12796 37100 12852
rect 37156 12796 37166 12852
rect 44146 12796 44156 12852
rect 44212 12796 46000 12852
rect 45200 12768 46000 12796
rect 18498 12684 18508 12740
rect 18564 12684 18574 12740
rect 22866 12684 22876 12740
rect 22932 12684 31500 12740
rect 31556 12684 31566 12740
rect 38882 12684 38892 12740
rect 38948 12684 41692 12740
rect 41748 12684 41758 12740
rect 16706 12348 16716 12404
rect 16772 12348 17500 12404
rect 17556 12348 17566 12404
rect 18508 12292 18564 12684
rect 28578 12572 28588 12628
rect 28644 12572 43708 12628
rect 43764 12572 43774 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 33954 12460 33964 12516
rect 34020 12460 36540 12516
rect 36596 12460 36606 12516
rect 21746 12348 21756 12404
rect 21812 12348 22092 12404
rect 22148 12348 22158 12404
rect 22978 12348 22988 12404
rect 23044 12348 23660 12404
rect 23716 12348 23726 12404
rect 34066 12348 34076 12404
rect 34132 12348 36316 12404
rect 36372 12348 38780 12404
rect 38836 12348 38846 12404
rect 18386 12236 18396 12292
rect 18452 12236 19852 12292
rect 19908 12236 28812 12292
rect 28868 12236 28878 12292
rect 30930 12236 30940 12292
rect 30996 12236 36148 12292
rect 41794 12236 41804 12292
rect 41860 12236 43260 12292
rect 43316 12236 43326 12292
rect 27906 12124 27916 12180
rect 27972 12124 28588 12180
rect 28644 12124 28654 12180
rect 16818 12012 16828 12068
rect 16884 12012 17612 12068
rect 17668 12012 17678 12068
rect 32386 12012 32396 12068
rect 32452 12012 33852 12068
rect 33908 12012 33918 12068
rect 36092 11844 36148 12236
rect 36082 11788 36092 11844
rect 36148 11788 36158 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 22418 11676 22428 11732
rect 22484 11676 22764 11732
rect 22820 11676 22830 11732
rect 19058 11564 19068 11620
rect 19124 11564 19628 11620
rect 19684 11564 21196 11620
rect 21252 11564 21262 11620
rect 21746 11564 21756 11620
rect 21812 11564 22092 11620
rect 22148 11564 22158 11620
rect 22316 11564 27692 11620
rect 27748 11564 30268 11620
rect 30324 11564 30334 11620
rect 32946 11564 32956 11620
rect 33012 11564 38220 11620
rect 38276 11564 38556 11620
rect 38612 11564 38622 11620
rect 22316 11508 22372 11564
rect 15092 11452 20748 11508
rect 20804 11452 21532 11508
rect 21588 11452 22372 11508
rect 24546 11452 24556 11508
rect 24612 11452 25676 11508
rect 25732 11452 25742 11508
rect 32834 11452 32844 11508
rect 32900 11452 33852 11508
rect 33908 11452 33918 11508
rect 35970 11452 35980 11508
rect 36036 11452 38108 11508
rect 38164 11452 38444 11508
rect 38500 11452 38510 11508
rect 15092 11172 15148 11452
rect 15810 11340 15820 11396
rect 15876 11340 22428 11396
rect 22484 11340 22494 11396
rect 22754 11340 22764 11396
rect 22820 11340 23996 11396
rect 24052 11340 24062 11396
rect 28018 11340 28028 11396
rect 28084 11340 29820 11396
rect 29876 11340 29886 11396
rect 35522 11340 35532 11396
rect 35588 11340 36764 11396
rect 36820 11340 37772 11396
rect 37828 11340 37838 11396
rect 38322 11340 38332 11396
rect 38388 11340 39228 11396
rect 39284 11340 39294 11396
rect 26562 11228 26572 11284
rect 26628 11228 27356 11284
rect 27412 11228 27422 11284
rect 29474 11228 29484 11284
rect 29540 11228 32620 11284
rect 32676 11228 33516 11284
rect 33572 11228 33582 11284
rect 12226 11116 12236 11172
rect 12292 11116 12796 11172
rect 12852 11116 13356 11172
rect 13412 11116 15148 11172
rect 22194 11116 22204 11172
rect 22260 11116 23996 11172
rect 24052 11116 24062 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 13122 10892 13132 10948
rect 13188 10892 15372 10948
rect 15428 10892 15438 10948
rect 34860 10892 36316 10948
rect 36372 10892 36382 10948
rect 34860 10836 34916 10892
rect 15250 10780 15260 10836
rect 15316 10780 15820 10836
rect 15876 10780 15886 10836
rect 32274 10780 32284 10836
rect 32340 10780 34860 10836
rect 34916 10780 34926 10836
rect 35308 10780 37548 10836
rect 37604 10780 37614 10836
rect 35308 10724 35364 10780
rect 10994 10668 11004 10724
rect 11060 10668 11900 10724
rect 11956 10668 12348 10724
rect 12404 10668 12796 10724
rect 12852 10668 13804 10724
rect 13860 10668 13870 10724
rect 21410 10668 21420 10724
rect 21476 10668 22204 10724
rect 22260 10668 23212 10724
rect 23268 10668 23278 10724
rect 31042 10668 31052 10724
rect 31108 10668 31724 10724
rect 31780 10668 35308 10724
rect 35364 10668 35374 10724
rect 36530 10668 36540 10724
rect 36596 10668 37436 10724
rect 37492 10668 37502 10724
rect 27682 10556 27692 10612
rect 27748 10556 29148 10612
rect 29204 10556 29214 10612
rect 35074 10556 35084 10612
rect 35140 10556 35150 10612
rect 36978 10556 36988 10612
rect 37044 10556 38332 10612
rect 38388 10556 38398 10612
rect 35084 10500 35140 10556
rect 29922 10444 29932 10500
rect 29988 10444 30940 10500
rect 30996 10444 31006 10500
rect 34738 10444 34748 10500
rect 34804 10444 39844 10500
rect 35522 10332 35532 10388
rect 35588 10332 38220 10388
rect 38276 10332 38286 10388
rect 39788 10276 39844 10444
rect 20962 10220 20972 10276
rect 21028 10220 21420 10276
rect 21476 10220 21486 10276
rect 39778 10220 39788 10276
rect 39844 10220 41804 10276
rect 41860 10220 44044 10276
rect 44100 10220 44110 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 18722 10108 18732 10164
rect 18788 10108 19516 10164
rect 19572 10108 19582 10164
rect 20626 10108 20636 10164
rect 20692 10108 22092 10164
rect 22148 10108 22158 10164
rect 21858 9996 21868 10052
rect 21924 9996 22428 10052
rect 22484 9996 22988 10052
rect 23044 9996 23054 10052
rect 30482 9996 30492 10052
rect 30548 9996 31948 10052
rect 34514 9996 34524 10052
rect 34580 9996 36316 10052
rect 36372 9996 36382 10052
rect 31892 9940 31948 9996
rect 16146 9884 16156 9940
rect 16212 9884 18844 9940
rect 18900 9884 19516 9940
rect 19572 9884 19582 9940
rect 31892 9884 38668 9940
rect 38724 9884 38734 9940
rect 9426 9772 9436 9828
rect 9492 9772 12460 9828
rect 12516 9772 13468 9828
rect 13524 9772 13534 9828
rect 35970 9772 35980 9828
rect 36036 9772 38108 9828
rect 38164 9772 38174 9828
rect 40674 9772 40684 9828
rect 40740 9772 42364 9828
rect 42420 9772 42430 9828
rect 12786 9660 12796 9716
rect 12852 9660 13580 9716
rect 13636 9660 13646 9716
rect 17490 9660 17500 9716
rect 17556 9660 18396 9716
rect 18452 9660 18462 9716
rect 18610 9660 18620 9716
rect 18676 9660 20636 9716
rect 20692 9660 20702 9716
rect 22754 9660 22764 9716
rect 22820 9660 26908 9716
rect 26964 9660 26974 9716
rect 30594 9548 30604 9604
rect 30660 9548 31388 9604
rect 31444 9548 32508 9604
rect 32564 9548 32574 9604
rect 45200 9492 46000 9520
rect 34514 9436 34524 9492
rect 34580 9436 38444 9492
rect 38500 9436 38510 9492
rect 43362 9436 43372 9492
rect 43428 9436 44156 9492
rect 44212 9436 46000 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 45200 9408 46000 9436
rect 27794 9324 27804 9380
rect 27860 9324 43708 9380
rect 43764 9324 43774 9380
rect 11218 9212 11228 9268
rect 11284 9212 12796 9268
rect 12852 9212 12862 9268
rect 14354 9212 14364 9268
rect 14420 9212 15820 9268
rect 15876 9212 15886 9268
rect 35074 9212 35084 9268
rect 35140 9212 37212 9268
rect 37268 9212 37278 9268
rect 24322 9100 24332 9156
rect 24388 9100 25340 9156
rect 25396 9100 25788 9156
rect 25844 9100 25854 9156
rect 29026 9100 29036 9156
rect 29092 9100 30940 9156
rect 30996 9100 31724 9156
rect 31780 9100 31790 9156
rect 34290 9100 34300 9156
rect 34356 9100 35868 9156
rect 35924 9100 35934 9156
rect 41010 9100 41020 9156
rect 41076 9100 42028 9156
rect 42084 9100 42094 9156
rect 13122 8988 13132 9044
rect 13188 8988 15260 9044
rect 15316 8988 15326 9044
rect 34178 8988 34188 9044
rect 34244 8988 36652 9044
rect 36708 8988 36718 9044
rect 37762 8988 37772 9044
rect 37828 8988 38556 9044
rect 38612 8988 40684 9044
rect 40740 8988 40750 9044
rect 13234 8876 13244 8932
rect 13300 8876 13804 8932
rect 13860 8876 16044 8932
rect 16100 8876 16110 8932
rect 19058 8876 19068 8932
rect 19124 8876 19740 8932
rect 19796 8876 19806 8932
rect 28466 8876 28476 8932
rect 28532 8876 29820 8932
rect 29876 8876 37212 8932
rect 37268 8876 37996 8932
rect 38052 8876 38062 8932
rect 39442 8876 39452 8932
rect 39508 8876 42140 8932
rect 42196 8876 42206 8932
rect 15586 8764 15596 8820
rect 15652 8764 18956 8820
rect 19012 8764 19022 8820
rect 20402 8764 20412 8820
rect 20468 8764 22652 8820
rect 22708 8764 24220 8820
rect 24276 8764 24286 8820
rect 35746 8764 35756 8820
rect 35812 8764 36988 8820
rect 37044 8764 37054 8820
rect 39452 8708 39508 8876
rect 12114 8652 12124 8708
rect 12180 8652 14140 8708
rect 14196 8652 14206 8708
rect 14914 8652 14924 8708
rect 14980 8652 22540 8708
rect 22596 8652 22606 8708
rect 23314 8652 23324 8708
rect 23380 8652 23772 8708
rect 23828 8652 23838 8708
rect 36306 8652 36316 8708
rect 36372 8652 36876 8708
rect 36932 8652 39508 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 21298 8540 21308 8596
rect 21364 8540 22764 8596
rect 22820 8540 22830 8596
rect 19618 8428 19628 8484
rect 19684 8428 20580 8484
rect 22838 8428 22876 8484
rect 22932 8428 22942 8484
rect 41010 8428 41020 8484
rect 41076 8428 41086 8484
rect 42018 8428 42028 8484
rect 42084 8428 42812 8484
rect 42868 8428 42878 8484
rect 20524 8372 20580 8428
rect 41020 8372 41076 8428
rect 9538 8316 9548 8372
rect 9604 8316 11228 8372
rect 11284 8316 11900 8372
rect 11956 8316 11966 8372
rect 18722 8316 18732 8372
rect 18788 8316 20300 8372
rect 20356 8316 20366 8372
rect 20524 8316 29260 8372
rect 29316 8316 30044 8372
rect 30100 8316 30110 8372
rect 38882 8316 38892 8372
rect 38948 8316 43372 8372
rect 43428 8316 43438 8372
rect 11330 8204 11340 8260
rect 11396 8204 12012 8260
rect 12068 8204 13692 8260
rect 13748 8204 13758 8260
rect 19506 8204 19516 8260
rect 19572 8204 21420 8260
rect 21476 8204 21486 8260
rect 21634 8204 21644 8260
rect 21700 8204 25116 8260
rect 25172 8204 25564 8260
rect 25620 8204 26908 8260
rect 35298 8204 35308 8260
rect 35364 8204 35868 8260
rect 35924 8204 38668 8260
rect 38724 8204 38734 8260
rect 42242 8204 42252 8260
rect 42308 8204 43148 8260
rect 43204 8204 43214 8260
rect 10882 8092 10892 8148
rect 10948 8092 13020 8148
rect 13076 8092 13086 8148
rect 13458 8092 13468 8148
rect 13524 8092 15820 8148
rect 15876 8092 15886 8148
rect 17042 8092 17052 8148
rect 17108 8092 25788 8148
rect 25844 8092 25854 8148
rect 12348 8036 12404 8092
rect 9314 7980 9324 8036
rect 9380 7980 10780 8036
rect 10836 7980 12124 8036
rect 12180 7980 12190 8036
rect 12338 7980 12348 8036
rect 12404 7980 12414 8036
rect 17378 7980 17388 8036
rect 17444 7980 18620 8036
rect 18676 7980 18686 8036
rect 19282 7980 19292 8036
rect 19348 7980 19740 8036
rect 19796 7980 19806 8036
rect 20738 7980 20748 8036
rect 20804 7980 21532 8036
rect 21588 7980 22316 8036
rect 22372 7980 22382 8036
rect 22530 7980 22540 8036
rect 22596 7980 22606 8036
rect 22754 7980 22764 8036
rect 22820 7980 23324 8036
rect 23380 7980 23390 8036
rect 17602 7868 17612 7924
rect 17668 7868 18508 7924
rect 18564 7868 18574 7924
rect 20178 7868 20188 7924
rect 20244 7868 21644 7924
rect 21700 7868 21710 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 22540 7812 22596 7980
rect 26852 7924 26908 8204
rect 31042 7980 31052 8036
rect 31108 7980 34076 8036
rect 34132 7980 34748 8036
rect 34804 7980 34814 8036
rect 41794 7980 41804 8036
rect 41860 7980 43036 8036
rect 43092 7980 43102 8036
rect 26852 7868 28812 7924
rect 28868 7868 28878 7924
rect 34850 7868 34860 7924
rect 34916 7868 35756 7924
rect 35812 7868 35822 7924
rect 15922 7756 15932 7812
rect 15988 7756 19516 7812
rect 19572 7756 19582 7812
rect 22540 7756 22764 7812
rect 22820 7756 22830 7812
rect 35634 7756 35644 7812
rect 35700 7756 37436 7812
rect 37492 7756 39004 7812
rect 39060 7756 40908 7812
rect 40964 7756 40974 7812
rect 24658 7644 24668 7700
rect 24724 7644 25228 7700
rect 25284 7644 25294 7700
rect 30370 7644 30380 7700
rect 30436 7644 31948 7700
rect 32004 7644 32396 7700
rect 32452 7644 32462 7700
rect 33282 7644 33292 7700
rect 33348 7644 35868 7700
rect 35924 7644 35934 7700
rect 39890 7644 39900 7700
rect 39956 7644 43596 7700
rect 43652 7644 43662 7700
rect 19058 7532 19068 7588
rect 19124 7532 22092 7588
rect 22148 7532 22158 7588
rect 22866 7532 22876 7588
rect 22932 7532 24556 7588
rect 24612 7532 24622 7588
rect 32610 7532 32620 7588
rect 32676 7532 33516 7588
rect 33572 7532 33582 7588
rect 16818 7420 16828 7476
rect 16884 7420 19964 7476
rect 20020 7420 20030 7476
rect 22306 7420 22316 7476
rect 22372 7420 24892 7476
rect 24948 7420 25228 7476
rect 25284 7420 25294 7476
rect 34066 7420 34076 7476
rect 34132 7420 34972 7476
rect 35028 7420 35038 7476
rect 16706 7308 16716 7364
rect 16772 7308 19292 7364
rect 19348 7308 19358 7364
rect 19506 7308 19516 7364
rect 19572 7308 19852 7364
rect 19908 7308 19918 7364
rect 32946 7308 32956 7364
rect 33012 7308 33964 7364
rect 34020 7308 34030 7364
rect 31378 7196 31388 7252
rect 31444 7196 31948 7252
rect 32004 7196 35308 7252
rect 35364 7196 35374 7252
rect 36418 7196 36428 7252
rect 36484 7196 40460 7252
rect 40516 7196 41020 7252
rect 41076 7196 41086 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 12114 6860 12124 6916
rect 12180 6860 16716 6916
rect 16772 6860 16782 6916
rect 12674 6748 12684 6804
rect 12740 6748 13468 6804
rect 13524 6748 14028 6804
rect 14084 6748 14094 6804
rect 18386 6748 18396 6804
rect 18452 6748 19628 6804
rect 19684 6748 19694 6804
rect 24546 6748 24556 6804
rect 24612 6748 25900 6804
rect 25956 6748 28588 6804
rect 28644 6748 28654 6804
rect 34290 6748 34300 6804
rect 34356 6748 36204 6804
rect 36260 6748 36270 6804
rect 11218 6636 11228 6692
rect 11284 6636 12572 6692
rect 12628 6636 12638 6692
rect 18050 6636 18060 6692
rect 18116 6636 20300 6692
rect 20356 6636 20366 6692
rect 21410 6636 21420 6692
rect 21476 6636 22764 6692
rect 22820 6636 22830 6692
rect 32386 6636 32396 6692
rect 32452 6636 33292 6692
rect 33348 6636 33358 6692
rect 35186 6636 35196 6692
rect 35252 6636 36988 6692
rect 37044 6636 37772 6692
rect 37828 6636 37838 6692
rect 39554 6636 39564 6692
rect 39620 6636 43820 6692
rect 43876 6636 43886 6692
rect 20300 6580 20356 6636
rect 20300 6524 22428 6580
rect 22484 6524 22494 6580
rect 33170 6524 33180 6580
rect 33236 6524 34076 6580
rect 34132 6524 34142 6580
rect 11778 6412 11788 6468
rect 11844 6412 12236 6468
rect 12292 6412 12302 6468
rect 13906 6412 13916 6468
rect 13972 6412 16492 6468
rect 16548 6412 17388 6468
rect 17444 6412 17454 6468
rect 24322 6412 24332 6468
rect 24388 6412 26908 6468
rect 26964 6412 26974 6468
rect 28130 6412 28140 6468
rect 28196 6412 29148 6468
rect 29204 6412 29214 6468
rect 32610 6412 32620 6468
rect 32676 6412 36092 6468
rect 36148 6412 36158 6468
rect 34402 6300 34412 6356
rect 34468 6300 34860 6356
rect 34916 6300 37436 6356
rect 37492 6300 40348 6356
rect 40404 6300 40414 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 45200 6132 46000 6160
rect 8866 6076 8876 6132
rect 8932 6076 13132 6132
rect 13188 6076 13198 6132
rect 18806 6076 18844 6132
rect 18900 6076 18910 6132
rect 22754 6076 22764 6132
rect 22820 6076 23772 6132
rect 23828 6076 23838 6132
rect 31892 6076 32620 6132
rect 32676 6076 32686 6132
rect 33282 6076 33292 6132
rect 33348 6076 34188 6132
rect 34244 6076 35532 6132
rect 35588 6076 35598 6132
rect 41458 6076 41468 6132
rect 41524 6076 42140 6132
rect 42196 6076 42206 6132
rect 43586 6076 43596 6132
rect 43652 6076 44156 6132
rect 44212 6076 46000 6132
rect 31892 6020 31948 6076
rect 45200 6048 46000 6076
rect 14354 5964 14364 6020
rect 14420 5964 17724 6020
rect 17780 5964 20188 6020
rect 20244 5964 20860 6020
rect 20916 5964 20926 6020
rect 22418 5964 22428 6020
rect 22484 5964 25228 6020
rect 25284 5964 25294 6020
rect 31602 5964 31612 6020
rect 31668 5964 31948 6020
rect 42914 5964 42924 6020
rect 42980 5964 43932 6020
rect 43988 5964 43998 6020
rect 24322 5852 24332 5908
rect 24388 5852 28028 5908
rect 28084 5852 29484 5908
rect 29540 5852 29550 5908
rect 38658 5852 38668 5908
rect 38724 5852 40908 5908
rect 40964 5852 41468 5908
rect 41524 5852 41534 5908
rect 37090 5740 37100 5796
rect 37156 5740 37996 5796
rect 38052 5740 38062 5796
rect 12450 5628 12460 5684
rect 12516 5628 13356 5684
rect 13412 5628 15148 5684
rect 15204 5628 15214 5684
rect 33058 5628 33068 5684
rect 33124 5628 34748 5684
rect 34804 5628 41692 5684
rect 41748 5628 41758 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 12562 5180 12572 5236
rect 12628 5180 14252 5236
rect 14308 5180 14318 5236
rect 14914 5180 14924 5236
rect 14980 5180 15708 5236
rect 15764 5180 21644 5236
rect 21700 5180 21710 5236
rect 26852 5180 30604 5236
rect 30660 5180 30670 5236
rect 31892 5180 38668 5236
rect 38724 5180 38734 5236
rect 14252 5124 14308 5180
rect 26852 5124 26908 5180
rect 31892 5124 31948 5180
rect 14252 5068 16380 5124
rect 16436 5068 16446 5124
rect 16706 5068 16716 5124
rect 16772 5068 17388 5124
rect 17444 5068 17454 5124
rect 22194 5068 22204 5124
rect 22260 5068 24444 5124
rect 24500 5068 26908 5124
rect 30034 5068 30044 5124
rect 30100 5068 31052 5124
rect 31108 5068 31948 5124
rect 35970 5068 35980 5124
rect 36036 5068 41580 5124
rect 41636 5068 41646 5124
rect 17938 4956 17948 5012
rect 18004 4956 18844 5012
rect 18900 4956 18910 5012
rect 20290 4844 20300 4900
rect 20356 4844 21084 4900
rect 21140 4844 21150 4900
rect 23202 4844 23212 4900
rect 23268 4844 25228 4900
rect 25284 4844 25294 4900
rect 33618 4844 33628 4900
rect 33684 4844 42476 4900
rect 42532 4844 42542 4900
rect 16370 4732 16380 4788
rect 16436 4732 17388 4788
rect 17444 4732 17454 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 19282 4396 19292 4452
rect 19348 4396 19852 4452
rect 19908 4396 24332 4452
rect 24388 4396 24398 4452
rect 21634 4284 21644 4340
rect 21700 4284 22316 4340
rect 22372 4284 22382 4340
rect 24658 4284 24668 4340
rect 24724 4284 25452 4340
rect 25508 4284 25518 4340
rect 21410 4172 21420 4228
rect 21476 4172 22988 4228
rect 23044 4172 28140 4228
rect 28196 4172 28206 4228
rect 28578 4172 28588 4228
rect 28644 4172 29484 4228
rect 29540 4172 29932 4228
rect 29988 4172 30492 4228
rect 30548 4172 39116 4228
rect 39172 4172 41020 4228
rect 41076 4172 41086 4228
rect 19506 4060 19516 4116
rect 19572 4060 23772 4116
rect 23828 4060 23838 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 35186 3612 35196 3668
rect 35252 3612 37772 3668
rect 37828 3612 37838 3668
rect 12674 3500 12684 3556
rect 12740 3500 14028 3556
rect 14084 3500 19516 3556
rect 19572 3500 19582 3556
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 45200 2772 46000 2800
rect 44146 2716 44156 2772
rect 44212 2716 46000 2772
rect 45200 2688 46000 2716
<< via3 >>
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 36316 42028 36372 42084
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 35868 40908 35924 40964
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 35868 40236 35924 40292
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 36316 39004 36372 39060
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 29148 27804 29204 27860
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 35644 23660 35700 23716
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 35644 23324 35700 23380
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 34524 22428 34580 22484
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 19068 21868 19124 21924
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 34524 20748 34580 20804
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 29372 20300 29428 20356
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19068 15708 19124 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 29372 15260 29428 15316
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 29148 14476 29204 14532
rect 18844 14252 18900 14308
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 19628 13580 19684 13636
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19516 9884 19572 9940
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19628 8428 19684 8484
rect 22876 8428 22932 8484
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 22876 7532 22932 7588
rect 19516 7308 19572 7364
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 18844 6076 18900 6132
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 41580 4768 42396
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 42364 20128 42396
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 35168 41580 35488 42396
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 36316 42084 36372 42094
rect 35868 40964 35924 40974
rect 35868 40292 35924 40908
rect 35868 40226 35924 40236
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 36316 39060 36372 42028
rect 36316 38994 36372 39004
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 19068 21924 19124 21934
rect 19068 15764 19124 21868
rect 19068 15698 19124 15708
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 18844 14308 18900 14318
rect 18844 6132 18900 14252
rect 19808 14140 20128 15652
rect 29148 27860 29204 27870
rect 29148 14532 29204 27804
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35644 23716 35700 23726
rect 35644 23380 35700 23660
rect 35644 23314 35700 23324
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 34524 22484 34580 22494
rect 34524 20804 34580 22428
rect 34524 20738 34580 20748
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 29372 20356 29428 20366
rect 29372 15316 29428 20300
rect 29372 15250 29428 15260
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 29148 14466 29204 14476
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19628 13636 19684 13646
rect 19516 9940 19572 9950
rect 19516 7364 19572 9884
rect 19628 8484 19684 13580
rect 19628 8418 19684 8428
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19516 7298 19572 7308
rect 19808 7868 20128 9380
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 18844 6066 18900 6076
rect 19808 6300 20128 7812
rect 22876 8484 22932 8494
rect 22876 7588 22932 8428
rect 22876 7522 22932 7532
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0537_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0538_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28336 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0539_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23184 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0540_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27328 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0541_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22512 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0542_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27440 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0543_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25648 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0544_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27216 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0545_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0546_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0547_
timestamp 1698431365
transform -1 0 33600 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0548_
timestamp 1698431365
transform -1 0 30128 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0549_
timestamp 1698431365
transform -1 0 27664 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0550_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0551_
timestamp 1698431365
transform -1 0 24752 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0552_
timestamp 1698431365
transform -1 0 28112 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0553_
timestamp 1698431365
transform 1 0 18368 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0554_
timestamp 1698431365
transform 1 0 26320 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0555_
timestamp 1698431365
transform 1 0 24192 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0556_
timestamp 1698431365
transform -1 0 32144 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0557_
timestamp 1698431365
transform -1 0 30576 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0558_
timestamp 1698431365
transform 1 0 25648 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0559_
timestamp 1698431365
transform -1 0 25760 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0560_
timestamp 1698431365
transform -1 0 24640 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0561_
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0562_
timestamp 1698431365
transform 1 0 25536 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0563_
timestamp 1698431365
transform 1 0 28336 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0564_
timestamp 1698431365
transform -1 0 28112 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0565_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25648 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0566_
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0567_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27888 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0568_
timestamp 1698431365
transform 1 0 28336 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0569_
timestamp 1698431365
transform -1 0 17696 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0570_
timestamp 1698431365
transform 1 0 15568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0571_
timestamp 1698431365
transform 1 0 17808 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0572_
timestamp 1698431365
transform -1 0 24304 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0573_
timestamp 1698431365
transform -1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0574_
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0575_
timestamp 1698431365
transform -1 0 15344 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0576_
timestamp 1698431365
transform 1 0 13776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0577_
timestamp 1698431365
transform 1 0 15568 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0578_
timestamp 1698431365
transform 1 0 24976 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0579_
timestamp 1698431365
transform -1 0 20048 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0580_
timestamp 1698431365
transform 1 0 25424 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0581_
timestamp 1698431365
transform -1 0 22512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0582_
timestamp 1698431365
transform -1 0 22960 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0583_
timestamp 1698431365
transform 1 0 17584 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0584_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16800 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0585_
timestamp 1698431365
transform -1 0 12880 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0586_
timestamp 1698431365
transform -1 0 11088 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0587_
timestamp 1698431365
transform -1 0 15456 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0588_
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0589_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0590_
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0591_
timestamp 1698431365
transform -1 0 20720 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0592_
timestamp 1698431365
transform -1 0 21616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0593_
timestamp 1698431365
transform -1 0 28224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0594_
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0595_
timestamp 1698431365
transform -1 0 23744 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0596_
timestamp 1698431365
transform 1 0 9520 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0597_
timestamp 1698431365
transform -1 0 12208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0598_
timestamp 1698431365
transform 1 0 10752 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0599_
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0600_
timestamp 1698431365
transform 1 0 6944 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0601_
timestamp 1698431365
transform 1 0 9520 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0602_
timestamp 1698431365
transform 1 0 3024 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0603_
timestamp 1698431365
transform -1 0 4592 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0604_
timestamp 1698431365
transform 1 0 7504 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0605_
timestamp 1698431365
transform -1 0 10752 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0606_
timestamp 1698431365
transform 1 0 11536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0607_
timestamp 1698431365
transform 1 0 29008 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0608_
timestamp 1698431365
transform -1 0 41888 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0609_
timestamp 1698431365
transform -1 0 37296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0610_
timestamp 1698431365
transform 1 0 37296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0611_
timestamp 1698431365
transform -1 0 35392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0612_
timestamp 1698431365
transform -1 0 37744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0613_
timestamp 1698431365
transform -1 0 39088 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0614_
timestamp 1698431365
transform 1 0 37968 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0615_
timestamp 1698431365
transform -1 0 42000 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0616_
timestamp 1698431365
transform -1 0 41216 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0617_
timestamp 1698431365
transform -1 0 39648 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0618_
timestamp 1698431365
transform -1 0 41216 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0619_
timestamp 1698431365
transform 1 0 30688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0620_
timestamp 1698431365
transform -1 0 37744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0621_
timestamp 1698431365
transform -1 0 40320 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0622_
timestamp 1698431365
transform -1 0 41440 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0623_
timestamp 1698431365
transform 1 0 40096 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0624_
timestamp 1698431365
transform -1 0 37296 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0625_
timestamp 1698431365
transform -1 0 38864 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0626_
timestamp 1698431365
transform 1 0 37632 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0627_
timestamp 1698431365
transform -1 0 41664 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0628_
timestamp 1698431365
transform 1 0 33936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0629_
timestamp 1698431365
transform -1 0 36288 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0630_
timestamp 1698431365
transform -1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0631_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11088 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0632_
timestamp 1698431365
transform -1 0 9184 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0633_
timestamp 1698431365
transform -1 0 10752 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0634_
timestamp 1698431365
transform 1 0 7728 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0635_
timestamp 1698431365
transform -1 0 10752 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0636_
timestamp 1698431365
transform -1 0 8848 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0637_
timestamp 1698431365
transform 1 0 17248 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0638_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _0639_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15680 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0640_
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0641_
timestamp 1698431365
transform -1 0 22176 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0642_
timestamp 1698431365
transform -1 0 24528 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0643_
timestamp 1698431365
transform -1 0 19040 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0644_
timestamp 1698431365
transform 1 0 19600 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0645_
timestamp 1698431365
transform -1 0 20272 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0646_
timestamp 1698431365
transform -1 0 19264 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0647_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19712 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0648_
timestamp 1698431365
transform 1 0 11536 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0649_
timestamp 1698431365
transform -1 0 23408 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0650_
timestamp 1698431365
transform -1 0 24752 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0651_
timestamp 1698431365
transform -1 0 23184 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0652_
timestamp 1698431365
transform 1 0 11088 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0653_
timestamp 1698431365
transform -1 0 16128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0654_
timestamp 1698431365
transform -1 0 14560 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0655_
timestamp 1698431365
transform 1 0 12544 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0656_
timestamp 1698431365
transform -1 0 13664 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0657_
timestamp 1698431365
transform 1 0 13888 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0658_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19264 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0659_
timestamp 1698431365
transform 1 0 18928 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0660_
timestamp 1698431365
transform -1 0 14112 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0661_
timestamp 1698431365
transform 1 0 12096 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0662_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12320 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0663_
timestamp 1698431365
transform 1 0 15232 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0664_
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0665_
timestamp 1698431365
transform 1 0 15680 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0666_
timestamp 1698431365
transform 1 0 15120 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0667_
timestamp 1698431365
transform 1 0 13888 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0668_
timestamp 1698431365
transform 1 0 11760 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0669_
timestamp 1698431365
transform 1 0 14112 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0670_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11760 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0671_
timestamp 1698431365
transform -1 0 11424 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0672_
timestamp 1698431365
transform -1 0 9744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0673_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9744 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0674_
timestamp 1698431365
transform 1 0 11200 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0675_
timestamp 1698431365
transform -1 0 11312 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0676_
timestamp 1698431365
transform 1 0 13552 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0677_
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0678_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0679_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0680_
timestamp 1698431365
transform 1 0 19152 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0681_
timestamp 1698431365
transform 1 0 35616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0682_
timestamp 1698431365
transform -1 0 34720 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _0683_
timestamp 1698431365
transform -1 0 38080 0 -1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0684_
timestamp 1698431365
transform -1 0 39536 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0685_
timestamp 1698431365
transform 1 0 37968 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0686_
timestamp 1698431365
transform -1 0 39200 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0687_
timestamp 1698431365
transform 1 0 37744 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0688_
timestamp 1698431365
transform -1 0 36624 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0689_
timestamp 1698431365
transform -1 0 32032 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0690_
timestamp 1698431365
transform -1 0 35728 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0691_
timestamp 1698431365
transform -1 0 34496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0692_
timestamp 1698431365
transform 1 0 33824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0693_
timestamp 1698431365
transform 1 0 34608 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0694_
timestamp 1698431365
transform 1 0 34272 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0695_
timestamp 1698431365
transform 1 0 35056 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0696_
timestamp 1698431365
transform 1 0 34384 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0697_
timestamp 1698431365
transform -1 0 37296 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0698_
timestamp 1698431365
transform 1 0 36176 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0699_
timestamp 1698431365
transform -1 0 37968 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0700_
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0701_
timestamp 1698431365
transform 1 0 35728 0 -1 10976
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0702_
timestamp 1698431365
transform -1 0 31136 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0703_
timestamp 1698431365
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0704_
timestamp 1698431365
transform 1 0 34832 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0705_
timestamp 1698431365
transform -1 0 36176 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0706_
timestamp 1698431365
transform 1 0 33488 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0707_
timestamp 1698431365
transform -1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0708_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0709_
timestamp 1698431365
transform -1 0 37184 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0710_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0711_
timestamp 1698431365
transform -1 0 31360 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0712_
timestamp 1698431365
transform -1 0 37856 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0713_
timestamp 1698431365
transform 1 0 33152 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0714_
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0715_
timestamp 1698431365
transform -1 0 34608 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0716_
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0717_
timestamp 1698431365
transform 1 0 33600 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0718_
timestamp 1698431365
transform 1 0 34608 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0719_
timestamp 1698431365
transform -1 0 36848 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0720_
timestamp 1698431365
transform -1 0 37296 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0721_
timestamp 1698431365
transform 1 0 34832 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0722_
timestamp 1698431365
transform 1 0 34832 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0723_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35840 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0724_
timestamp 1698431365
transform -1 0 32144 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0725_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0726_
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0727_
timestamp 1698431365
transform -1 0 39424 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0728_
timestamp 1698431365
transform -1 0 38976 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0729_
timestamp 1698431365
transform -1 0 43008 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0730_
timestamp 1698431365
transform -1 0 42336 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0731_
timestamp 1698431365
transform -1 0 40096 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0732_
timestamp 1698431365
transform 1 0 39200 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0733_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0734_
timestamp 1698431365
transform -1 0 38192 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0735_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0736_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0737_
timestamp 1698431365
transform 1 0 39872 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0738_
timestamp 1698431365
transform 1 0 39424 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0739_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0740_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43904 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0741_
timestamp 1698431365
transform -1 0 41440 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0742_
timestamp 1698431365
transform -1 0 42560 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0743_
timestamp 1698431365
transform 1 0 42560 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0744_
timestamp 1698431365
transform 1 0 40096 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0745_
timestamp 1698431365
transform -1 0 40992 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0746_
timestamp 1698431365
transform -1 0 40544 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0747_
timestamp 1698431365
transform 1 0 39424 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0748_
timestamp 1698431365
transform 1 0 41104 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0749_
timestamp 1698431365
transform 1 0 43456 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0750_
timestamp 1698431365
transform -1 0 41104 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0751_
timestamp 1698431365
transform 1 0 38864 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0752_
timestamp 1698431365
transform 1 0 43456 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0753_
timestamp 1698431365
transform 1 0 39984 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0754_
timestamp 1698431365
transform 1 0 42896 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0755_
timestamp 1698431365
transform 1 0 42336 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0756_
timestamp 1698431365
transform 1 0 40880 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0757_
timestamp 1698431365
transform 1 0 43008 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0758_
timestamp 1698431365
transform -1 0 39760 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0759_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38976 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0760_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40208 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0761_
timestamp 1698431365
transform -1 0 39872 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0762_
timestamp 1698431365
transform -1 0 38864 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0763_
timestamp 1698431365
transform -1 0 34496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0764_
timestamp 1698431365
transform 1 0 34608 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0765_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38640 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0766_
timestamp 1698431365
transform -1 0 38192 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0767_
timestamp 1698431365
transform 1 0 36512 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0768_
timestamp 1698431365
transform -1 0 39872 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0769_
timestamp 1698431365
transform 1 0 38640 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0770_
timestamp 1698431365
transform -1 0 30240 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0771_
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0772_
timestamp 1698431365
transform 1 0 20272 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0773_
timestamp 1698431365
transform -1 0 21392 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0774_
timestamp 1698431365
transform 1 0 18032 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0775_
timestamp 1698431365
transform 1 0 17360 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0776_
timestamp 1698431365
transform -1 0 18816 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0777_
timestamp 1698431365
transform -1 0 17808 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0778_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15456 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0779_
timestamp 1698431365
transform 1 0 30576 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0780_
timestamp 1698431365
transform -1 0 17136 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0781_
timestamp 1698431365
transform -1 0 15232 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0782_
timestamp 1698431365
transform -1 0 40208 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0783_
timestamp 1698431365
transform -1 0 38864 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0784_
timestamp 1698431365
transform -1 0 38976 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0785_
timestamp 1698431365
transform -1 0 38192 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0786_
timestamp 1698431365
transform -1 0 37520 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0787_
timestamp 1698431365
transform 1 0 37744 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0788_
timestamp 1698431365
transform 1 0 37968 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0789_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25200 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0790_
timestamp 1698431365
transform -1 0 26544 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0791_
timestamp 1698431365
transform 1 0 27776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0792_
timestamp 1698431365
transform 1 0 30576 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _0793_
timestamp 1698431365
transform 1 0 36624 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0794_
timestamp 1698431365
transform -1 0 31360 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0795_
timestamp 1698431365
transform 1 0 25088 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0796_
timestamp 1698431365
transform 1 0 24304 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0797_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26544 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0798_
timestamp 1698431365
transform -1 0 37520 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0799_
timestamp 1698431365
transform -1 0 36624 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0800_
timestamp 1698431365
transform 1 0 31808 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0801_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25312 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0802_
timestamp 1698431365
transform -1 0 24864 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0803_
timestamp 1698431365
transform -1 0 25200 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0804_
timestamp 1698431365
transform -1 0 24864 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0805_
timestamp 1698431365
transform 1 0 28560 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0806_
timestamp 1698431365
transform 1 0 26768 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0807_
timestamp 1698431365
transform 1 0 25872 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0808_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26656 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0809_
timestamp 1698431365
transform 1 0 29120 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0810_
timestamp 1698431365
transform -1 0 36400 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0811_
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0812_
timestamp 1698431365
transform -1 0 37968 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0813_
timestamp 1698431365
transform 1 0 26544 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0814_
timestamp 1698431365
transform -1 0 26656 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0815_
timestamp 1698431365
transform -1 0 29904 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0816_
timestamp 1698431365
transform -1 0 29232 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0817_
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0818_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37520 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0819_
timestamp 1698431365
transform 1 0 35392 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0820_
timestamp 1698431365
transform -1 0 35392 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0821_
timestamp 1698431365
transform 1 0 34944 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0822_
timestamp 1698431365
transform 1 0 29568 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0823_
timestamp 1698431365
transform 1 0 30128 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0824_
timestamp 1698431365
transform 1 0 33264 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0825_
timestamp 1698431365
transform -1 0 30128 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0826_
timestamp 1698431365
transform 1 0 29232 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0827_
timestamp 1698431365
transform 1 0 30688 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0828_
timestamp 1698431365
transform 1 0 35280 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0829_
timestamp 1698431365
transform 1 0 33152 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0830_
timestamp 1698431365
transform 1 0 30800 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0831_
timestamp 1698431365
transform -1 0 37520 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0832_
timestamp 1698431365
transform -1 0 32704 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0833_
timestamp 1698431365
transform 1 0 34944 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0834_
timestamp 1698431365
transform -1 0 33488 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0835_
timestamp 1698431365
transform -1 0 34944 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0836_
timestamp 1698431365
transform 1 0 33488 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0837_
timestamp 1698431365
transform -1 0 36400 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0838_
timestamp 1698431365
transform -1 0 35616 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0839_
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0840_
timestamp 1698431365
transform -1 0 36288 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0841_
timestamp 1698431365
transform -1 0 36624 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0842_
timestamp 1698431365
transform -1 0 34384 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0843_
timestamp 1698431365
transform -1 0 34608 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0844_
timestamp 1698431365
transform -1 0 34272 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0845_
timestamp 1698431365
transform 1 0 31136 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0846_
timestamp 1698431365
transform -1 0 32704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0847_
timestamp 1698431365
transform 1 0 32032 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0848_
timestamp 1698431365
transform -1 0 30352 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0849_
timestamp 1698431365
transform 1 0 29904 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0850_
timestamp 1698431365
transform -1 0 27216 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0851_
timestamp 1698431365
transform -1 0 28784 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0852_
timestamp 1698431365
transform 1 0 29904 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0853_
timestamp 1698431365
transform -1 0 27888 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0854_
timestamp 1698431365
transform 1 0 30240 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0855_
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0856_
timestamp 1698431365
transform 1 0 29456 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0857_
timestamp 1698431365
transform 1 0 29680 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0858_
timestamp 1698431365
transform 1 0 30128 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0859_
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0860_
timestamp 1698431365
transform -1 0 32704 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0861_
timestamp 1698431365
transform -1 0 35840 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0862_
timestamp 1698431365
transform 1 0 8288 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0863_
timestamp 1698431365
transform -1 0 18032 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0864_
timestamp 1698431365
transform -1 0 21840 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0865_
timestamp 1698431365
transform -1 0 16912 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0866_
timestamp 1698431365
transform -1 0 15120 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0867_
timestamp 1698431365
transform 1 0 15344 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0868_
timestamp 1698431365
transform -1 0 15232 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0869_
timestamp 1698431365
transform -1 0 16464 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0870_
timestamp 1698431365
transform 1 0 17808 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0871_
timestamp 1698431365
transform -1 0 18480 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0872_
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0873_
timestamp 1698431365
transform -1 0 16128 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0874_
timestamp 1698431365
transform 1 0 18480 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0875_
timestamp 1698431365
transform -1 0 20720 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0876_
timestamp 1698431365
transform -1 0 25872 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0877_
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0878_
timestamp 1698431365
transform -1 0 21952 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0879_
timestamp 1698431365
transform -1 0 31024 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0880_
timestamp 1698431365
transform 1 0 21952 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0881_
timestamp 1698431365
transform -1 0 21952 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0882_
timestamp 1698431365
transform -1 0 22400 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0883_
timestamp 1698431365
transform -1 0 30464 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0884_
timestamp 1698431365
transform 1 0 21504 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0885_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0886_
timestamp 1698431365
transform -1 0 32256 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0887_
timestamp 1698431365
transform 1 0 22624 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0888_
timestamp 1698431365
transform -1 0 23408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0889_
timestamp 1698431365
transform 1 0 31024 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0890_
timestamp 1698431365
transform 1 0 21952 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0891_
timestamp 1698431365
transform 1 0 23408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0892_
timestamp 1698431365
transform -1 0 19824 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0893_
timestamp 1698431365
transform -1 0 21280 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0894_
timestamp 1698431365
transform -1 0 13328 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0895_
timestamp 1698431365
transform -1 0 12544 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0896_
timestamp 1698431365
transform 1 0 10864 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0897_
timestamp 1698431365
transform 1 0 19264 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0898_
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0899_
timestamp 1698431365
transform 1 0 11760 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0900_
timestamp 1698431365
transform 1 0 15344 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0901_
timestamp 1698431365
transform 1 0 14112 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0902_
timestamp 1698431365
transform -1 0 15568 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0903_
timestamp 1698431365
transform 1 0 13664 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0904_
timestamp 1698431365
transform -1 0 28672 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0905_
timestamp 1698431365
transform -1 0 26880 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0906_
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0907_
timestamp 1698431365
transform 1 0 22624 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0908_
timestamp 1698431365
transform -1 0 21616 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0909_
timestamp 1698431365
transform -1 0 22736 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0910_
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0911_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0912_
timestamp 1698431365
transform -1 0 20272 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0913_
timestamp 1698431365
transform -1 0 22064 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0914_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0915_
timestamp 1698431365
transform -1 0 25760 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0916_
timestamp 1698431365
transform -1 0 31808 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0917_
timestamp 1698431365
transform -1 0 31136 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0918_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25200 0 1 15680
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0919_
timestamp 1698431365
transform -1 0 24192 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0920_
timestamp 1698431365
transform -1 0 19264 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0921_
timestamp 1698431365
transform -1 0 19376 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0922_
timestamp 1698431365
transform 1 0 18704 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0923_
timestamp 1698431365
transform -1 0 28336 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0924_
timestamp 1698431365
transform 1 0 27776 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0925_
timestamp 1698431365
transform -1 0 29008 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0926_
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0927_
timestamp 1698431365
transform -1 0 27440 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0928_
timestamp 1698431365
transform -1 0 22400 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0929_
timestamp 1698431365
transform 1 0 21952 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0930_
timestamp 1698431365
transform -1 0 23408 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0931_
timestamp 1698431365
transform -1 0 21952 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0932_
timestamp 1698431365
transform -1 0 21616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0933_
timestamp 1698431365
transform -1 0 18144 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0934_
timestamp 1698431365
transform 1 0 15344 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0935_
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0936_
timestamp 1698431365
transform -1 0 15344 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0937_
timestamp 1698431365
transform -1 0 14336 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0938_
timestamp 1698431365
transform -1 0 24752 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0939_
timestamp 1698431365
transform -1 0 13104 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0940_
timestamp 1698431365
transform -1 0 12768 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0941_
timestamp 1698431365
transform 1 0 13664 0 1 3136
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0942_
timestamp 1698431365
transform 1 0 14336 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0943_
timestamp 1698431365
transform -1 0 20384 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0944_
timestamp 1698431365
transform -1 0 18704 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0945_
timestamp 1698431365
transform 1 0 23408 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0946_
timestamp 1698431365
transform -1 0 25760 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0947_
timestamp 1698431365
transform 1 0 30464 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0948_
timestamp 1698431365
transform -1 0 30464 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0949_
timestamp 1698431365
transform -1 0 29680 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0950_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0951_
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0952_
timestamp 1698431365
transform -1 0 29904 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0953_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0954_
timestamp 1698431365
transform -1 0 22736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0955_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19712 0 -1 23520
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0956_
timestamp 1698431365
transform -1 0 6720 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0957_
timestamp 1698431365
transform 1 0 7952 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0958_
timestamp 1698431365
transform 1 0 10416 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0959_
timestamp 1698431365
transform -1 0 12768 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0960_
timestamp 1698431365
transform 1 0 9408 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0961_
timestamp 1698431365
transform -1 0 14448 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0962_
timestamp 1698431365
transform 1 0 10752 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0963_
timestamp 1698431365
transform 1 0 12320 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0964_
timestamp 1698431365
transform -1 0 7952 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0965_
timestamp 1698431365
transform 1 0 8064 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0966_
timestamp 1698431365
transform -1 0 11200 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0967_
timestamp 1698431365
transform -1 0 6720 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0968_
timestamp 1698431365
transform 1 0 6048 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0969_
timestamp 1698431365
transform -1 0 8848 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0970_
timestamp 1698431365
transform 1 0 6272 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0971_
timestamp 1698431365
transform -1 0 8176 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0972_
timestamp 1698431365
transform 1 0 3920 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0973_
timestamp 1698431365
transform -1 0 6160 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0974_
timestamp 1698431365
transform -1 0 8064 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0975_
timestamp 1698431365
transform -1 0 6832 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0976_
timestamp 1698431365
transform -1 0 5264 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0977_
timestamp 1698431365
transform -1 0 6720 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0978_
timestamp 1698431365
transform 1 0 4592 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0979_
timestamp 1698431365
transform 1 0 6720 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0980_
timestamp 1698431365
transform 1 0 8176 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0981_
timestamp 1698431365
transform 1 0 6720 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0982_
timestamp 1698431365
transform 1 0 9408 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0983_
timestamp 1698431365
transform 1 0 26992 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0984_
timestamp 1698431365
transform -1 0 27440 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0985_
timestamp 1698431365
transform 1 0 25760 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0986_
timestamp 1698431365
transform 1 0 25088 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0987_
timestamp 1698431365
transform 1 0 27440 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0988_
timestamp 1698431365
transform 1 0 28112 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0989_
timestamp 1698431365
transform -1 0 30016 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0990_
timestamp 1698431365
transform 1 0 29120 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0991_
timestamp 1698431365
transform 1 0 30016 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0992_
timestamp 1698431365
transform -1 0 14000 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0993_
timestamp 1698431365
transform 1 0 12096 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0994_
timestamp 1698431365
transform -1 0 13552 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0995_
timestamp 1698431365
transform -1 0 13888 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0996_
timestamp 1698431365
transform -1 0 9184 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0997_
timestamp 1698431365
transform 1 0 15344 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0998_
timestamp 1698431365
transform -1 0 15680 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0999_
timestamp 1698431365
transform -1 0 13104 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1000_
timestamp 1698431365
transform -1 0 13664 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1001_
timestamp 1698431365
transform 1 0 21616 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1002_
timestamp 1698431365
transform 1 0 21280 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1003_
timestamp 1698431365
transform 1 0 19152 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1004_
timestamp 1698431365
transform -1 0 20272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1005_
timestamp 1698431365
transform 1 0 18480 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1006_
timestamp 1698431365
transform -1 0 17024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1007_
timestamp 1698431365
transform -1 0 19488 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1008_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1009_
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1010_
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1011_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28112 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1012_
timestamp 1698431365
transform 1 0 30240 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1013_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30800 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1014_
timestamp 1698431365
transform -1 0 41552 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1015_
timestamp 1698431365
transform -1 0 41664 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1016_
timestamp 1698431365
transform 1 0 40880 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1017_
timestamp 1698431365
transform -1 0 43008 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1018_
timestamp 1698431365
transform -1 0 39760 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1019_
timestamp 1698431365
transform -1 0 38752 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1020_
timestamp 1698431365
transform 1 0 38192 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1021_
timestamp 1698431365
transform 1 0 39312 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1022_
timestamp 1698431365
transform -1 0 39312 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1023_
timestamp 1698431365
transform -1 0 38080 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1024_
timestamp 1698431365
transform 1 0 39424 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1025_
timestamp 1698431365
transform 1 0 40544 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1026_
timestamp 1698431365
transform 1 0 42560 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1027_
timestamp 1698431365
transform -1 0 42560 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1028_
timestamp 1698431365
transform -1 0 40544 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1029_
timestamp 1698431365
transform -1 0 42896 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1030_
timestamp 1698431365
transform -1 0 41664 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1031_
timestamp 1698431365
transform 1 0 41776 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1032_
timestamp 1698431365
transform -1 0 43792 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1033_
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1034_
timestamp 1698431365
transform 1 0 42448 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1035_
timestamp 1698431365
transform -1 0 43792 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1036_
timestamp 1698431365
transform -1 0 43904 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1037_
timestamp 1698431365
transform -1 0 43008 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1038_
timestamp 1698431365
transform 1 0 41440 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1039_
timestamp 1698431365
transform -1 0 43568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1040_
timestamp 1698431365
transform 1 0 41664 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1041_
timestamp 1698431365
transform -1 0 44128 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1042_
timestamp 1698431365
transform -1 0 20272 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1043_
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1044_
timestamp 1698431365
transform -1 0 16912 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1045_
timestamp 1698431365
transform -1 0 19600 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1046_
timestamp 1698431365
transform 1 0 18032 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1047_
timestamp 1698431365
transform 1 0 14560 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1048_
timestamp 1698431365
transform -1 0 12992 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1049_
timestamp 1698431365
transform 1 0 27328 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1050_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1051_
timestamp 1698431365
transform 1 0 34272 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1052_
timestamp 1698431365
transform 1 0 34048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1053_
timestamp 1698431365
transform -1 0 32704 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1054_
timestamp 1698431365
transform -1 0 32816 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1055_
timestamp 1698431365
transform 1 0 34944 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1056_
timestamp 1698431365
transform 1 0 32480 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1057_
timestamp 1698431365
transform 1 0 31696 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1058_
timestamp 1698431365
transform -1 0 32704 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1059_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30352 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1060_
timestamp 1698431365
transform 1 0 28336 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1061_
timestamp 1698431365
transform 1 0 27664 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1062_
timestamp 1698431365
transform 1 0 31696 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1063_
timestamp 1698431365
transform 1 0 32144 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1064_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1065_
timestamp 1698431365
transform 1 0 30016 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1066_
timestamp 1698431365
transform -1 0 30128 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1067_
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1068_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1069_
timestamp 1698431365
transform -1 0 24304 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1070_
timestamp 1698431365
transform 1 0 28336 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1071_
timestamp 1698431365
transform -1 0 39200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1072_
timestamp 1698431365
transform 1 0 39648 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1073_
timestamp 1698431365
transform 1 0 38976 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1074_
timestamp 1698431365
transform -1 0 41440 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1075_
timestamp 1698431365
transform -1 0 42896 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1076_
timestamp 1698431365
transform -1 0 42448 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1077_
timestamp 1698431365
transform -1 0 43120 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1078_
timestamp 1698431365
transform -1 0 43680 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1079_
timestamp 1698431365
transform 1 0 42448 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1080_
timestamp 1698431365
transform 1 0 41440 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1081_
timestamp 1698431365
transform 1 0 42896 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1082_
timestamp 1698431365
transform 1 0 39648 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1083_
timestamp 1698431365
transform -1 0 42224 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1084_
timestamp 1698431365
transform -1 0 40544 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1085_
timestamp 1698431365
transform 1 0 41104 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1086_
timestamp 1698431365
transform -1 0 43792 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1087_
timestamp 1698431365
transform -1 0 43568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1088_
timestamp 1698431365
transform 1 0 41104 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1089_
timestamp 1698431365
transform -1 0 42448 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1090_
timestamp 1698431365
transform 1 0 41216 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1091_
timestamp 1698431365
transform 1 0 42560 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1092_
timestamp 1698431365
transform -1 0 39872 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1093_
timestamp 1698431365
transform -1 0 38752 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1094_
timestamp 1698431365
transform -1 0 39984 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1095_
timestamp 1698431365
transform -1 0 39424 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1096_
timestamp 1698431365
transform -1 0 38304 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1097_
timestamp 1698431365
transform -1 0 37744 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1098_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28672 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1099_
timestamp 1698431365
transform 1 0 27104 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1100_
timestamp 1698431365
transform 1 0 26432 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1101_
timestamp 1698431365
transform 1 0 29680 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1102_
timestamp 1698431365
transform 1 0 30128 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1103_
timestamp 1698431365
transform 1 0 30688 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1104_
timestamp 1698431365
transform 1 0 30352 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1105_
timestamp 1698431365
transform 1 0 30688 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1106_
timestamp 1698431365
transform 1 0 28112 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1107_
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1108_
timestamp 1698431365
transform 1 0 33824 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1109_
timestamp 1698431365
transform 1 0 34832 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1110_
timestamp 1698431365
transform 1 0 31248 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1111_
timestamp 1698431365
transform -1 0 31472 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1112_
timestamp 1698431365
transform 1 0 32368 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1113_
timestamp 1698431365
transform -1 0 34720 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1114_
timestamp 1698431365
transform 1 0 32032 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1115_
timestamp 1698431365
transform -1 0 34832 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1116_
timestamp 1698431365
transform -1 0 28448 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1117_
timestamp 1698431365
transform 1 0 25872 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1118_
timestamp 1698431365
transform -1 0 25760 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1119_
timestamp 1698431365
transform 1 0 28112 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1120_
timestamp 1698431365
transform 1 0 29344 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1121_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1122_
timestamp 1698431365
transform 1 0 26096 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1123_
timestamp 1698431365
transform 1 0 25312 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1124_
timestamp 1698431365
transform 1 0 29904 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1125_
timestamp 1698431365
transform 1 0 30576 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1126_
timestamp 1698431365
transform -1 0 27216 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1127_
timestamp 1698431365
transform -1 0 27776 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1128_
timestamp 1698431365
transform 1 0 25760 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1129_
timestamp 1698431365
transform -1 0 28560 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1130_
timestamp 1698431365
transform -1 0 29008 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1131_
timestamp 1698431365
transform -1 0 28336 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1132_
timestamp 1698431365
transform -1 0 20832 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1133_
timestamp 1698431365
transform -1 0 20048 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1134_
timestamp 1698431365
transform -1 0 21616 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1135_
timestamp 1698431365
transform 1 0 22288 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1136_
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1137_
timestamp 1698431365
transform -1 0 18032 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1138_
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1139_
timestamp 1698431365
transform 1 0 16128 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1140_
timestamp 1698431365
transform -1 0 17696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1141_
timestamp 1698431365
transform 1 0 18032 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1142_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44016 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1143_
timestamp 1698431365
transform 1 0 35616 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1144_
timestamp 1698431365
transform -1 0 42448 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1145_
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1146_
timestamp 1698431365
transform -1 0 44016 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1147_
timestamp 1698431365
transform 1 0 40992 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1148_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1149_
timestamp 1698431365
transform 1 0 41104 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1150_
timestamp 1698431365
transform -1 0 44240 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1151_
timestamp 1698431365
transform -1 0 44240 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1152_
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1153_
timestamp 1698431365
transform 1 0 40992 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1154_
timestamp 1698431365
transform 1 0 17248 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1155_
timestamp 1698431365
transform -1 0 17248 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1156_
timestamp 1698431365
transform -1 0 16576 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1157_
timestamp 1698431365
transform 1 0 37408 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1158_
timestamp 1698431365
transform 1 0 37856 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1159_
timestamp 1698431365
transform 1 0 31808 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1160_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1161_
timestamp 1698431365
transform 1 0 31360 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1162_
timestamp 1698431365
transform 1 0 34496 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1163_
timestamp 1698431365
transform 1 0 32592 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1164_
timestamp 1698431365
transform 1 0 31472 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1165_
timestamp 1698431365
transform 1 0 32256 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1166_
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1167_
timestamp 1698431365
transform -1 0 37520 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1168_
timestamp 1698431365
transform 1 0 31584 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1169_
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1170_
timestamp 1698431365
transform 1 0 26656 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1171_
timestamp 1698431365
transform 1 0 26992 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1172_
timestamp 1698431365
transform -1 0 34048 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1173_
timestamp 1698431365
transform -1 0 10416 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1174_
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1175_
timestamp 1698431365
transform 1 0 20048 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1176_
timestamp 1698431365
transform 1 0 21056 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1177_
timestamp 1698431365
transform 1 0 19936 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1178_
timestamp 1698431365
transform 1 0 8400 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1179_
timestamp 1698431365
transform 1 0 7504 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1180_
timestamp 1698431365
transform -1 0 9184 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1181_
timestamp 1698431365
transform 1 0 7056 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1182_
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1183_
timestamp 1698431365
transform 1 0 7392 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _1184_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1185_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10752 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _1186_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1187_
timestamp 1698431365
transform 1 0 10864 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _1188_
timestamp 1698431365
transform 1 0 12432 0 -1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1189_
timestamp 1698431365
transform 1 0 15344 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _1190_
timestamp 1698431365
transform -1 0 18480 0 1 32928
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _1191_
timestamp 1698431365
transform 1 0 16128 0 1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1192_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1193_
timestamp 1698431365
transform 1 0 19712 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1194_
timestamp 1698431365
transform -1 0 21504 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1195_
timestamp 1698431365
transform 1 0 22512 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1196_
timestamp 1698431365
transform 1 0 22624 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1197_
timestamp 1698431365
transform 1 0 9184 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1198_
timestamp 1698431365
transform -1 0 12656 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1199_
timestamp 1698431365
transform 1 0 13776 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1200_
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1201_
timestamp 1698431365
transform 1 0 22400 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1202_
timestamp 1698431365
transform 1 0 19824 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1203_
timestamp 1698431365
transform 1 0 19264 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1204_
timestamp 1698431365
transform 1 0 23744 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1205_
timestamp 1698431365
transform 1 0 17696 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1206_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1207_
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1208_
timestamp 1698431365
transform 1 0 20048 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1209_
timestamp 1698431365
transform 1 0 17136 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1210_
timestamp 1698431365
transform 1 0 13216 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1211_
timestamp 1698431365
transform 1 0 10528 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1212_
timestamp 1698431365
transform 1 0 8624 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1213_
timestamp 1698431365
transform 1 0 11872 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1214_
timestamp 1698431365
transform -1 0 20608 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1215_
timestamp 1698431365
transform -1 0 26208 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1216_
timestamp 1698431365
transform 1 0 24976 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1217_
timestamp 1698431365
transform -1 0 13104 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1218_
timestamp 1698431365
transform 1 0 9968 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1219_
timestamp 1698431365
transform 1 0 10640 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1220_
timestamp 1698431365
transform -1 0 12208 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1221_
timestamp 1698431365
transform -1 0 9072 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1222_
timestamp 1698431365
transform -1 0 9520 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1223_
timestamp 1698431365
transform -1 0 5376 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1224_
timestamp 1698431365
transform 1 0 1904 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1225_
timestamp 1698431365
transform 1 0 3696 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1226_
timestamp 1698431365
transform 1 0 6720 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1227_
timestamp 1698431365
transform -1 0 14112 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1228_
timestamp 1698431365
transform 1 0 19712 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1229_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25200 0 -1 36064
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1230_
timestamp 1698431365
transform -1 0 26768 0 1 36064
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1231_
timestamp 1698431365
transform 1 0 21728 0 1 34496
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1232_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1233_
timestamp 1698431365
transform 1 0 28336 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1234_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1235_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1236_
timestamp 1698431365
transform 1 0 8848 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1237_
timestamp 1698431365
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1238_
timestamp 1698431365
transform 1 0 9744 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1239_
timestamp 1698431365
transform 1 0 19712 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1240_
timestamp 1698431365
transform -1 0 18480 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1241_
timestamp 1698431365
transform -1 0 18368 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1242_
timestamp 1698431365
transform 1 0 19824 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1243_
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1244_
timestamp 1698431365
transform 1 0 34496 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1245_
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1246_
timestamp 1698431365
transform 1 0 34048 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1247_
timestamp 1698431365
transform 1 0 35952 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1248_
timestamp 1698431365
transform 1 0 37968 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1249_
timestamp 1698431365
transform 1 0 38640 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1250_
timestamp 1698431365
transform 1 0 40544 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1251_
timestamp 1698431365
transform 1 0 39648 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1252_
timestamp 1698431365
transform 1 0 38640 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1253_
timestamp 1698431365
transform 1 0 36736 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1254_
timestamp 1698431365
transform 1 0 29456 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1255_
timestamp 1698431365
transform 1 0 14784 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1256_
timestamp 1698431365
transform -1 0 19264 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1257_
timestamp 1698431365
transform 1 0 10752 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1258_
timestamp 1698431365
transform 1 0 33376 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1259_
timestamp 1698431365
transform 1 0 31024 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1260_
timestamp 1698431365
transform 1 0 32928 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1261_
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1262_
timestamp 1698431365
transform 1 0 27440 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1263_
timestamp 1698431365
transform 1 0 31808 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1264_
timestamp 1698431365
transform 1 0 28896 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1265_
timestamp 1698431365
transform 1 0 33152 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1266_
timestamp 1698431365
transform 1 0 36624 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1267_
timestamp 1698431365
transform 1 0 38640 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1268_
timestamp 1698431365
transform 1 0 40432 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1269_
timestamp 1698431365
transform 1 0 40544 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1270_
timestamp 1698431365
transform 1 0 35952 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1271_
timestamp 1698431365
transform 1 0 37968 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1272_
timestamp 1698431365
transform 1 0 38864 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1273_
timestamp 1698431365
transform 1 0 40544 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1274_
timestamp 1698431365
transform 1 0 34384 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1275_
timestamp 1698431365
transform 1 0 34832 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1276_
timestamp 1698431365
transform 1 0 32816 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1277_
timestamp 1698431365
transform -1 0 32704 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1278_
timestamp 1698431365
transform 1 0 26768 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1279_
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1280_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1281_
timestamp 1698431365
transform 1 0 33376 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1282_
timestamp 1698431365
transform 1 0 30016 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1283_
timestamp 1698431365
transform 1 0 33040 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1284_
timestamp 1698431365
transform 1 0 33264 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1285_
timestamp 1698431365
transform 1 0 23856 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1286_
timestamp 1698431365
transform 1 0 28784 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1287_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1288_
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1289_
timestamp 1698431365
transform 1 0 40992 0 -1 26656
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _1290_
timestamp 1698431365
transform 1 0 40992 0 1 26656
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1291_
timestamp 1698431365
transform 1 0 24080 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1292_
timestamp 1698431365
transform 1 0 24976 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1293_
timestamp 1698431365
transform 1 0 23184 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1294_
timestamp 1698431365
transform 1 0 23296 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1295_
timestamp 1698431365
transform 1 0 16016 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1296_
timestamp 1698431365
transform -1 0 19040 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _1297_
timestamp 1698431365
transform 1 0 18256 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1298_
timestamp 1698431365
transform 1 0 20608 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1299_
timestamp 1698431365
transform 1 0 18480 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1300_
timestamp 1698431365
transform 1 0 15680 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1301_
timestamp 1698431365
transform 1 0 13552 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1302_
timestamp 1698431365
transform -1 0 16800 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _1303_
timestamp 1698431365
transform 1 0 16016 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0537__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0540__A1
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0540__A2
timestamp 1698431365
transform 1 0 27664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0542__A1
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0542__A2
timestamp 1698431365
transform 1 0 27440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0545__I0
timestamp 1698431365
transform 1 0 29232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0550__I0
timestamp 1698431365
transform -1 0 27664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0553__I
timestamp 1698431365
transform -1 0 18368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0554__I0
timestamp 1698431365
transform 1 0 23968 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0556__I
timestamp 1698431365
transform 1 0 33040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0558__I0
timestamp 1698431365
transform 1 0 27552 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0577__I
timestamp 1698431365
transform 1 0 15344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0578__A2
timestamp 1698431365
transform -1 0 26432 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0579__I
timestamp 1698431365
transform 1 0 20272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0726__I
timestamp 1698431365
transform -1 0 38864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0763__I
timestamp 1698431365
transform -1 0 34048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__I1
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__A1
timestamp 1698431365
transform 1 0 17808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0780__A1
timestamp 1698431365
transform -1 0 17584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0845__A1
timestamp 1698431365
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__I
timestamp 1698431365
transform 1 0 34720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__I
timestamp 1698431365
transform 1 0 9184 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__I
timestamp 1698431365
transform 1 0 18256 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__I
timestamp 1698431365
transform 1 0 19376 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__I
timestamp 1698431365
transform -1 0 31248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__A1
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0884__A1
timestamp 1698431365
transform 1 0 22400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0887__A1
timestamp 1698431365
transform -1 0 23744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__I
timestamp 1698431365
transform -1 0 32144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__A1
timestamp 1698431365
transform 1 0 22848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0895__A1
timestamp 1698431365
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0897__I
timestamp 1698431365
transform 1 0 20160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0898__A1
timestamp 1698431365
transform 1 0 13552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0900__I1
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0902__A1
timestamp 1698431365
transform 1 0 15792 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__I
timestamp 1698431365
transform -1 0 29456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__A1
timestamp 1698431365
transform -1 0 27104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__I0
timestamp 1698431365
transform 1 0 24864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A1
timestamp 1698431365
transform 1 0 23408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__A1
timestamp 1698431365
transform -1 0 18928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0914__I0
timestamp 1698431365
transform 1 0 26880 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0916__I
timestamp 1698431365
transform -1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__A1
timestamp 1698431365
transform 1 0 19040 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__A2
timestamp 1698431365
transform 1 0 18144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A1
timestamp 1698431365
transform 1 0 29904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0926__A1
timestamp 1698431365
transform 1 0 29456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__A1
timestamp 1698431365
transform -1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__A2
timestamp 1698431365
transform -1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__B
timestamp 1698431365
transform -1 0 21840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0964__I
timestamp 1698431365
transform -1 0 7056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__I
timestamp 1698431365
transform 1 0 8288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__I0
timestamp 1698431365
transform 1 0 29568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A1
timestamp 1698431365
transform 1 0 27888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0990__A1
timestamp 1698431365
transform 1 0 30688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0992__I
timestamp 1698431365
transform -1 0 14224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0993__A1
timestamp 1698431365
transform 1 0 14224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__A1
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0997__I1
timestamp 1698431365
transform 1 0 17696 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0997__S
timestamp 1698431365
transform 1 0 17248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0999__I1
timestamp 1698431365
transform -1 0 14336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0999__S
timestamp 1698431365
transform -1 0 14672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1002__I0
timestamp 1698431365
transform 1 0 23184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1005__A1
timestamp 1698431365
transform -1 0 19376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__A1
timestamp 1698431365
transform -1 0 19824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__I0
timestamp 1698431365
transform 1 0 23072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1013__A1
timestamp 1698431365
transform -1 0 29456 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A1
timestamp 1698431365
transform 1 0 40992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1024__I
timestamp 1698431365
transform 1 0 39200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__I0
timestamp 1698431365
transform 1 0 19824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1045__A1
timestamp 1698431365
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__I0
timestamp 1698431365
transform 1 0 17136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__I0
timestamp 1698431365
transform 1 0 30800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A1
timestamp 1698431365
transform 1 0 31472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__I1
timestamp 1698431365
transform 1 0 30016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A1
timestamp 1698431365
transform -1 0 32256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__I1
timestamp 1698431365
transform 1 0 32480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__A1
timestamp 1698431365
transform 1 0 33712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A1
timestamp 1698431365
transform 1 0 28112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A1
timestamp 1698431365
transform 1 0 38752 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__A1
timestamp 1698431365
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__I1
timestamp 1698431365
transform 1 0 30240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__A1
timestamp 1698431365
transform 1 0 29232 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__A1
timestamp 1698431365
transform 1 0 31136 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1110__I0
timestamp 1698431365
transform 1 0 31696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__A1
timestamp 1698431365
transform 1 0 31808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__I0
timestamp 1698431365
transform 1 0 27776 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A1
timestamp 1698431365
transform -1 0 29792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__I0
timestamp 1698431365
transform 1 0 29120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1124__A1
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__I
timestamp 1698431365
transform 1 0 27888 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__CLK
timestamp 1698431365
transform 1 0 32368 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__CLK
timestamp 1698431365
transform 1 0 34272 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__CLK
timestamp 1698431365
transform 1 0 20944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__CLK
timestamp 1698431365
transform -1 0 13216 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1221__CLK
timestamp 1698431365
transform 1 0 9072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1247__CLK
timestamp 1698431365
transform 1 0 35728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__CLK
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1289__D
timestamp 1698431365
transform 1 0 44128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1290__CLKN
timestamp 1698431365
transform 1 0 40768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1290__D
timestamp 1698431365
transform -1 0 43232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1302__CLKN
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout24_I
timestamp 1698431365
transform 1 0 20272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout41_I
timestamp 1698431365
transform 1 0 37072 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout47_I
timestamp 1698431365
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout52_I
timestamp 1698431365
transform 1 0 32480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout61_I
timestamp 1698431365
transform 1 0 43792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 44352 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 43456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 44352 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 43680 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 44352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 44352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 43680 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 43680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout14
timestamp 1698431365
transform -1 0 28336 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout15
timestamp 1698431365
transform 1 0 19600 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout16
timestamp 1698431365
transform -1 0 10976 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout17
timestamp 1698431365
transform -1 0 7504 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout18
timestamp 1698431365
transform -1 0 11760 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout19
timestamp 1698431365
transform -1 0 11648 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout20
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout21
timestamp 1698431365
transform -1 0 16352 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout22
timestamp 1698431365
transform -1 0 19152 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout23
timestamp 1698431365
transform -1 0 19824 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout24
timestamp 1698431365
transform -1 0 19600 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout25
timestamp 1698431365
transform -1 0 20496 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout26
timestamp 1698431365
transform -1 0 10640 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout27
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout28
timestamp 1698431365
transform -1 0 15344 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout29
timestamp 1698431365
transform -1 0 19376 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout30
timestamp 1698431365
transform 1 0 18928 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout31
timestamp 1698431365
transform -1 0 20048 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout32
timestamp 1698431365
transform -1 0 20720 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout33
timestamp 1698431365
transform -1 0 20720 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout34
timestamp 1698431365
transform -1 0 22064 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout35
timestamp 1698431365
transform -1 0 21392 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout36
timestamp 1698431365
transform -1 0 24640 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout37
timestamp 1698431365
transform -1 0 29680 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout38
timestamp 1698431365
transform -1 0 32928 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout39
timestamp 1698431365
transform 1 0 32032 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout40
timestamp 1698431365
transform -1 0 33376 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout41
timestamp 1698431365
transform -1 0 36400 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout42
timestamp 1698431365
transform -1 0 24192 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout43
timestamp 1698431365
transform -1 0 24976 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout44
timestamp 1698431365
transform -1 0 26208 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout45
timestamp 1698431365
transform 1 0 32928 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout46
timestamp 1698431365
transform -1 0 33264 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout47
timestamp 1698431365
transform -1 0 33600 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout48
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout49
timestamp 1698431365
transform -1 0 30800 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout50
timestamp 1698431365
transform -1 0 32368 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout51
timestamp 1698431365
transform 1 0 31360 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout52
timestamp 1698431365
transform -1 0 33376 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout53
timestamp 1698431365
transform -1 0 32592 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout54
timestamp 1698431365
transform -1 0 40544 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout55
timestamp 1698431365
transform -1 0 43904 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout56
timestamp 1698431365
transform 1 0 38640 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout57
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout58
timestamp 1698431365
transform 1 0 39872 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout59
timestamp 1698431365
transform -1 0 40544 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout60
timestamp 1698431365
transform 1 0 39872 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout61
timestamp 1698431365
transform -1 0 42336 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_104 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_108 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_123 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15120 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_131
timestamp 1698431365
transform 1 0 16016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_181
timestamp 1698431365
transform 1 0 21616 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_189
timestamp 1698431365
transform 1 0 22512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_197
timestamp 1698431365
transform 1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_274 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_290
timestamp 1698431365
transform 1 0 33824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_298
timestamp 1698431365
transform 1 0 34720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_304
timestamp 1698431365
transform 1 0 35392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_316
timestamp 1698431365
transform 1 0 36736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_320
timestamp 1698431365
transform 1 0 37184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_334
timestamp 1698431365
transform 1 0 38752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_338
timestamp 1698431365
transform 1 0 39200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_88
timestamp 1698431365
transform 1 0 11200 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_92
timestamp 1698431365
transform 1 0 11648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_128
timestamp 1698431365
transform 1 0 15680 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_132
timestamp 1698431365
transform 1 0 16128 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_154
timestamp 1698431365
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698431365
transform 1 0 18816 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_170
timestamp 1698431365
transform 1 0 20384 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_218
timestamp 1698431365
transform 1 0 25760 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_234
timestamp 1698431365
transform 1 0 27552 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_249
timestamp 1698431365
transform 1 0 29232 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_253
timestamp 1698431365
transform 1 0 29680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_257
timestamp 1698431365
transform 1 0 30128 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_266
timestamp 1698431365
transform 1 0 31136 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_274
timestamp 1698431365
transform 1 0 32032 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698431365
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_290
timestamp 1698431365
transform 1 0 33824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_345
timestamp 1698431365
transform 1 0 39984 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_356
timestamp 1698431365
transform 1 0 41216 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_362
timestamp 1698431365
transform 1 0 41888 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_378
timestamp 1698431365
transform 1 0 43680 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_69
timestamp 1698431365
transform 1 0 9072 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_85
timestamp 1698431365
transform 1 0 10864 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_89
timestamp 1698431365
transform 1 0 11312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_91
timestamp 1698431365
transform 1 0 11536 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_111
timestamp 1698431365
transform 1 0 13776 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_138
timestamp 1698431365
transform 1 0 16800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_140
timestamp 1698431365
transform 1 0 17024 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_179
timestamp 1698431365
transform 1 0 21392 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_222
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_230
timestamp 1698431365
transform 1 0 27104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_268
timestamp 1698431365
transform 1 0 31360 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_276
timestamp 1698431365
transform 1 0 32256 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_280
timestamp 1698431365
transform 1 0 32704 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_351
timestamp 1698431365
transform 1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_372
timestamp 1698431365
transform 1 0 43008 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_380
timestamp 1698431365
transform 1 0 43904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_88
timestamp 1698431365
transform 1 0 11200 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_102
timestamp 1698431365
transform 1 0 12768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_144
timestamp 1698431365
transform 1 0 17472 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_163
timestamp 1698431365
transform 1 0 19600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_216
timestamp 1698431365
transform 1 0 25536 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_224
timestamp 1698431365
transform 1 0 26432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_226
timestamp 1698431365
transform 1 0 26656 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_253
timestamp 1698431365
transform 1 0 29680 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_261
timestamp 1698431365
transform 1 0 30576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_265
timestamp 1698431365
transform 1 0 31024 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_272
timestamp 1698431365
transform 1 0 31808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_290
timestamp 1698431365
transform 1 0 33824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_343
timestamp 1698431365
transform 1 0 39760 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_347
timestamp 1698431365
transform 1 0 40208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_373
timestamp 1698431365
transform 1 0 43120 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_375
timestamp 1698431365
transform 1 0 43344 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_53
timestamp 1698431365
transform 1 0 7280 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_61
timestamp 1698431365
transform 1 0 8176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698431365
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_109
timestamp 1698431365
transform 1 0 13552 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_126
timestamp 1698431365
transform 1 0 15456 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_313
timestamp 1698431365
transform 1 0 36400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_325
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_382
timestamp 1698431365
transform 1 0 44128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_80
timestamp 1698431365
transform 1 0 10304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_116
timestamp 1698431365
transform 1 0 14336 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_132
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_169
timestamp 1698431365
transform 1 0 20272 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_193
timestamp 1698431365
transform 1 0 22960 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_201
timestamp 1698431365
transform 1 0 23856 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_205
timestamp 1698431365
transform 1 0 24304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_294
timestamp 1698431365
transform 1 0 34272 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_296
timestamp 1698431365
transform 1 0 34496 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_310
timestamp 1698431365
transform 1 0 36064 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_356
timestamp 1698431365
transform 1 0 41216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_377
timestamp 1698431365
transform 1 0 43568 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_381
timestamp 1698431365
transform 1 0 44016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_383
timestamp 1698431365
transform 1 0 44240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_77
timestamp 1698431365
transform 1 0 9968 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_81
timestamp 1698431365
transform 1 0 10416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_118
timestamp 1698431365
transform 1 0 14560 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_126
timestamp 1698431365
transform 1 0 15456 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_160
timestamp 1698431365
transform 1 0 19264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_162
timestamp 1698431365
transform 1 0 19488 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_195
timestamp 1698431365
transform 1 0 23184 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_211
timestamp 1698431365
transform 1 0 24976 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_219
timestamp 1698431365
transform 1 0 25872 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_235
timestamp 1698431365
transform 1 0 27664 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_243
timestamp 1698431365
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_270
timestamp 1698431365
transform 1 0 31584 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_380
timestamp 1698431365
transform 1 0 43904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_110
timestamp 1698431365
transform 1 0 13664 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_132
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_197
timestamp 1698431365
transform 1 0 23408 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_201
timestamp 1698431365
transform 1 0 23856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_207
timestamp 1698431365
transform 1 0 24528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_221
timestamp 1698431365
transform 1 0 26096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_225
timestamp 1698431365
transform 1 0 26544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_277
timestamp 1698431365
transform 1 0 32368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_287
timestamp 1698431365
transform 1 0 33488 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_291
timestamp 1698431365
transform 1 0 33936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_328
timestamp 1698431365
transform 1 0 38080 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_342
timestamp 1698431365
transform 1 0 39648 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_356
timestamp 1698431365
transform 1 0 41216 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_364
timestamp 1698431365
transform 1 0 42112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_372
timestamp 1698431365
transform 1 0 43008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_99
timestamp 1698431365
transform 1 0 12432 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_136
timestamp 1698431365
transform 1 0 16576 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_140
timestamp 1698431365
transform 1 0 17024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_158
timestamp 1698431365
transform 1 0 19040 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_166
timestamp 1698431365
transform 1 0 19936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_170
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_185
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_218
timestamp 1698431365
transform 1 0 25760 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_234
timestamp 1698431365
transform 1 0 27552 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_242
timestamp 1698431365
transform 1 0 28448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_276
timestamp 1698431365
transform 1 0 32256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_280
timestamp 1698431365
transform 1 0 32704 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_288
timestamp 1698431365
transform 1 0 33600 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_292
timestamp 1698431365
transform 1 0 34048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_310
timestamp 1698431365
transform 1 0 36064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_341
timestamp 1698431365
transform 1 0 39536 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_349
timestamp 1698431365
transform 1 0 40432 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_84
timestamp 1698431365
transform 1 0 10752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_107
timestamp 1698431365
transform 1 0 13328 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_109
timestamp 1698431365
transform 1 0 13552 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_118
timestamp 1698431365
transform 1 0 14560 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_127
timestamp 1698431365
transform 1 0 15568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_131
timestamp 1698431365
transform 1 0 16016 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_150
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_188
timestamp 1698431365
transform 1 0 22400 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_228
timestamp 1698431365
transform 1 0 26880 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_232
timestamp 1698431365
transform 1 0 27328 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_274
timestamp 1698431365
transform 1 0 32032 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_278
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_286
timestamp 1698431365
transform 1 0 33376 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_288
timestamp 1698431365
transform 1 0 33600 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_334
timestamp 1698431365
transform 1 0 38752 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_363
timestamp 1698431365
transform 1 0 42000 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_379
timestamp 1698431365
transform 1 0 43792 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_383
timestamp 1698431365
transform 1 0 44240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_85
timestamp 1698431365
transform 1 0 10864 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_93
timestamp 1698431365
transform 1 0 11760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_100
timestamp 1698431365
transform 1 0 12544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_111
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_127
timestamp 1698431365
transform 1 0 15568 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_160
timestamp 1698431365
transform 1 0 19264 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_168
timestamp 1698431365
transform 1 0 20160 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_172
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_219
timestamp 1698431365
transform 1 0 25872 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_223
timestamp 1698431365
transform 1 0 26320 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_264
timestamp 1698431365
transform 1 0 30912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_268
timestamp 1698431365
transform 1 0 31360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_331
timestamp 1698431365
transform 1 0 38416 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_373
timestamp 1698431365
transform 1 0 43120 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_383
timestamp 1698431365
transform 1 0 44240 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_104
timestamp 1698431365
transform 1 0 12992 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_108
timestamp 1698431365
transform 1 0 13440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_110
timestamp 1698431365
transform 1 0 13664 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_163
timestamp 1698431365
transform 1 0 19600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_167
timestamp 1698431365
transform 1 0 20048 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_175
timestamp 1698431365
transform 1 0 20944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_177
timestamp 1698431365
transform 1 0 21168 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_196
timestamp 1698431365
transform 1 0 23296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_200
timestamp 1698431365
transform 1 0 23744 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_230
timestamp 1698431365
transform 1 0 27104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_232
timestamp 1698431365
transform 1 0 27328 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_256
timestamp 1698431365
transform 1 0 30016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_266
timestamp 1698431365
transform 1 0 31136 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_270
timestamp 1698431365
transform 1 0 31584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_321
timestamp 1698431365
transform 1 0 37296 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_325
timestamp 1698431365
transform 1 0 37744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_331
timestamp 1698431365
transform 1 0 38416 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_337
timestamp 1698431365
transform 1 0 39088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_345
timestamp 1698431365
transform 1 0 39984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_379
timestamp 1698431365
transform 1 0 43792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_381
timestamp 1698431365
transform 1 0 44016 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_69
timestamp 1698431365
transform 1 0 9072 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_85
timestamp 1698431365
transform 1 0 10864 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_93
timestamp 1698431365
transform 1 0 11760 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_97
timestamp 1698431365
transform 1 0 12208 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_111
timestamp 1698431365
transform 1 0 13776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_113
timestamp 1698431365
transform 1 0 14000 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_163
timestamp 1698431365
transform 1 0 19600 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_167
timestamp 1698431365
transform 1 0 20048 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_170
timestamp 1698431365
transform 1 0 20384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_186
timestamp 1698431365
transform 1 0 22176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_190
timestamp 1698431365
transform 1 0 22624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_194
timestamp 1698431365
transform 1 0 23072 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_210
timestamp 1698431365
transform 1 0 24864 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_214
timestamp 1698431365
transform 1 0 25312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_233
timestamp 1698431365
transform 1 0 27440 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_237
timestamp 1698431365
transform 1 0 27888 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_251
timestamp 1698431365
transform 1 0 29456 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_255
timestamp 1698431365
transform 1 0 29904 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_258
timestamp 1698431365
transform 1 0 30240 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_262
timestamp 1698431365
transform 1 0 30688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_264
timestamp 1698431365
transform 1 0 30912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_267
timestamp 1698431365
transform 1 0 31248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_271
timestamp 1698431365
transform 1 0 31696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_275
timestamp 1698431365
transform 1 0 32144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_277
timestamp 1698431365
transform 1 0 32368 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_374
timestamp 1698431365
transform 1 0 43232 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_113
timestamp 1698431365
transform 1 0 14000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_117
timestamp 1698431365
transform 1 0 14448 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_146
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_154
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_178
timestamp 1698431365
transform 1 0 21280 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_186
timestamp 1698431365
transform 1 0 22176 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_196
timestamp 1698431365
transform 1 0 23296 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_204
timestamp 1698431365
transform 1 0 24192 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_288
timestamp 1698431365
transform 1 0 33600 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_306
timestamp 1698431365
transform 1 0 35616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_308
timestamp 1698431365
transform 1 0 35840 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_343
timestamp 1698431365
transform 1 0 39760 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_354
timestamp 1698431365
transform 1 0 40992 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_376
timestamp 1698431365
transform 1 0 43456 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_53
timestamp 1698431365
transform 1 0 7280 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_61
timestamp 1698431365
transform 1 0 8176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_65
timestamp 1698431365
transform 1 0 8624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_112
timestamp 1698431365
transform 1 0 13888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_116
timestamp 1698431365
transform 1 0 14336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_143
timestamp 1698431365
transform 1 0 17360 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_147
timestamp 1698431365
transform 1 0 17808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_149
timestamp 1698431365
transform 1 0 18032 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_227
timestamp 1698431365
transform 1 0 26768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_229
timestamp 1698431365
transform 1 0 26992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_263
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_300
timestamp 1698431365
transform 1 0 34944 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_304
timestamp 1698431365
transform 1 0 35392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_306
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_309
timestamp 1698431365
transform 1 0 35952 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_313
timestamp 1698431365
transform 1 0 36400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_349
timestamp 1698431365
transform 1 0 40432 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_371
timestamp 1698431365
transform 1 0 42896 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_379
timestamp 1698431365
transform 1 0 43792 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_383
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_34
timestamp 1698431365
transform 1 0 5152 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_50
timestamp 1698431365
transform 1 0 6944 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_58
timestamp 1698431365
transform 1 0 7840 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_109
timestamp 1698431365
transform 1 0 13552 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_115
timestamp 1698431365
transform 1 0 14224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_119
timestamp 1698431365
transform 1 0 14672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_121
timestamp 1698431365
transform 1 0 14896 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_128
timestamp 1698431365
transform 1 0 15680 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_264
timestamp 1698431365
transform 1 0 30912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_314
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698431365
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_379
timestamp 1698431365
transform 1 0 43792 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_383
timestamp 1698431365
transform 1 0 44240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_45
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_49
timestamp 1698431365
transform 1 0 6832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_54
timestamp 1698431365
transform 1 0 7392 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_62
timestamp 1698431365
transform 1 0 8288 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_66
timestamp 1698431365
transform 1 0 8736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_68
timestamp 1698431365
transform 1 0 8960 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_85
timestamp 1698431365
transform 1 0 10864 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_140
timestamp 1698431365
transform 1 0 17024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_144
timestamp 1698431365
transform 1 0 17472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_148
timestamp 1698431365
transform 1 0 17920 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_152
timestamp 1698431365
transform 1 0 18368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_154
timestamp 1698431365
transform 1 0 18592 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_191
timestamp 1698431365
transform 1 0 22736 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_208
timestamp 1698431365
transform 1 0 24640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_212
timestamp 1698431365
transform 1 0 25088 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_267
timestamp 1698431365
transform 1 0 31248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_281
timestamp 1698431365
transform 1 0 32816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_285
timestamp 1698431365
transform 1 0 33264 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_289
timestamp 1698431365
transform 1 0 33712 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_296
timestamp 1698431365
transform 1 0 34496 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_333
timestamp 1698431365
transform 1 0 38640 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_383
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_34
timestamp 1698431365
transform 1 0 5152 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_74
timestamp 1698431365
transform 1 0 9632 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698431365
transform 1 0 13664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_204
timestamp 1698431365
transform 1 0 24192 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_227
timestamp 1698431365
transform 1 0 26768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_257
timestamp 1698431365
transform 1 0 30128 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_261
timestamp 1698431365
transform 1 0 30576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_265
timestamp 1698431365
transform 1 0 31024 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_273
timestamp 1698431365
transform 1 0 31920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_284
timestamp 1698431365
transform 1 0 33152 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_314
timestamp 1698431365
transform 1 0 36512 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_360
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_367
timestamp 1698431365
transform 1 0 42448 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_375
timestamp 1698431365
transform 1 0 43344 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_83
timestamp 1698431365
transform 1 0 10640 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_87
timestamp 1698431365
transform 1 0 11088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_99
timestamp 1698431365
transform 1 0 12432 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_103
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_141
timestamp 1698431365
transform 1 0 17136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_145
timestamp 1698431365
transform 1 0 17584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_149
timestamp 1698431365
transform 1 0 18032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_153
timestamp 1698431365
transform 1 0 18480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_195
timestamp 1698431365
transform 1 0 23184 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_199
timestamp 1698431365
transform 1 0 23632 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_267
timestamp 1698431365
transform 1 0 31248 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_271
timestamp 1698431365
transform 1 0 31696 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_273
timestamp 1698431365
transform 1 0 31920 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_373
timestamp 1698431365
transform 1 0 43120 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_381
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_383
timestamp 1698431365
transform 1 0 44240 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_36
timestamp 1698431365
transform 1 0 5376 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_40
timestamp 1698431365
transform 1 0 5824 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_54
timestamp 1698431365
transform 1 0 7392 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_67
timestamp 1698431365
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_78
timestamp 1698431365
transform 1 0 10080 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_101
timestamp 1698431365
transform 1 0 12656 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_113
timestamp 1698431365
transform 1 0 14000 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_115
timestamp 1698431365
transform 1 0 14224 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_124
timestamp 1698431365
transform 1 0 15232 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_134
timestamp 1698431365
transform 1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_147
timestamp 1698431365
transform 1 0 17808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_149
timestamp 1698431365
transform 1 0 18032 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_156
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_164
timestamp 1698431365
transform 1 0 19712 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_168
timestamp 1698431365
transform 1 0 20160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_170
timestamp 1698431365
transform 1 0 20384 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_179
timestamp 1698431365
transform 1 0 21392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_199
timestamp 1698431365
transform 1 0 23632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_201
timestamp 1698431365
transform 1 0 23856 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_218
timestamp 1698431365
transform 1 0 25760 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_226
timestamp 1698431365
transform 1 0 26656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_230
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_234
timestamp 1698431365
transform 1 0 27552 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_236
timestamp 1698431365
transform 1 0 27776 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_260
timestamp 1698431365
transform 1 0 30464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_268
timestamp 1698431365
transform 1 0 31360 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_288
timestamp 1698431365
transform 1 0 33600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_290
timestamp 1698431365
transform 1 0 33824 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_317
timestamp 1698431365
transform 1 0 36848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_321
timestamp 1698431365
transform 1 0 37296 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_337
timestamp 1698431365
transform 1 0 39088 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_341
timestamp 1698431365
transform 1 0 39536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_343
timestamp 1698431365
transform 1 0 39760 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_348
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_377
timestamp 1698431365
transform 1 0 43568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_381
timestamp 1698431365
transform 1 0 44016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_383
timestamp 1698431365
transform 1 0 44240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_10
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_14
timestamp 1698431365
transform 1 0 2912 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_19
timestamp 1698431365
transform 1 0 3472 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_43
timestamp 1698431365
transform 1 0 6160 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_56
timestamp 1698431365
transform 1 0 7616 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_88
timestamp 1698431365
transform 1 0 11200 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_92
timestamp 1698431365
transform 1 0 11648 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_102
timestamp 1698431365
transform 1 0 12768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_111
timestamp 1698431365
transform 1 0 13776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_190
timestamp 1698431365
transform 1 0 22624 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_222
timestamp 1698431365
transform 1 0 26208 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_226
timestamp 1698431365
transform 1 0 26656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_276
timestamp 1698431365
transform 1 0 32256 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698431365
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_321
timestamp 1698431365
transform 1 0 37296 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_337
timestamp 1698431365
transform 1 0 39088 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_345
timestamp 1698431365
transform 1 0 39984 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_4
timestamp 1698431365
transform 1 0 1792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_39
timestamp 1698431365
transform 1 0 5712 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_55
timestamp 1698431365
transform 1 0 7504 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_63
timestamp 1698431365
transform 1 0 8400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_92
timestamp 1698431365
transform 1 0 11648 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_127
timestamp 1698431365
transform 1 0 15568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_135
timestamp 1698431365
transform 1 0 16464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_193
timestamp 1698431365
transform 1 0 22960 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_216
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_231
timestamp 1698431365
transform 1 0 27216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_239
timestamp 1698431365
transform 1 0 28112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_288
timestamp 1698431365
transform 1 0 33600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_298
timestamp 1698431365
transform 1 0 34720 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_343
timestamp 1698431365
transform 1 0 39760 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_18
timestamp 1698431365
transform 1 0 3360 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_22
timestamp 1698431365
transform 1 0 3808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_24
timestamp 1698431365
transform 1 0 4032 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_49
timestamp 1698431365
transform 1 0 6832 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_57
timestamp 1698431365
transform 1 0 7728 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_61
timestamp 1698431365
transform 1 0 8176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_97
timestamp 1698431365
transform 1 0 12208 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_119
timestamp 1698431365
transform 1 0 14672 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_153
timestamp 1698431365
transform 1 0 18480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_155
timestamp 1698431365
transform 1 0 18704 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_162
timestamp 1698431365
transform 1 0 19488 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_193
timestamp 1698431365
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_197
timestamp 1698431365
transform 1 0 23408 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_205
timestamp 1698431365
transform 1 0 24304 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_209
timestamp 1698431365
transform 1 0 24752 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_211
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698431365
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_264
timestamp 1698431365
transform 1 0 30912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_266
timestamp 1698431365
transform 1 0 31136 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_326
timestamp 1698431365
transform 1 0 37856 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_361
timestamp 1698431365
transform 1 0 41776 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_379
timestamp 1698431365
transform 1 0 43792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_381
timestamp 1698431365
transform 1 0 44016 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_18
timestamp 1698431365
transform 1 0 3360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_20
timestamp 1698431365
transform 1 0 3584 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_59
timestamp 1698431365
transform 1 0 7952 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_67
timestamp 1698431365
transform 1 0 8848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_110
timestamp 1698431365
transform 1 0 13664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_121
timestamp 1698431365
transform 1 0 14896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_123
timestamp 1698431365
transform 1 0 15120 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_152
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_194
timestamp 1698431365
transform 1 0 23072 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_246
timestamp 1698431365
transform 1 0 28896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_250
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_254
timestamp 1698431365
transform 1 0 29792 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_262
timestamp 1698431365
transform 1 0 30688 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_269
timestamp 1698431365
transform 1 0 31472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698431365
transform 1 0 31920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698431365
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_321
timestamp 1698431365
transform 1 0 37296 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_337
timestamp 1698431365
transform 1 0 39088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_341
timestamp 1698431365
transform 1 0 39536 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_354
timestamp 1698431365
transform 1 0 40992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_368
timestamp 1698431365
transform 1 0 42560 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_18
timestamp 1698431365
transform 1 0 3360 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_26
timestamp 1698431365
transform 1 0 4256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_39
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_88
timestamp 1698431365
transform 1 0 11200 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_90
timestamp 1698431365
transform 1 0 11424 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_95
timestamp 1698431365
transform 1 0 11984 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_116
timestamp 1698431365
transform 1 0 14336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_120
timestamp 1698431365
transform 1 0 14784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_122
timestamp 1698431365
transform 1 0 15008 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_152
timestamp 1698431365
transform 1 0 18368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_156
timestamp 1698431365
transform 1 0 18816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_158
timestamp 1698431365
transform 1 0 19040 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_161
timestamp 1698431365
transform 1 0 19376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_165
timestamp 1698431365
transform 1 0 19824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_192
timestamp 1698431365
transform 1 0 22848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_196
timestamp 1698431365
transform 1 0 23296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_198
timestamp 1698431365
transform 1 0 23520 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_205
timestamp 1698431365
transform 1 0 24304 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_213
timestamp 1698431365
transform 1 0 25200 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_220
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_236
timestamp 1698431365
transform 1 0 27776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_238
timestamp 1698431365
transform 1 0 28000 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_249
timestamp 1698431365
transform 1 0 29232 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_285
timestamp 1698431365
transform 1 0 33264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_287
timestamp 1698431365
transform 1 0 33488 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_308
timestamp 1698431365
transform 1 0 35840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_326
timestamp 1698431365
transform 1 0 37856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_330
timestamp 1698431365
transform 1 0 38304 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_369
timestamp 1698431365
transform 1 0 42672 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_377
timestamp 1698431365
transform 1 0 43568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_34
timestamp 1698431365
transform 1 0 5152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_67
timestamp 1698431365
transform 1 0 8848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_80
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_82
timestamp 1698431365
transform 1 0 10528 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_117
timestamp 1698431365
transform 1 0 14448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698431365
transform 1 0 16240 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698431365
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_144
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_164
timestamp 1698431365
transform 1 0 19712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_166
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_185
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_201
timestamp 1698431365
transform 1 0 23856 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_250
timestamp 1698431365
transform 1 0 29344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_254
timestamp 1698431365
transform 1 0 29792 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_275
timestamp 1698431365
transform 1 0 32144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_298
timestamp 1698431365
transform 1 0 34720 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_320
timestamp 1698431365
transform 1 0 37184 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_328
timestamp 1698431365
transform 1 0 38080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_338
timestamp 1698431365
transform 1 0 39200 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_377
timestamp 1698431365
transform 1 0 43568 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_78
timestamp 1698431365
transform 1 0 10080 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_94
timestamp 1698431365
transform 1 0 11872 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_158
timestamp 1698431365
transform 1 0 19040 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_167
timestamp 1698431365
transform 1 0 20048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_193
timestamp 1698431365
transform 1 0 22960 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_230
timestamp 1698431365
transform 1 0 27104 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_238
timestamp 1698431365
transform 1 0 28000 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_288
timestamp 1698431365
transform 1 0 33600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_296
timestamp 1698431365
transform 1 0 34496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_298
timestamp 1698431365
transform 1 0 34720 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_308
timestamp 1698431365
transform 1 0 35840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_341
timestamp 1698431365
transform 1 0 39536 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_349
timestamp 1698431365
transform 1 0 40432 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_34
timestamp 1698431365
transform 1 0 5152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_42
timestamp 1698431365
transform 1 0 6048 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_46
timestamp 1698431365
transform 1 0 6496 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_48
timestamp 1698431365
transform 1 0 6720 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_67
timestamp 1698431365
transform 1 0 8848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_114
timestamp 1698431365
transform 1 0 14112 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_130
timestamp 1698431365
transform 1 0 15904 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_146
timestamp 1698431365
transform 1 0 17696 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_185
timestamp 1698431365
transform 1 0 22064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_191
timestamp 1698431365
transform 1 0 22736 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698431365
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_218
timestamp 1698431365
transform 1 0 25760 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_234
timestamp 1698431365
transform 1 0 27552 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_238
timestamp 1698431365
transform 1 0 28000 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_242
timestamp 1698431365
transform 1 0 28448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_244
timestamp 1698431365
transform 1 0 28672 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_286
timestamp 1698431365
transform 1 0 33376 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_333
timestamp 1698431365
transform 1 0 38640 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_354
timestamp 1698431365
transform 1 0 40992 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_374
timestamp 1698431365
transform 1 0 43232 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_382
timestamp 1698431365
transform 1 0 44128 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_49
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_51
timestamp 1698431365
transform 1 0 7056 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_60
timestamp 1698431365
transform 1 0 8064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_64
timestamp 1698431365
transform 1 0 8512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_68
timestamp 1698431365
transform 1 0 8960 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_70
timestamp 1698431365
transform 1 0 9184 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_123
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_181
timestamp 1698431365
transform 1 0 21616 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_191
timestamp 1698431365
transform 1 0 22736 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_199
timestamp 1698431365
transform 1 0 23632 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_205
timestamp 1698431365
transform 1 0 24304 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_209
timestamp 1698431365
transform 1 0 24752 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_220
timestamp 1698431365
transform 1 0 25984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_224
timestamp 1698431365
transform 1 0 26432 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_232
timestamp 1698431365
transform 1 0 27328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_236
timestamp 1698431365
transform 1 0 27776 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_251
timestamp 1698431365
transform 1 0 29456 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_267
timestamp 1698431365
transform 1 0 31248 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_275
timestamp 1698431365
transform 1 0 32144 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_279
timestamp 1698431365
transform 1 0 32592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_330
timestamp 1698431365
transform 1 0 38304 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_344
timestamp 1698431365
transform 1 0 39872 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_352
timestamp 1698431365
transform 1 0 40768 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_360
timestamp 1698431365
transform 1 0 41664 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_367
timestamp 1698431365
transform 1 0 42448 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_375
timestamp 1698431365
transform 1 0 43344 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_379
timestamp 1698431365
transform 1 0 43792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_34
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_50
timestamp 1698431365
transform 1 0 6944 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_58
timestamp 1698431365
transform 1 0 7840 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_117
timestamp 1698431365
transform 1 0 14448 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_133
timestamp 1698431365
transform 1 0 16240 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_137
timestamp 1698431365
transform 1 0 16688 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_154
timestamp 1698431365
transform 1 0 18592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_156
timestamp 1698431365
transform 1 0 18816 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_167
timestamp 1698431365
transform 1 0 20048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_171
timestamp 1698431365
transform 1 0 20496 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_216
timestamp 1698431365
transform 1 0 25536 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_232
timestamp 1698431365
transform 1 0 27328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_236
timestamp 1698431365
transform 1 0 27776 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_252
timestamp 1698431365
transform 1 0 29568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_260
timestamp 1698431365
transform 1 0 30464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_266
timestamp 1698431365
transform 1 0 31136 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698431365
transform 1 0 32032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_290
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_329
timestamp 1698431365
transform 1 0 38192 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_331
timestamp 1698431365
transform 1 0 38416 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_345
timestamp 1698431365
transform 1 0 39984 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_349
timestamp 1698431365
transform 1 0 40432 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_69
timestamp 1698431365
transform 1 0 9072 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_102
timestamp 1698431365
transform 1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_123
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_165
timestamp 1698431365
transform 1 0 19824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_181
timestamp 1698431365
transform 1 0 21616 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_197
timestamp 1698431365
transform 1 0 23408 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_201
timestamp 1698431365
transform 1 0 23856 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_237
timestamp 1698431365
transform 1 0 27888 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_280
timestamp 1698431365
transform 1 0 32704 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_296
timestamp 1698431365
transform 1 0 34496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_321
timestamp 1698431365
transform 1 0 37296 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_325
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_327
timestamp 1698431365
transform 1 0 37968 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_340
timestamp 1698431365
transform 1 0 39424 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_348
timestamp 1698431365
transform 1 0 40320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_80
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_97
timestamp 1698431365
transform 1 0 12208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_101
timestamp 1698431365
transform 1 0 12656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_103
timestamp 1698431365
transform 1 0 12880 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_148
timestamp 1698431365
transform 1 0 17920 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_187
timestamp 1698431365
transform 1 0 22288 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_195
timestamp 1698431365
transform 1 0 23184 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_199
timestamp 1698431365
transform 1 0 23632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_201
timestamp 1698431365
transform 1 0 23856 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_243
timestamp 1698431365
transform 1 0 28560 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_368
timestamp 1698431365
transform 1 0 42560 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_374
timestamp 1698431365
transform 1 0 43232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_53
timestamp 1698431365
transform 1 0 7280 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_83
timestamp 1698431365
transform 1 0 10640 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_99
timestamp 1698431365
transform 1 0 12432 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_103
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_123
timestamp 1698431365
transform 1 0 15120 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_127
timestamp 1698431365
transform 1 0 15568 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_162
timestamp 1698431365
transform 1 0 19488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_166
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_193
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_201
timestamp 1698431365
transform 1 0 23856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_251
timestamp 1698431365
transform 1 0 29456 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_292
timestamp 1698431365
transform 1 0 34048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_296
timestamp 1698431365
transform 1 0 34496 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_349
timestamp 1698431365
transform 1 0 40432 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_353
timestamp 1698431365
transform 1 0 40880 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_383
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_34
timestamp 1698431365
transform 1 0 5152 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_38
timestamp 1698431365
transform 1 0 5600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_40
timestamp 1698431365
transform 1 0 5824 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_108
timestamp 1698431365
transform 1 0 13440 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_110
timestamp 1698431365
transform 1 0 13664 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_115
timestamp 1698431365
transform 1 0 14224 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_119
timestamp 1698431365
transform 1 0 14672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_125
timestamp 1698431365
transform 1 0 15344 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_129
timestamp 1698431365
transform 1 0 15792 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_131
timestamp 1698431365
transform 1 0 16016 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_149
timestamp 1698431365
transform 1 0 18032 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_154
timestamp 1698431365
transform 1 0 18592 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_162
timestamp 1698431365
transform 1 0 19488 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_193
timestamp 1698431365
transform 1 0 22960 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_197
timestamp 1698431365
transform 1 0 23408 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_247
timestamp 1698431365
transform 1 0 29008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_266
timestamp 1698431365
transform 1 0 31136 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_270
timestamp 1698431365
transform 1 0 31584 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_288
timestamp 1698431365
transform 1 0 33600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_325
timestamp 1698431365
transform 1 0 37744 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_341
timestamp 1698431365
transform 1 0 39536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_343
timestamp 1698431365
transform 1 0 39760 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_381
timestamp 1698431365
transform 1 0 44016 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_383
timestamp 1698431365
transform 1 0 44240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_143
timestamp 1698431365
transform 1 0 17360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_145
timestamp 1698431365
transform 1 0 17584 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_183
timestamp 1698431365
transform 1 0 21840 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_191
timestamp 1698431365
transform 1 0 22736 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_195
timestamp 1698431365
transform 1 0 23184 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_269
timestamp 1698431365
transform 1 0 31472 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_303
timestamp 1698431365
transform 1 0 35280 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_331
timestamp 1698431365
transform 1 0 38416 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_335
timestamp 1698431365
transform 1 0 38864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_337
timestamp 1698431365
transform 1 0 39088 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_380
timestamp 1698431365
transform 1 0 43904 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_34
timestamp 1698431365
transform 1 0 5152 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_50
timestamp 1698431365
transform 1 0 6944 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_58
timestamp 1698431365
transform 1 0 7840 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_60
timestamp 1698431365
transform 1 0 8064 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_67
timestamp 1698431365
transform 1 0 8848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_123
timestamp 1698431365
transform 1 0 15120 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_131
timestamp 1698431365
transform 1 0 16016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_158
timestamp 1698431365
transform 1 0 19040 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_162
timestamp 1698431365
transform 1 0 19488 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_173
timestamp 1698431365
transform 1 0 20720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_181
timestamp 1698431365
transform 1 0 21616 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_197
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_201
timestamp 1698431365
transform 1 0 23856 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_222
timestamp 1698431365
transform 1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_224
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_231
timestamp 1698431365
transform 1 0 27216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_235
timestamp 1698431365
transform 1 0 27664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_239
timestamp 1698431365
transform 1 0 28112 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_255
timestamp 1698431365
transform 1 0 29904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_273
timestamp 1698431365
transform 1 0 31920 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_277
timestamp 1698431365
transform 1 0 32368 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_288
timestamp 1698431365
transform 1 0 33600 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_296
timestamp 1698431365
transform 1 0 34496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_381
timestamp 1698431365
transform 1 0 44016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_383
timestamp 1698431365
transform 1 0 44240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_45
timestamp 1698431365
transform 1 0 6384 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_49
timestamp 1698431365
transform 1 0 6832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_80
timestamp 1698431365
transform 1 0 10304 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_84
timestamp 1698431365
transform 1 0 10752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_92
timestamp 1698431365
transform 1 0 11648 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_100
timestamp 1698431365
transform 1 0 12544 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_149
timestamp 1698431365
transform 1 0 18032 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_153
timestamp 1698431365
transform 1 0 18480 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_169
timestamp 1698431365
transform 1 0 20272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_173
timestamp 1698431365
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_255
timestamp 1698431365
transform 1 0 29904 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_259
timestamp 1698431365
transform 1 0 30352 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_261
timestamp 1698431365
transform 1 0 30576 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_275
timestamp 1698431365
transform 1 0 32144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_308
timestamp 1698431365
transform 1 0 35840 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_327
timestamp 1698431365
transform 1 0 37968 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_34
timestamp 1698431365
transform 1 0 5152 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_38
timestamp 1698431365
transform 1 0 5600 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_40
timestamp 1698431365
transform 1 0 5824 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_84
timestamp 1698431365
transform 1 0 10752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_124
timestamp 1698431365
transform 1 0 15232 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_135
timestamp 1698431365
transform 1 0 16464 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_146
timestamp 1698431365
transform 1 0 17696 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_153
timestamp 1698431365
transform 1 0 18480 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_161
timestamp 1698431365
transform 1 0 19376 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_165
timestamp 1698431365
transform 1 0 19824 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_195
timestamp 1698431365
transform 1 0 23184 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_203
timestamp 1698431365
transform 1 0 24080 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_240
timestamp 1698431365
transform 1 0 28224 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_255
timestamp 1698431365
transform 1 0 29904 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_271
timestamp 1698431365
transform 1 0 31696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_273
timestamp 1698431365
transform 1 0 31920 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_292
timestamp 1698431365
transform 1 0 34048 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_329
timestamp 1698431365
transform 1 0 38192 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_380
timestamp 1698431365
transform 1 0 43904 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_84
timestamp 1698431365
transform 1 0 10752 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_100
timestamp 1698431365
transform 1 0 12544 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_115
timestamp 1698431365
transform 1 0 14224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_158
timestamp 1698431365
transform 1 0 19040 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_206
timestamp 1698431365
transform 1 0 24416 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_259
timestamp 1698431365
transform 1 0 30352 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_267
timestamp 1698431365
transform 1 0 31248 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_298
timestamp 1698431365
transform 1 0 34720 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_302
timestamp 1698431365
transform 1 0 35168 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_329
timestamp 1698431365
transform 1 0 38192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_336
timestamp 1698431365
transform 1 0 38976 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_356
timestamp 1698431365
transform 1 0 41216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_34
timestamp 1698431365
transform 1 0 5152 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_50
timestamp 1698431365
transform 1 0 6944 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_54
timestamp 1698431365
transform 1 0 7392 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_56
timestamp 1698431365
transform 1 0 7616 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_63
timestamp 1698431365
transform 1 0 8400 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_74
timestamp 1698431365
transform 1 0 9632 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_93
timestamp 1698431365
transform 1 0 11760 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_97
timestamp 1698431365
transform 1 0 12208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_135
timestamp 1698431365
transform 1 0 16464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_269
timestamp 1698431365
transform 1 0 31472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_271
timestamp 1698431365
transform 1 0 31696 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_327
timestamp 1698431365
transform 1 0 37968 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_335
timestamp 1698431365
transform 1 0 38864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_337
timestamp 1698431365
transform 1 0 39088 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_358
timestamp 1698431365
transform 1 0 41440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_377
timestamp 1698431365
transform 1 0 43568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_381
timestamp 1698431365
transform 1 0 44016 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_383
timestamp 1698431365
transform 1 0 44240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_53
timestamp 1698431365
transform 1 0 7280 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_61
timestamp 1698431365
transform 1 0 8176 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_92
timestamp 1698431365
transform 1 0 11648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_100
timestamp 1698431365
transform 1 0 12544 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_123
timestamp 1698431365
transform 1 0 15120 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_181
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_257
timestamp 1698431365
transform 1 0 30128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_261
timestamp 1698431365
transform 1 0 30576 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_297
timestamp 1698431365
transform 1 0 34608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_313
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_335
timestamp 1698431365
transform 1 0 38864 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_347
timestamp 1698431365
transform 1 0 40208 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_86
timestamp 1698431365
transform 1 0 10976 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_118
timestamp 1698431365
transform 1 0 14560 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_126
timestamp 1698431365
transform 1 0 15456 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_165
timestamp 1698431365
transform 1 0 19824 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_200
timestamp 1698431365
transform 1 0 23744 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_255
timestamp 1698431365
transform 1 0 29904 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_277
timestamp 1698431365
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_290
timestamp 1698431365
transform 1 0 33824 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_298
timestamp 1698431365
transform 1 0 34720 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_302
timestamp 1698431365
transform 1 0 35168 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_381
timestamp 1698431365
transform 1 0 44016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_383
timestamp 1698431365
transform 1 0 44240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_45
timestamp 1698431365
transform 1 0 6384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_49
timestamp 1698431365
transform 1 0 6832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_51
timestamp 1698431365
transform 1 0 7056 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_81
timestamp 1698431365
transform 1 0 10416 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_97
timestamp 1698431365
transform 1 0 12208 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_123
timestamp 1698431365
transform 1 0 15120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_159
timestamp 1698431365
transform 1 0 19152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_163
timestamp 1698431365
transform 1 0 19600 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_193
timestamp 1698431365
transform 1 0 22960 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_263
timestamp 1698431365
transform 1 0 30800 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_271
timestamp 1698431365
transform 1 0 31696 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_301
timestamp 1698431365
transform 1 0 35056 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_309
timestamp 1698431365
transform 1 0 35952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_383
timestamp 1698431365
transform 1 0 44240 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_216
timestamp 1698431365
transform 1 0 25536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_218
timestamp 1698431365
transform 1 0 25760 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_241
timestamp 1698431365
transform 1 0 28336 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_249
timestamp 1698431365
transform 1 0 29232 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_258
timestamp 1698431365
transform 1 0 30240 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_274
timestamp 1698431365
transform 1 0 32032 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_286
timestamp 1698431365
transform 1 0 33376 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_293
timestamp 1698431365
transform 1 0 34160 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_309
timestamp 1698431365
transform 1 0 35952 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_313
timestamp 1698431365
transform 1 0 36400 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_320
timestamp 1698431365
transform 1 0 37184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_322
timestamp 1698431365
transform 1 0 37408 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_343
timestamp 1698431365
transform 1 0 39760 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_347
timestamp 1698431365
transform 1 0 40208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_263
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_271
timestamp 1698431365
transform 1 0 31696 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_274
timestamp 1698431365
transform 1 0 32032 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_278
timestamp 1698431365
transform 1 0 32480 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_280
timestamp 1698431365
transform 1 0 32704 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_306
timestamp 1698431365
transform 1 0 35616 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1698431365
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_323
timestamp 1698431365
transform 1 0 37520 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_339
timestamp 1698431365
transform 1 0 39312 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_343
timestamp 1698431365
transform 1 0 39760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_381
timestamp 1698431365
transform 1 0 44016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_383
timestamp 1698431365
transform 1 0 44240 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_228
timestamp 1698431365
transform 1 0 26880 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_315
timestamp 1698431365
transform 1 0 36624 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_323
timestamp 1698431365
transform 1 0 37520 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_347
timestamp 1698431365
transform 1 0 40208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_349
timestamp 1698431365
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_209
timestamp 1698431365
transform 1 0 24752 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_313
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_351
timestamp 1698431365
transform 1 0 40656 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_353
timestamp 1698431365
transform 1 0 40880 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_383
timestamp 1698431365
transform 1 0 44240 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_220
timestamp 1698431365
transform 1 0 25984 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_224
timestamp 1698431365
transform 1 0 26432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_263
timestamp 1698431365
transform 1 0 30800 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_267
timestamp 1698431365
transform 1 0 31248 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_323
timestamp 1698431365
transform 1 0 37520 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_381
timestamp 1698431365
transform 1 0 44016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_383
timestamp 1698431365
transform 1 0 44240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_259
timestamp 1698431365
transform 1 0 30352 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_267
timestamp 1698431365
transform 1 0 31248 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_269
timestamp 1698431365
transform 1 0 31472 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_312
timestamp 1698431365
transform 1 0 36288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_36
timestamp 1698431365
transform 1 0 5376 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_70
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_104
timestamp 1698431365
transform 1 0 12992 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_138
timestamp 1698431365
transform 1 0 16800 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_172
timestamp 1698431365
transform 1 0 20608 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_240
timestamp 1698431365
transform 1 0 28224 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_274
timestamp 1698431365
transform 1 0 32032 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_286
timestamp 1698431365
transform 1 0 33376 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_295
timestamp 1698431365
transform 1 0 34384 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_303
timestamp 1698431365
transform 1 0 35280 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_305
timestamp 1698431365
transform 1 0 35504 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_308
timestamp 1698431365
transform 1 0 35840 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_342
timestamp 1698431365
transform 1 0 39648 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_346
timestamp 1698431365
transform 1 0 40096 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_381
timestamp 1698431365
transform 1 0 44016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_383
timestamp 1698431365
transform 1 0 44240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 44352 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2
timestamp 1698431365
transform -1 0 44352 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform -1 0 44352 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform -1 0 44352 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 44352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 44352 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698431365
transform -1 0 44352 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform -1 0 44352 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44352 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698431365
transform -1 0 44352 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698431365
transform 1 0 41440 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698431365
transform -1 0 44352 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform -1 0 43232 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_50 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 44576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 44576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 44576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 44576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 44576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 44576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 44576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 44576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 44576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_60
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 44576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 44576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 44576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 44576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 44576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 44576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 44576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 44576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 44576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 44576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 44576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 44576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 44576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 44576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 44576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 44576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 44576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 44576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 44576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 44576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 44576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 44576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 44576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 44576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 44576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 44576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 44576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 44576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 44576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 44576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 44576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 44576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 44576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 44576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 44576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 44576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 44576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 44576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_111
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_112
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_113
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_114
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_115
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_117
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_118
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_119
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_120
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_121
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_122
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_123
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_124
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_125
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_126
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_127
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_128
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_129
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_130
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_131
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_132
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_133
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_134
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_135
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_136
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_137
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_138
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_139
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_140
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_141
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_142
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_143
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_144
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_145
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_146
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_147
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_148
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_149
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_150
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_151
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_152
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_153
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_154
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_155
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_156
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_157
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_158
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_159
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_160
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_161
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_162
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_163
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_164
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_165
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_166
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_167
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_168
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_169
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_170
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_171
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_172
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_173
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_174
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_175
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_176
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_177
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_178
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_179
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_180
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_181
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_182
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_183
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_184
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_185
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_186
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_187
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_188
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_189
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_190
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_191
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_192
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_193
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_194
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_195
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_196
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_197
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_198
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_199
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_200
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_201
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_202
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_204
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_205
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_209
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_210
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_212
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_213
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_214
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_215
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_216
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_217
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_218
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_219
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_220
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_221
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_222
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_223
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_224
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_225
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_226
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_227
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_228
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_229
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_230
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_231
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_232
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_233
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_234
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_235
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_236
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_237
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_238
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_239
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_240
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_241
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_242
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_243
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_244
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_245
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_246
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_247
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_248
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_249
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_250
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_251
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_252
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_253
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_254
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_255
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_256
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_257
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_258
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_259
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_260
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_261
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_262
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_263
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_264
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_265
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_266
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_267
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_268
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_269
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_270
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_271
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_272
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_273
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_274
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_275
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_276
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_277
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_278
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_279
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_280
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_281
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_282
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_283
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_284
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_285
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_286
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_287
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_288
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_289
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_290
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_291
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_292
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_293
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_294
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_295
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_296
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_297
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_298
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_299
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_300
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_301
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_302
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_303
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_304
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_305
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_306
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_307
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_308
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_309
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_310
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_311
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_312
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_313
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_314
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_315
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_316
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_317
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_318
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_319
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_320
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_321
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_322
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_323
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_324
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_325
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_326
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_327
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_328
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_329
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_330
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_331
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_332
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_333
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_334
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_335
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_336
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_337
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_338
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_339
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_340
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_341
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_342
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_343
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_344
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_345
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_346
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_347
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_348
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_349
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_350
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_351
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_352
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_353
timestamp 1698431365
transform 1 0 12768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_354
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_355
timestamp 1698431365
transform 1 0 20384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_356
timestamp 1698431365
transform 1 0 24192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_357
timestamp 1698431365
transform 1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_358
timestamp 1698431365
transform 1 0 31808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_359
timestamp 1698431365
transform 1 0 35616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_360
timestamp 1698431365
transform 1 0 39424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_361
timestamp 1698431365
transform 1 0 43232 0 -1 42336
box -86 -86 310 870
<< labels >>
flabel metal3 s 45200 2688 46000 2800 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 45200 9408 46000 9520 0 FreeSans 448 0 0 0 io_in[0]
port 1 nsew signal input
flabel metal3 s 45200 12768 46000 12880 0 FreeSans 448 0 0 0 io_in[1]
port 2 nsew signal input
flabel metal3 s 45200 16128 46000 16240 0 FreeSans 448 0 0 0 io_in[2]
port 3 nsew signal input
flabel metal3 s 45200 19488 46000 19600 0 FreeSans 448 0 0 0 io_in[3]
port 4 nsew signal input
flabel metal3 s 45200 22848 46000 22960 0 FreeSans 448 0 0 0 io_in[4]
port 5 nsew signal input
flabel metal3 s 45200 26208 46000 26320 0 FreeSans 448 0 0 0 io_in[5]
port 6 nsew signal input
flabel metal3 s 45200 29568 46000 29680 0 FreeSans 448 0 0 0 io_out[0]
port 7 nsew signal tristate
flabel metal3 s 45200 32928 46000 33040 0 FreeSans 448 0 0 0 io_out[1]
port 8 nsew signal tristate
flabel metal3 s 45200 36288 46000 36400 0 FreeSans 448 0 0 0 io_out[2]
port 9 nsew signal tristate
flabel metal3 s 45200 39648 46000 39760 0 FreeSans 448 0 0 0 io_out[3]
port 10 nsew signal tristate
flabel metal3 s 45200 43008 46000 43120 0 FreeSans 448 0 0 0 io_out[4]
port 11 nsew signal tristate
flabel metal3 s 45200 6048 46000 6160 0 FreeSans 448 0 0 0 rst_n
port 12 nsew signal input
flabel metal4 s 4448 3076 4768 42396 0 FreeSans 1280 90 0 0 vdd
port 13 nsew power bidirectional
flabel metal4 s 35168 3076 35488 42396 0 FreeSans 1280 90 0 0 vdd
port 13 nsew power bidirectional
flabel metal4 s 19808 3076 20128 42396 0 FreeSans 1280 90 0 0 vss
port 14 nsew ground bidirectional
rlabel metal1 22960 41552 22960 41552 0 vdd
rlabel metal1 22960 42336 22960 42336 0 vss
rlabel metal2 30968 29288 30968 29288 0 CIRCUIT_2223.CLK
rlabel metal2 25816 13720 25816 13720 0 CIRCUIT_2223.GATES_1.input1\[0\]
rlabel metal3 23688 15176 23688 15176 0 CIRCUIT_2223.GATES_1.input1\[1\]
rlabel metal2 22344 16072 22344 16072 0 CIRCUIT_2223.GATES_1.input1\[2\]
rlabel metal2 25704 16912 25704 16912 0 CIRCUIT_2223.GATES_1.input1\[3\]
rlabel metal2 24024 25984 24024 25984 0 CIRCUIT_2223.GATES_11.input2
rlabel metal2 18536 24416 18536 24416 0 CIRCUIT_2223.GATES_11.result
rlabel metal3 27048 27272 27048 27272 0 CIRCUIT_2223.GATES_2.input2
rlabel metal3 27832 28616 27832 28616 0 CIRCUIT_2223.GATES_3.input2
rlabel metal2 25816 33040 25816 33040 0 CIRCUIT_2223.GATES_4.input1\[0\]
rlabel metal2 25256 35168 25256 35168 0 CIRCUIT_2223.GATES_4.input1\[1\]
rlabel metal2 24136 34832 24136 34832 0 CIRCUIT_2223.GATES_4.input1\[2\]
rlabel metal3 25032 32536 25032 32536 0 CIRCUIT_2223.GATES_4.input1\[3\]
rlabel metal2 27384 31836 27384 31836 0 CIRCUIT_2223.GATES_5.input2
rlabel metal2 16744 25760 16744 25760 0 CIRCUIT_2223.MEMORY_18.clock
rlabel metal2 16632 27160 16632 27160 0 CIRCUIT_2223.MEMORY_18.d
rlabel metal2 16688 27832 16688 27832 0 CIRCUIT_2223.MEMORY_18.s_currentState
rlabel metal2 16072 28168 16072 28168 0 CIRCUIT_2223.MEMORY_19.d
rlabel metal3 13496 29288 13496 29288 0 CIRCUIT_2223.MEMORY_19.s_currentState
rlabel metal2 15064 29904 15064 29904 0 CIRCUIT_2223.MEMORY_20.d
rlabel metal2 15176 29904 15176 29904 0 CIRCUIT_2223.MEMORY_20.s_currentState
rlabel metal2 16408 28896 16408 28896 0 CIRCUIT_2223.MEMORY_21.d
rlabel metal2 19208 29008 19208 29008 0 CIRCUIT_2223.MEMORY_21.s_currentState
rlabel metal2 20216 27552 20216 27552 0 CIRCUIT_2223.MEMORY_22.d
rlabel metal2 20328 27440 20328 27440 0 CIRCUIT_2223.MEMORY_22.s_currentState
rlabel metal2 24136 25872 24136 25872 0 CIRCUIT_2223.MEMORY_23.s_currentState
rlabel metal3 18480 24696 18480 24696 0 CIRCUIT_2223.MEMORY_24.d
rlabel metal3 21168 24920 21168 24920 0 CIRCUIT_2223.MEMORY_24.s_currentState
rlabel metal2 18312 24192 18312 24192 0 CIRCUIT_2223.MEMORY_25.d
rlabel metal2 15736 24696 15736 24696 0 CIRCUIT_2223.MEMORY_25.s_currentState
rlabel metal2 17528 25928 17528 25928 0 CIRCUIT_2223.MEMORY_26.s_currentState
rlabel metal2 26880 31752 26880 31752 0 CIRCUIT_2223.s_logisimNet48
rlabel metal2 8456 33824 8456 33824 0 CIRCUIT_2223.tone_generator_1.GATES_1.result
rlabel metal2 8232 33432 8232 33432 0 CIRCUIT_2223.tone_generator_1.GATES_2.result
rlabel metal2 8288 29512 8288 29512 0 CIRCUIT_2223.tone_generator_1.GATES_3.result
rlabel metal2 6104 29008 6104 29008 0 CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState
rlabel metal2 10472 29064 10472 29064 0 CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState
rlabel metal3 12376 29624 12376 29624 0 CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState
rlabel metal2 14504 31472 14504 31472 0 CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState
rlabel metal3 20524 32424 20524 32424 0 CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState
rlabel metal3 13888 32536 13888 32536 0 CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState
rlabel metal2 16296 35392 16296 35392 0 CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState
rlabel metal2 17752 33712 17752 33712 0 CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState
rlabel metal2 14616 34216 14616 34216 0 CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState
rlabel metal2 21000 35112 21000 35112 0 CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState
rlabel metal2 21056 34328 21056 34328 0 CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState
rlabel metal2 7336 35784 7336 35784 0 CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState
rlabel metal2 10584 34552 10584 34552 0 CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState
rlabel metal2 10584 32984 10584 32984 0 CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState
rlabel metal3 7056 31864 7056 31864 0 CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState
rlabel metal2 10136 31360 10136 31360 0 CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState
rlabel metal2 13272 8960 13272 8960 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2
rlabel metal2 12488 8232 12488 8232 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2
rlabel metal3 10416 8344 10416 8344 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2
rlabel metal2 16744 12040 16744 12040 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2
rlabel metal2 15960 8344 15960 8344 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2
rlabel metal2 22792 8736 22792 8736 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2
rlabel metal2 18872 8792 18872 8792 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2
rlabel metal3 25088 9128 25088 9128 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2
rlabel metal2 21000 30520 21000 30520 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result
rlabel metal2 24584 11088 24584 11088 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2
rlabel metal2 17864 10920 17864 10920 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2
rlabel metal3 17528 9912 17528 9912 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2
rlabel metal2 25704 8736 25704 8736 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock
rlabel metal3 24976 7672 24976 7672 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d
rlabel metal2 24584 7168 24584 7168 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState
rlabel metal2 25424 5096 25424 5096 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d
rlabel metal3 19208 6664 19208 6664 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState
rlabel metal3 18424 7448 18424 7448 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d
rlabel metal2 12152 5600 12152 5600 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState
rlabel metal2 12488 4984 12488 4984 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d
rlabel metal2 15400 5376 15400 5376 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState
rlabel metal3 10080 8008 10080 8008 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d
rlabel metal3 11984 8120 11984 8120 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState
rlabel metal2 11256 7056 11256 7056 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d
rlabel metal2 14056 7672 14056 7672 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState
rlabel metal2 13944 6160 13944 6160 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d
rlabel metal2 16688 5768 16688 5768 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState
rlabel metal2 18088 5880 18088 5880 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d
rlabel metal2 14392 7056 14392 7056 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState
rlabel metal3 21168 8008 21168 8008 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d
rlabel metal2 22792 6720 22792 6720 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState
rlabel metal2 22176 7224 22176 7224 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d
rlabel metal2 22288 7448 22288 7448 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState
rlabel metal2 28840 7784 28840 7784 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState
rlabel metal2 18648 30464 18648 30464 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d
rlabel metal2 20776 31108 20776 31108 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState
rlabel metal2 31864 10192 31864 10192 0 CIRCUIT_2223.tone_generator_2_1.GATES_10.input2
rlabel metal2 37128 12096 37128 12096 0 CIRCUIT_2223.tone_generator_2_1.GATES_11.input2
rlabel metal2 34104 14840 34104 14840 0 CIRCUIT_2223.tone_generator_2_1.GATES_12.input2
rlabel metal3 37072 11480 37072 11480 0 CIRCUIT_2223.tone_generator_2_1.GATES_13.input2
rlabel metal2 36456 11536 36456 11536 0 CIRCUIT_2223.tone_generator_2_1.GATES_14.input2
rlabel metal2 30464 10472 30464 10472 0 CIRCUIT_2223.tone_generator_2_1.GATES_15.input2
rlabel metal2 35784 7728 35784 7728 0 CIRCUIT_2223.tone_generator_2_1.GATES_16.input2
rlabel metal2 31416 8176 31416 8176 0 CIRCUIT_2223.tone_generator_2_1.GATES_17.input2
rlabel metal3 29400 27832 29400 27832 0 CIRCUIT_2223.tone_generator_2_1.GATES_27.result
rlabel metal2 34328 6384 34328 6384 0 CIRCUIT_2223.tone_generator_2_1.GATES_7.input2
rlabel metal3 29176 8904 29176 8904 0 CIRCUIT_2223.tone_generator_2_1.GATES_8.input2
rlabel metal2 32984 7056 32984 7056 0 CIRCUIT_2223.tone_generator_2_1.GATES_9.input2
rlabel metal3 39984 7784 39984 7784 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock
rlabel metal2 41608 4816 41608 4816 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d
rlabel metal2 34776 5768 34776 5768 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState
rlabel metal3 37408 6664 37408 6664 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d
rlabel metal2 37128 5824 37128 5824 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState
rlabel metal2 37576 5768 37576 5768 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d
rlabel metal2 37464 6440 37464 6440 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState
rlabel metal2 35112 4032 35112 4032 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d
rlabel metal2 37800 4704 37800 4704 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState
rlabel metal2 37464 13216 37464 13216 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d
rlabel metal2 38248 12992 38248 12992 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState
rlabel metal2 36344 12264 36344 12264 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d
rlabel metal2 38920 12488 38920 12488 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState
rlabel via2 38360 11368 38360 11368 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d
rlabel metal3 38192 9016 38192 9016 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState
rlabel metal2 41272 10080 41272 10080 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d
rlabel metal2 44072 10080 44072 10080 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState
rlabel metal2 40376 7532 40376 7532 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d
rlabel metal3 42224 8344 42224 8344 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState
rlabel metal2 39368 8512 39368 8512 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d
rlabel metal3 40824 8904 40824 8904 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState
rlabel metal3 38472 7224 38472 7224 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState
rlabel metal3 29848 27720 29848 27720 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d
rlabel metal2 30296 28280 30296 28280 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState
rlabel metal2 31192 18872 31192 18872 0 CIRCUIT_2223.tone_generator_2_2.GATES_10.input2
rlabel metal2 36680 18816 36680 18816 0 CIRCUIT_2223.tone_generator_2_2.GATES_11.input2
rlabel metal3 32536 22456 32536 22456 0 CIRCUIT_2223.tone_generator_2_2.GATES_12.input2
rlabel metal2 36008 20944 36008 20944 0 CIRCUIT_2223.tone_generator_2_2.GATES_13.input2
rlabel metal2 36344 17136 36344 17136 0 CIRCUIT_2223.tone_generator_2_2.GATES_14.input2
rlabel metal2 26992 24024 26992 24024 0 CIRCUIT_2223.tone_generator_2_2.GATES_15.input2
rlabel metal2 32032 24584 32032 24584 0 CIRCUIT_2223.tone_generator_2_2.GATES_16.input2
rlabel metal2 26712 22232 26712 22232 0 CIRCUIT_2223.tone_generator_2_2.GATES_17.input2
rlabel metal3 32032 23352 32032 23352 0 CIRCUIT_2223.tone_generator_2_2.GATES_27.result
rlabel metal2 33152 24024 33152 24024 0 CIRCUIT_2223.tone_generator_2_2.GATES_7.input2
rlabel metal2 26376 21392 26376 21392 0 CIRCUIT_2223.tone_generator_2_2.GATES_8.input2
rlabel metal3 31920 19880 31920 19880 0 CIRCUIT_2223.tone_generator_2_2.GATES_9.input2
rlabel metal2 34216 22960 34216 22960 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock
rlabel metal2 37408 16856 37408 16856 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d
rlabel metal2 38920 17360 38920 17360 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState
rlabel metal2 39928 21700 39928 21700 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d
rlabel metal2 42168 18032 42168 18032 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState
rlabel metal2 41160 17136 41160 17136 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d
rlabel metal2 43960 17136 43960 17136 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState
rlabel metal2 41160 18928 41160 18928 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d
rlabel metal3 43876 19320 43876 19320 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState
rlabel metal3 36008 19992 36008 19992 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d
rlabel metal2 38136 21168 38136 21168 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState
rlabel metal2 38696 21392 38696 21392 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d
rlabel metal2 39144 21616 39144 21616 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState
rlabel metal3 37240 23240 37240 23240 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d
rlabel metal2 40712 23184 40712 23184 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState
rlabel metal2 41272 24584 41272 24584 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d
rlabel metal2 44072 24808 44072 24808 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState
rlabel metal2 35000 26376 35000 26376 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d
rlabel metal3 36008 26152 36008 26152 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState
rlabel metal2 36008 25760 36008 25760 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d
rlabel metal2 35000 24304 35000 24304 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState
rlabel metal2 36344 23632 36344 23632 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState
rlabel metal2 31360 26936 31360 26936 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d
rlabel metal2 30184 28952 30184 28952 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState
rlabel metal2 12712 21336 12712 21336 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2
rlabel metal3 11704 16184 11704 16184 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2
rlabel metal3 10752 15960 10752 15960 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2
rlabel metal2 14840 19768 14840 19768 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2
rlabel metal3 11704 18424 11704 18424 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2
rlabel metal2 14056 21448 14056 21448 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2
rlabel metal2 15400 20552 15400 20552 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2
rlabel metal2 15848 21952 15848 21952 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2
rlabel metal2 19712 29400 19712 29400 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result
rlabel metal2 12544 22232 12544 22232 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2
rlabel metal2 13832 19824 13832 19824 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2
rlabel metal2 14168 19600 14168 19600 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2
rlabel metal2 12712 23520 12712 23520 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock
rlabel metal2 12376 25760 12376 25760 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d
rlabel metal2 9632 26152 9632 26152 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState
rlabel metal2 10752 26264 10752 26264 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d
rlabel metal2 10808 22624 10808 22624 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState
rlabel metal2 11088 21784 11088 21784 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d
rlabel metal2 14168 22288 14168 22288 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState
rlabel metal2 11592 20832 11592 20832 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d
rlabel metal3 9912 20104 9912 20104 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState
rlabel metal2 7224 16632 7224 16632 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d
rlabel metal2 7112 16520 7112 16520 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState
rlabel metal2 9800 18200 9800 18200 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d
rlabel metal2 5208 18088 5208 18088 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState
rlabel metal2 4816 18424 4816 18424 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d
rlabel metal2 2072 19320 2072 19320 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState
rlabel metal2 2632 19936 2632 19936 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d
rlabel metal2 4368 20888 4368 20888 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState
rlabel metal3 6104 21560 6104 21560 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d
rlabel metal2 7224 21896 7224 21896 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState
rlabel metal2 10472 20944 10472 20944 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d
rlabel metal2 13664 22344 13664 22344 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState
rlabel metal2 11704 21952 11704 21952 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState
rlabel metal2 20664 29736 20664 29736 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d
rlabel metal3 22120 30856 22120 30856 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState
rlabel metal2 25872 36456 25872 36456 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock
rlabel metal2 26040 35952 26040 35952 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d
rlabel metal3 26768 34664 26768 34664 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState
rlabel metal2 22904 34888 22904 34888 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock
rlabel metal3 25928 35672 25928 35672 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState
rlabel metal2 24920 35112 24920 35112 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState
rlabel metal2 41048 26992 41048 26992 0 _0000_
rlabel metal2 41048 23800 41048 23800 0 _0001_
rlabel metal2 11032 27888 11032 27888 0 _0002_
rlabel metal2 14504 30968 14504 30968 0 _0003_
rlabel metal2 16184 31836 16184 31836 0 _0004_
rlabel metal2 14392 32760 14392 32760 0 _0005_
rlabel metal2 15960 32928 15960 32928 0 _0006_
rlabel metal2 17752 36064 17752 36064 0 _0007_
rlabel metal2 15624 33992 15624 33992 0 _0008_
rlabel metal2 18984 34104 18984 34104 0 _0009_
rlabel metal2 20216 34496 20216 34496 0 _0010_
rlabel metal2 28504 6888 28504 6888 0 _0011_
rlabel metal2 26936 6272 26936 6272 0 _0012_
rlabel metal2 22904 4704 22904 4704 0 _0013_
rlabel metal2 21112 4144 21112 4144 0 _0014_
rlabel metal2 16520 5320 16520 5320 0 _0015_
rlabel metal2 13832 7112 13832 7112 0 _0016_
rlabel metal2 12264 6272 12264 6272 0 _0017_
rlabel metal2 14840 5488 14840 5488 0 _0018_
rlabel metal2 18200 6160 18200 6160 0 _0019_
rlabel metal2 25256 4704 25256 4704 0 _0020_
rlabel metal2 29176 6272 29176 6272 0 _0021_
rlabel metal3 11256 26936 11256 26936 0 _0022_
rlabel metal3 13552 26488 13552 26488 0 _0023_
rlabel metal2 12824 23520 12824 23520 0 _0024_
rlabel metal2 10696 22008 10696 22008 0 _0025_
rlabel metal2 8344 18144 8344 18144 0 _0026_
rlabel metal2 7672 18032 7672 18032 0 _0027_
rlabel metal2 5656 18816 5656 18816 0 _0028_
rlabel metal2 4816 20552 4816 20552 0 _0029_
rlabel metal2 5096 21896 5096 21896 0 _0030_
rlabel metal2 8680 22736 8680 22736 0 _0031_
rlabel metal2 9912 24360 9912 24360 0 _0032_
rlabel metal3 38080 4872 38080 4872 0 _0033_
rlabel metal2 38192 3416 38192 3416 0 _0034_
rlabel metal2 39816 4704 39816 4704 0 _0035_
rlabel metal2 37576 3976 37576 3976 0 _0036_
rlabel metal2 39928 13944 39928 13944 0 _0037_
rlabel metal2 41160 12544 41160 12544 0 _0038_
rlabel metal2 41832 11704 41832 11704 0 _0039_
rlabel metal2 42952 10416 42952 10416 0 _0040_
rlabel metal2 42616 7476 42616 7476 0 _0041_
rlabel metal2 43064 7840 43064 7840 0 _0042_
rlabel metal2 43624 7112 43624 7112 0 _0043_
rlabel metal3 40376 15512 40376 15512 0 _0044_
rlabel metal2 41888 17080 41888 17080 0 _0045_
rlabel metal2 42952 16688 42952 16688 0 _0046_
rlabel metal2 43456 18648 43456 18648 0 _0047_
rlabel metal3 39592 20104 39592 20104 0 _0048_
rlabel metal3 42224 20552 42224 20552 0 _0049_
rlabel metal2 41944 23688 41944 23688 0 _0050_
rlabel metal2 43064 24304 43064 24304 0 _0051_
rlabel metal2 37576 26656 37576 26656 0 _0052_
rlabel metal2 38920 26600 38920 26600 0 _0053_
rlabel metal2 37240 24360 37240 24360 0 _0054_
rlabel metal2 26040 27272 26040 27272 0 _0055_
rlabel metal2 28056 28224 28056 28224 0 _0056_
rlabel metal2 28672 29176 28672 29176 0 _0057_
rlabel metal3 27160 29960 27160 29960 0 _0058_
rlabel metal3 23128 24472 23128 24472 0 _0059_
rlabel metal2 16072 24528 16072 24528 0 _0060_
rlabel metal2 21336 25088 21336 25088 0 _0061_
rlabel metal2 22568 26040 22568 26040 0 _0062_
rlabel metal2 21448 27608 21448 27608 0 _0063_
rlabel metal2 18536 28504 18536 28504 0 _0064_
rlabel metal2 16464 29624 16464 29624 0 _0065_
rlabel metal3 15624 27944 15624 27944 0 _0066_
rlabel metal3 18648 26936 18648 26936 0 _0067_
rlabel metal2 41832 39984 41832 39984 0 _0068_
rlabel metal3 36848 30072 36848 30072 0 _0069_
rlabel metal2 41608 30184 41608 30184 0 _0070_
rlabel metal2 41720 29736 41720 29736 0 _0071_
rlabel metal2 43064 31696 43064 31696 0 _0072_
rlabel metal2 40152 39368 40152 39368 0 _0073_
rlabel metal2 41608 39144 41608 39144 0 _0074_
rlabel metal2 39368 40824 39368 40824 0 _0075_
rlabel metal2 43232 38248 43232 38248 0 _0076_
rlabel metal2 43512 35336 43512 35336 0 _0077_
rlabel metal2 38360 36848 38360 36848 0 _0078_
rlabel metal2 41944 29512 41944 29512 0 _0079_
rlabel metal2 18200 19712 18200 19712 0 _0080_
rlabel metal2 15736 18872 15736 18872 0 _0081_
rlabel metal2 14952 18032 14952 18032 0 _0082_
rlabel metal2 38360 39928 38360 39928 0 _0083_
rlabel metal2 38248 40824 38248 40824 0 _0084_
rlabel metal2 31080 35672 31080 35672 0 _0085_
rlabel metal3 32984 33992 32984 33992 0 _0086_
rlabel metal3 32760 35000 32760 35000 0 _0087_
rlabel metal2 35504 29512 35504 29512 0 _0088_
rlabel metal2 33544 31892 33544 31892 0 _0089_
rlabel metal2 32424 32984 32424 32984 0 _0090_
rlabel metal2 33208 38808 33208 38808 0 _0091_
rlabel metal2 33768 38052 33768 38052 0 _0092_
rlabel metal2 36568 40544 36568 40544 0 _0093_
rlabel metal2 32536 40824 32536 40824 0 _0094_
rlabel metal3 28392 39704 28392 39704 0 _0095_
rlabel metal2 27608 39984 27608 39984 0 _0096_
rlabel metal3 28616 38136 28616 38136 0 _0097_
rlabel metal2 33152 28728 33152 28728 0 _0098_
rlabel metal2 20608 9128 20608 9128 0 _0099_
rlabel metal2 21448 9968 21448 9968 0 _0100_
rlabel metal2 23464 9968 23464 9968 0 _0101_
rlabel metal2 23632 10808 23632 10808 0 _0102_
rlabel metal2 10136 10024 10136 10024 0 _0103_
rlabel metal2 11704 9688 11704 9688 0 _0104_
rlabel metal2 14728 12488 14728 12488 0 _0105_
rlabel metal2 14280 9968 14280 9968 0 _0106_
rlabel metal2 23128 14168 23128 14168 0 _0107_
rlabel metal2 20776 15344 20776 15344 0 _0108_
rlabel metal2 21784 16352 21784 16352 0 _0109_
rlabel metal2 24696 17920 24696 17920 0 _0110_
rlabel metal2 25872 20552 25872 20552 0 _0111_
rlabel metal2 29288 20160 29288 20160 0 _0112_
rlabel metal2 29960 19768 29960 19768 0 _0113_
rlabel metal3 11816 15176 11816 15176 0 _0114_
rlabel metal2 9800 14728 9800 14728 0 _0115_
rlabel metal2 15064 16128 15064 16128 0 _0116_
rlabel metal2 10696 16800 10696 16800 0 _0117_
rlabel metal3 20160 20104 20160 20104 0 _0118_
rlabel metal2 17528 21168 17528 21168 0 _0119_
rlabel metal2 17472 21784 17472 21784 0 _0120_
rlabel metal2 20776 21056 20776 21056 0 _0121_
rlabel metal2 15792 13048 15792 13048 0 _0122_
rlabel metal2 18256 11480 18256 11480 0 _0123_
rlabel metal3 12096 12824 12096 12824 0 _0124_
rlabel metal2 34328 13328 34328 13328 0 _0125_
rlabel metal2 32032 15512 32032 15512 0 _0126_
rlabel metal3 33376 11480 33376 11480 0 _0127_
rlabel metal3 33152 12040 33152 12040 0 _0128_
rlabel metal2 28392 11480 28392 11480 0 _0129_
rlabel metal2 33208 7896 33208 7896 0 _0130_
rlabel metal2 29848 7784 29848 7784 0 _0131_
rlabel metal2 33208 6328 33208 6328 0 _0132_
rlabel metal2 27720 9576 27720 9576 0 _0133_
rlabel metal2 30912 6776 30912 6776 0 _0134_
rlabel metal2 29960 10192 29960 10192 0 _0135_
rlabel metal3 34720 17528 34720 17528 0 _0136_
rlabel metal2 30968 22008 30968 22008 0 _0137_
rlabel metal2 33992 19376 33992 19376 0 _0138_
rlabel metal2 34328 16968 34328 16968 0 _0139_
rlabel metal2 24808 24416 24808 24416 0 _0140_
rlabel metal2 29288 24304 29288 24304 0 _0141_
rlabel metal2 25816 22624 25816 22624 0 _0142_
rlabel metal2 30856 23576 30856 23576 0 _0143_
rlabel metal2 24808 27496 24808 27496 0 _0144_
rlabel metal2 24920 28056 24920 28056 0 _0145_
rlabel metal2 24248 31472 24248 31472 0 _0146_
rlabel metal2 24360 29904 24360 29904 0 _0147_
rlabel metal2 27944 29456 27944 29456 0 _0148_
rlabel metal3 26880 31640 26880 31640 0 _0149_
rlabel metal2 22904 16912 22904 16912 0 _0150_
rlabel metal2 23128 16520 23128 16520 0 _0151_
rlabel metal2 26824 20888 26824 20888 0 _0152_
rlabel metal3 26152 14336 26152 14336 0 _0153_
rlabel metal2 26712 17192 26712 17192 0 _0154_
rlabel metal2 27384 27440 27384 27440 0 _0155_
rlabel metal3 25872 29400 25872 29400 0 _0156_
rlabel metal2 35504 13720 35504 13720 0 _0157_
rlabel metal2 26264 29624 26264 29624 0 _0158_
rlabel metal2 26152 30856 26152 30856 0 _0159_
rlabel metal3 24976 29624 24976 29624 0 _0160_
rlabel metal2 18480 17080 18480 17080 0 _0161_
rlabel metal2 27496 27832 27496 27832 0 _0162_
rlabel metal3 25536 27832 25536 27832 0 _0163_
rlabel metal2 34664 14756 34664 14756 0 _0164_
rlabel metal2 24360 15680 24360 15680 0 _0165_
rlabel metal2 25704 27832 25704 27832 0 _0166_
rlabel metal3 24640 16072 24640 16072 0 _0167_
rlabel metal2 27216 13944 27216 13944 0 _0168_
rlabel metal2 25704 16072 25704 16072 0 _0169_
rlabel metal2 28616 14392 28616 14392 0 _0170_
rlabel metal2 25816 19264 25816 19264 0 _0171_
rlabel metal2 28112 14504 28112 14504 0 _0172_
rlabel metal2 28168 19208 28168 19208 0 _0173_
rlabel metal2 29288 14616 29288 14616 0 _0174_
rlabel metal2 9464 34104 9464 34104 0 _0175_
rlabel metal2 8008 33376 8008 33376 0 _0176_
rlabel metal2 9128 30968 9128 30968 0 _0177_
rlabel metal2 17528 8624 17528 8624 0 _0178_
rlabel metal2 17080 8176 17080 8176 0 _0179_
rlabel metal2 17976 7952 17976 7952 0 _0180_
rlabel metal2 21560 9632 21560 9632 0 _0181_
rlabel metal2 21448 8288 21448 8288 0 _0182_
rlabel metal3 22344 8792 22344 8792 0 _0183_
rlabel metal2 18648 10024 18648 10024 0 _0184_
rlabel metal3 19544 8344 19544 8344 0 _0185_
rlabel metal2 19712 7672 19712 7672 0 _0186_
rlabel metal2 18536 8680 18536 8680 0 _0187_
rlabel metal2 18480 7448 18480 7448 0 _0188_
rlabel metal3 13160 8680 13160 8680 0 _0189_
rlabel metal2 23072 9240 23072 9240 0 _0190_
rlabel metal2 23800 9632 23800 9632 0 _0191_
rlabel metal2 22568 8512 22568 8512 0 _0192_
rlabel metal3 12880 8232 12880 8232 0 _0193_
rlabel metal2 14168 8316 14168 8316 0 _0194_
rlabel metal2 14056 8736 14056 8736 0 _0195_
rlabel metal2 12824 9128 12824 9128 0 _0196_
rlabel metal3 14224 9016 14224 9016 0 _0197_
rlabel metal2 18984 8176 18984 8176 0 _0198_
rlabel metal2 19208 9744 19208 9744 0 _0199_
rlabel metal3 13216 20664 13216 20664 0 _0200_
rlabel metal2 12936 22120 12936 22120 0 _0201_
rlabel metal2 13720 21224 13720 21224 0 _0202_
rlabel metal2 13720 21952 13720 21952 0 _0203_
rlabel metal3 13216 21112 13216 21112 0 _0204_
rlabel metal2 14728 21616 14728 21616 0 _0205_
rlabel metal2 14784 20440 14784 20440 0 _0206_
rlabel metal3 13384 21448 13384 21448 0 _0207_
rlabel metal2 12208 19320 12208 19320 0 _0208_
rlabel metal3 13328 19992 13328 19992 0 _0209_
rlabel metal3 13328 20104 13328 20104 0 _0210_
rlabel metal2 11144 15680 11144 15680 0 _0211_
rlabel metal3 9128 15848 9128 15848 0 _0212_
rlabel metal2 10472 16408 10472 16408 0 _0213_
rlabel metal2 11872 21000 11872 21000 0 _0214_
rlabel metal3 11256 18312 11256 18312 0 _0215_
rlabel metal2 13832 17976 13832 17976 0 _0216_
rlabel metal2 12096 17752 12096 17752 0 _0217_
rlabel metal2 14168 20468 14168 20468 0 _0218_
rlabel metal2 14616 21840 14616 21840 0 _0219_
rlabel metal3 34608 7672 34608 7672 0 _0220_
rlabel metal2 34216 9744 34216 9744 0 _0221_
rlabel metal2 36568 9912 36568 9912 0 _0222_
rlabel metal2 38360 10248 38360 10248 0 _0223_
rlabel metal3 35616 11592 35616 11592 0 _0224_
rlabel metal2 38640 9240 38640 9240 0 _0225_
rlabel metal2 35448 9800 35448 9800 0 _0226_
rlabel metal2 34888 10696 34888 10696 0 _0227_
rlabel metal3 31416 10696 31416 10696 0 _0228_
rlabel metal2 35224 10920 35224 10920 0 _0229_
rlabel metal2 35448 7840 35448 7840 0 _0230_
rlabel metal2 34104 7840 34104 7840 0 _0231_
rlabel metal2 34888 7672 34888 7672 0 _0232_
rlabel metal2 35896 10136 35896 10136 0 _0233_
rlabel metal3 36400 8792 36400 8792 0 _0234_
rlabel metal3 36176 9240 36176 9240 0 _0235_
rlabel metal3 35784 13160 35784 13160 0 _0236_
rlabel metal2 37464 10192 37464 10192 0 _0237_
rlabel metal2 37688 10248 37688 10248 0 _0238_
rlabel metal3 37072 9800 37072 9800 0 _0239_
rlabel metal3 36120 12040 36120 12040 0 _0240_
rlabel metal2 32312 24192 32312 24192 0 _0241_
rlabel metal2 35448 23352 35448 23352 0 _0242_
rlabel metal2 35000 22792 35000 22792 0 _0243_
rlabel metal2 35056 22344 35056 22344 0 _0244_
rlabel metal3 36736 21000 36736 21000 0 _0245_
rlabel metal2 34720 21560 34720 21560 0 _0246_
rlabel metal2 34440 21728 34440 21728 0 _0247_
rlabel metal2 37128 20384 37128 20384 0 _0248_
rlabel metal2 35224 20048 35224 20048 0 _0249_
rlabel metal3 35672 20888 35672 20888 0 _0250_
rlabel metal2 33432 23464 33432 23464 0 _0251_
rlabel metal2 32536 20384 32536 20384 0 _0252_
rlabel metal2 33992 21224 33992 21224 0 _0253_
rlabel metal3 34776 22344 34776 22344 0 _0254_
rlabel metal2 35000 21784 35000 21784 0 _0255_
rlabel metal2 35280 20888 35280 20888 0 _0256_
rlabel metal2 36568 18648 36568 18648 0 _0257_
rlabel metal2 35448 21616 35448 21616 0 _0258_
rlabel metal2 35560 20776 35560 20776 0 _0259_
rlabel metal2 36120 22064 36120 22064 0 _0260_
rlabel metal2 31864 22568 31864 22568 0 _0261_
rlabel metal3 39928 31304 39928 31304 0 _0262_
rlabel metal3 39200 31864 39200 31864 0 _0263_
rlabel metal2 38808 31416 38808 31416 0 _0264_
rlabel metal3 39760 31528 39760 31528 0 _0265_
rlabel metal2 42504 35952 42504 35952 0 _0266_
rlabel metal2 37240 30856 37240 30856 0 _0267_
rlabel metal2 39704 32984 39704 32984 0 _0268_
rlabel metal2 31472 30744 31472 30744 0 _0269_
rlabel metal2 37688 35784 37688 35784 0 _0270_
rlabel metal2 37576 31024 37576 31024 0 _0271_
rlabel metal3 40712 32312 40712 32312 0 _0272_
rlabel metal2 40432 31192 40432 31192 0 _0273_
rlabel metal3 41944 30184 41944 30184 0 _0274_
rlabel metal2 42504 32312 42504 32312 0 _0275_
rlabel metal2 40824 35336 40824 35336 0 _0276_
rlabel metal2 41384 39032 41384 39032 0 _0277_
rlabel metal2 41216 38024 41216 38024 0 _0278_
rlabel metal2 44016 38024 44016 38024 0 _0279_
rlabel metal2 40600 38864 40600 38864 0 _0280_
rlabel metal2 43736 40376 43736 40376 0 _0281_
rlabel metal3 41776 37912 41776 37912 0 _0282_
rlabel metal2 43288 35168 43288 35168 0 _0283_
rlabel metal2 43176 34888 43176 34888 0 _0284_
rlabel metal3 38864 37240 38864 37240 0 _0285_
rlabel metal2 39816 36960 39816 36960 0 _0286_
rlabel metal2 37352 34552 37352 34552 0 _0287_
rlabel metal2 38808 36232 38808 36232 0 _0288_
rlabel metal2 38304 35112 38304 35112 0 _0289_
rlabel metal3 33376 29624 33376 29624 0 _0290_
rlabel metal2 35112 30408 35112 30408 0 _0291_
rlabel metal2 36792 37408 36792 37408 0 _0292_
rlabel metal2 38920 32592 38920 32592 0 _0293_
rlabel metal2 39368 33600 39368 33600 0 _0294_
rlabel metal2 18592 19768 18592 19768 0 _0295_
rlabel metal2 19656 15232 19656 15232 0 _0296_
rlabel metal2 20944 17640 20944 17640 0 _0297_
rlabel metal3 19656 18424 19656 18424 0 _0298_
rlabel metal3 17976 19992 17976 19992 0 _0299_
rlabel metal3 16632 18536 16632 18536 0 _0300_
rlabel metal3 16800 18424 16800 18424 0 _0301_
rlabel metal2 31192 11760 31192 11760 0 _0302_
rlabel metal2 14504 18144 14504 18144 0 _0303_
rlabel metal2 39648 38696 39648 38696 0 _0304_
rlabel metal2 38080 34664 38080 34664 0 _0305_
rlabel metal2 37464 36568 37464 36568 0 _0306_
rlabel metal2 30800 38024 30800 38024 0 _0307_
rlabel metal2 38584 39088 38584 39088 0 _0308_
rlabel metal2 27384 33824 27384 33824 0 _0309_
rlabel metal3 26992 32424 26992 32424 0 _0310_
rlabel metal2 28056 33208 28056 33208 0 _0311_
rlabel metal2 30968 34496 30968 34496 0 _0312_
rlabel metal2 37128 35112 37128 35112 0 _0313_
rlabel metal2 25592 34328 25592 34328 0 _0314_
rlabel metal3 26544 34104 26544 34104 0 _0315_
rlabel metal3 30464 34104 30464 34104 0 _0316_
rlabel metal2 35616 34888 35616 34888 0 _0317_
rlabel metal2 32536 34888 32536 34888 0 _0318_
rlabel metal2 29176 35280 29176 35280 0 _0319_
rlabel metal2 26712 32592 26712 32592 0 _0320_
rlabel metal2 24696 33040 24696 33040 0 _0321_
rlabel metal3 26544 35560 26544 35560 0 _0322_
rlabel metal2 29512 33264 29512 33264 0 _0323_
rlabel metal2 27272 35616 27272 35616 0 _0324_
rlabel metal2 27048 35952 27048 35952 0 _0325_
rlabel metal3 29064 34776 29064 34776 0 _0326_
rlabel metal2 30408 35000 30408 35000 0 _0327_
rlabel metal2 35448 34944 35448 34944 0 _0328_
rlabel metal2 36456 32872 36456 32872 0 _0329_
rlabel metal2 29400 35000 29400 35000 0 _0330_
rlabel metal2 29736 35224 29736 35224 0 _0331_
rlabel metal2 29904 33320 29904 33320 0 _0332_
rlabel metal2 28952 32816 28952 32816 0 _0333_
rlabel metal2 35672 32872 35672 32872 0 _0334_
rlabel metal3 36400 32648 36400 32648 0 _0335_
rlabel metal2 36344 32480 36344 32480 0 _0336_
rlabel metal2 35000 31080 35000 31080 0 _0337_
rlabel metal2 31752 29904 31752 29904 0 _0338_
rlabel metal2 30688 29624 30688 29624 0 _0339_
rlabel metal2 31304 30688 31304 30688 0 _0340_
rlabel metal2 29400 33656 29400 33656 0 _0341_
rlabel metal3 30408 31864 30408 31864 0 _0342_
rlabel metal2 33208 32256 33208 32256 0 _0343_
rlabel metal2 33880 32872 33880 32872 0 _0344_
rlabel metal2 31864 31472 31864 31472 0 _0345_
rlabel metal2 32536 33152 32536 33152 0 _0346_
rlabel metal3 33712 38024 33712 38024 0 _0347_
rlabel metal2 33656 37632 33656 37632 0 _0348_
rlabel metal2 36120 39984 36120 39984 0 _0349_
rlabel metal2 34888 40264 34888 40264 0 _0350_
rlabel metal2 37016 39816 37016 39816 0 _0351_
rlabel metal4 36344 40544 36344 40544 0 _0352_
rlabel metal2 32480 38808 32480 38808 0 _0353_
rlabel metal2 27048 31304 27048 31304 0 _0354_
rlabel metal2 30072 38248 30072 38248 0 _0355_
rlabel metal3 31976 38696 31976 38696 0 _0356_
rlabel metal2 31976 39704 31976 39704 0 _0357_
rlabel metal2 30072 39984 30072 39984 0 _0358_
rlabel metal2 30240 38136 30240 38136 0 _0359_
rlabel metal2 27776 39368 27776 39368 0 _0360_
rlabel metal2 27720 40040 27720 40040 0 _0361_
rlabel metal3 30128 38920 30128 38920 0 _0362_
rlabel metal2 27496 30128 27496 30128 0 _0363_
rlabel metal2 30352 37240 30352 37240 0 _0364_
rlabel metal2 31304 29792 31304 29792 0 _0365_
rlabel metal3 31780 5992 31780 5992 0 _0366_
rlabel metal2 8344 25928 8344 25928 0 _0367_
rlabel metal3 16856 32648 16856 32648 0 _0368_
rlabel metal3 21000 28616 21000 28616 0 _0369_
rlabel metal3 15680 31864 15680 31864 0 _0370_
rlabel metal2 18312 35280 18312 35280 0 _0371_
rlabel metal2 20552 34048 20552 34048 0 _0372_
rlabel metal3 27832 14448 27832 14448 0 _0373_
rlabel metal2 21784 12880 21784 12880 0 _0374_
rlabel metal3 21840 10696 21840 10696 0 _0375_
rlabel metal2 30296 13104 30296 13104 0 _0376_
rlabel metal2 21728 11592 21728 11592 0 _0377_
rlabel metal2 21672 10920 21672 10920 0 _0378_
rlabel metal2 18872 22176 18872 22176 0 _0379_
rlabel metal2 21952 9800 21952 9800 0 _0380_
rlabel metal2 18984 20832 18984 20832 0 _0381_
rlabel metal2 22792 10864 22792 10864 0 _0382_
rlabel metal2 31528 13272 31528 13272 0 _0383_
rlabel metal2 24024 10864 24024 10864 0 _0384_
rlabel metal2 18984 13776 18984 13776 0 _0385_
rlabel metal2 13160 10864 13160 10864 0 _0386_
rlabel metal3 13328 10696 13328 10696 0 _0387_
rlabel metal2 11704 10864 11704 10864 0 _0388_
rlabel metal2 30240 8008 30240 8008 0 _0389_
rlabel metal2 12600 10192 12600 10192 0 _0390_
rlabel metal2 14392 13216 14392 13216 0 _0391_
rlabel metal2 14784 10584 14784 10584 0 _0392_
rlabel metal2 26488 14224 26488 14224 0 _0393_
rlabel metal2 26432 15624 26432 15624 0 _0394_
rlabel metal2 23184 15064 23184 15064 0 _0395_
rlabel metal2 21560 17696 21560 17696 0 _0396_
rlabel metal3 21000 16072 21000 16072 0 _0397_
rlabel metal2 21896 17696 21896 17696 0 _0398_
rlabel metal2 21336 16128 21336 16128 0 _0399_
rlabel metal2 25368 17752 25368 17752 0 _0400_
rlabel metal2 30632 5152 30632 5152 0 _0401_
rlabel metal3 30240 4200 30240 4200 0 _0402_
rlabel metal3 24024 16800 24024 16800 0 _0403_
rlabel metal2 23856 16632 23856 16632 0 _0404_
rlabel metal2 18760 14000 18760 14000 0 _0405_
rlabel metal4 18872 10192 18872 10192 0 _0406_
rlabel metal2 29512 5544 29512 5544 0 _0407_
rlabel metal2 28168 4704 28168 4704 0 _0408_
rlabel metal2 28728 4984 28728 4984 0 _0409_
rlabel metal2 27272 5488 27272 5488 0 _0410_
rlabel metal2 14952 5152 14952 5152 0 _0411_
rlabel metal2 23128 3808 23128 3808 0 _0412_
rlabel metal2 21336 3808 21336 3808 0 _0413_
rlabel metal3 13440 5208 13440 5208 0 _0414_
rlabel metal2 16688 4312 16688 4312 0 _0415_
rlabel metal2 14168 5936 14168 5936 0 _0416_
rlabel metal3 13384 3528 13384 3528 0 _0417_
rlabel metal2 12376 5600 12376 5600 0 _0418_
rlabel metal2 14504 5152 14504 5152 0 _0419_
rlabel metal2 18424 5152 18424 5152 0 _0420_
rlabel metal3 25088 4312 25088 4312 0 _0421_
rlabel metal2 31080 5152 31080 5152 0 _0422_
rlabel metal2 29400 5600 29400 5600 0 _0423_
rlabel metal2 26152 17920 26152 17920 0 _0424_
rlabel metal2 26264 16800 26264 16800 0 _0425_
rlabel metal3 14392 15512 14392 15512 0 _0426_
rlabel metal2 20496 17416 20496 17416 0 _0427_
rlabel metal2 6552 23016 6552 23016 0 _0428_
rlabel metal2 7784 24304 7784 24304 0 _0429_
rlabel metal2 8736 24584 8736 24584 0 _0430_
rlabel metal2 12488 27384 12488 27384 0 _0431_
rlabel metal2 14168 26320 14168 26320 0 _0432_
rlabel metal2 12488 25088 12488 25088 0 _0433_
rlabel metal2 7224 24360 7224 24360 0 _0434_
rlabel metal2 10920 22680 10920 22680 0 _0435_
rlabel metal2 5992 21616 5992 21616 0 _0436_
rlabel metal3 7896 18424 7896 18424 0 _0437_
rlabel metal2 7896 18760 7896 18760 0 _0438_
rlabel metal3 5544 19208 5544 19208 0 _0439_
rlabel metal2 6104 21952 6104 21952 0 _0440_
rlabel metal2 5376 20664 5376 20664 0 _0441_
rlabel metal3 5208 22344 5208 22344 0 _0442_
rlabel metal2 8120 23128 8120 23128 0 _0443_
rlabel metal3 8736 23800 8736 23800 0 _0444_
rlabel metal2 27832 21336 27832 21336 0 _0445_
rlabel metal2 27608 19712 27608 19712 0 _0446_
rlabel metal2 25704 20776 25704 20776 0 _0447_
rlabel metal2 29960 20776 29960 20776 0 _0448_
rlabel metal2 28392 19992 28392 19992 0 _0449_
rlabel metal2 29624 18480 29624 18480 0 _0450_
rlabel metal2 12264 14952 12264 14952 0 _0451_
rlabel metal2 12600 14896 12600 14896 0 _0452_
rlabel metal2 13608 15008 13608 15008 0 _0453_
rlabel metal2 15512 15624 15512 15624 0 _0454_
rlabel metal2 12824 16352 12824 16352 0 _0455_
rlabel metal2 22120 21448 22120 21448 0 _0456_
rlabel metal2 21560 21280 21560 21280 0 _0457_
rlabel metal2 17136 21560 17136 21560 0 _0458_
rlabel metal3 17584 21560 17584 21560 0 _0459_
rlabel metal2 19208 20944 19208 20944 0 _0460_
rlabel metal2 20552 20832 20552 20832 0 _0461_
rlabel metal3 28560 14616 28560 14616 0 _0462_
rlabel metal2 30520 14728 30520 14728 0 _0463_
rlabel metal2 42728 14112 42728 14112 0 _0464_
rlabel metal2 42168 6552 42168 6552 0 _0465_
rlabel metal2 38584 5880 38584 5880 0 _0466_
rlabel metal2 42448 5096 42448 5096 0 _0467_
rlabel metal2 38584 4592 38584 4592 0 _0468_
rlabel metal2 39480 5488 39480 5488 0 _0469_
rlabel metal2 37968 3528 37968 3528 0 _0470_
rlabel metal2 43120 20776 43120 20776 0 _0471_
rlabel metal3 41664 14504 41664 14504 0 _0472_
rlabel metal2 41832 14056 41832 14056 0 _0473_
rlabel metal3 40824 13720 40824 13720 0 _0474_
rlabel metal2 41552 12264 41552 12264 0 _0475_
rlabel metal2 43512 12488 43512 12488 0 _0476_
rlabel metal2 42616 11648 42616 11648 0 _0477_
rlabel metal2 42280 6664 42280 6664 0 _0478_
rlabel metal2 42728 8736 42728 8736 0 _0479_
rlabel metal2 43288 7392 43288 7392 0 _0480_
rlabel metal2 43960 6272 43960 6272 0 _0481_
rlabel metal2 18088 13272 18088 13272 0 _0482_
rlabel metal3 17136 12376 17136 12376 0 _0483_
rlabel metal2 19096 12992 19096 12992 0 _0484_
rlabel metal2 12824 13608 12824 13608 0 _0485_
rlabel metal2 31864 13888 31864 13888 0 _0486_
rlabel metal2 34216 14112 34216 14112 0 _0487_
rlabel metal2 34776 14224 34776 14224 0 _0488_
rlabel metal2 32424 15792 32424 15792 0 _0489_
rlabel metal2 33208 13216 33208 13216 0 _0490_
rlabel metal2 32088 12488 32088 12488 0 _0491_
rlabel metal2 29176 12320 29176 12320 0 _0492_
rlabel metal3 28280 12152 28280 12152 0 _0493_
rlabel metal2 33096 6776 33096 6776 0 _0494_
rlabel metal3 33096 7560 33096 7560 0 _0495_
rlabel metal2 30128 8792 30128 8792 0 _0496_
rlabel metal2 33544 7112 33544 7112 0 _0497_
rlabel metal2 24024 22792 24024 22792 0 _0498_
rlabel metal2 38920 23296 38920 23296 0 _0499_
rlabel metal2 38808 25368 38808 25368 0 _0500_
rlabel metal2 42056 15624 42056 15624 0 _0501_
rlabel metal2 41160 15344 41160 15344 0 _0502_
rlabel metal2 41944 15960 41944 15960 0 _0503_
rlabel metal2 42392 20944 42392 20944 0 _0504_
rlabel metal2 42616 18144 42616 18144 0 _0505_
rlabel metal2 42896 18424 42896 18424 0 _0506_
rlabel metal2 41720 23800 41720 23800 0 _0507_
rlabel metal3 40656 20104 40656 20104 0 _0508_
rlabel metal2 43512 21056 43512 21056 0 _0509_
rlabel metal2 39480 25872 39480 25872 0 _0510_
rlabel metal2 42280 24976 42280 24976 0 _0511_
rlabel metal2 42728 23968 42728 23968 0 _0512_
rlabel metal2 38584 26320 38584 26320 0 _0513_
rlabel metal2 39256 26488 39256 26488 0 _0514_
rlabel metal2 37576 24808 37576 24808 0 _0515_
rlabel metal2 28056 12768 28056 12768 0 _0516_
rlabel metal3 26992 11256 26992 11256 0 _0517_
rlabel metal2 30688 8008 30688 8008 0 _0518_
rlabel metal2 30968 8232 30968 8232 0 _0519_
rlabel metal2 31304 10864 31304 10864 0 _0520_
rlabel metal3 30576 18424 30576 18424 0 _0521_
rlabel metal2 33432 18424 33432 18424 0 _0522_
rlabel metal2 34328 16520 34328 16520 0 _0523_
rlabel metal2 31528 21280 31528 21280 0 _0524_
rlabel metal2 32872 19712 32872 19712 0 _0525_
rlabel metal2 34104 18368 34104 18368 0 _0526_
rlabel metal2 27160 23520 27160 23520 0 _0527_
rlabel metal2 25872 24696 25872 24696 0 _0528_
rlabel metal3 29064 22232 29064 22232 0 _0529_
rlabel metal2 29624 23184 29624 23184 0 _0530_
rlabel metal2 25592 22176 25592 22176 0 _0531_
rlabel metal2 31192 23016 31192 23016 0 _0532_
rlabel metal3 27160 28056 27160 28056 0 _0533_
rlabel metal3 27160 27944 27160 27944 0 _0534_
rlabel metal2 20384 28392 20384 28392 0 _0535_
rlabel metal3 16912 29512 16912 29512 0 _0536_
rlabel metal2 44184 3080 44184 3080 0 clk
rlabel metal2 44184 9352 44184 9352 0 io_in[0]
rlabel metal3 44730 12824 44730 12824 0 io_in[1]
rlabel metal3 45304 16688 45304 16688 0 io_in[2]
rlabel metal3 44786 19544 44786 19544 0 io_in[3]
rlabel metal2 44184 23016 44184 23016 0 io_in[4]
rlabel metal2 44632 26992 44632 26992 0 io_in[5]
rlabel metal3 45304 30016 45304 30016 0 io_out[0]
rlabel metal3 44478 32984 44478 32984 0 io_out[1]
rlabel metal3 45304 36736 45304 36736 0 io_out[2]
rlabel metal2 43176 39368 43176 39368 0 io_out[3]
rlabel metal2 41944 42448 41944 42448 0 io_out[4]
rlabel metal2 43848 4592 43848 4592 0 net1
rlabel metal2 44072 34160 44072 34160 0 net10
rlabel metal2 40824 36904 40824 36904 0 net11
rlabel metal2 44184 27328 44184 27328 0 net12
rlabel metal2 44184 26656 44184 26656 0 net13
rlabel metal2 26488 36120 26488 36120 0 net14
rlabel metal2 20216 31136 20216 31136 0 net15
rlabel metal2 10472 36120 10472 36120 0 net16
rlabel metal2 7224 31836 7224 31836 0 net17
rlabel metal2 10920 32872 10920 32872 0 net18
rlabel metal2 8904 29008 8904 29008 0 net19
rlabel metal2 27496 11984 27496 11984 0 net2
rlabel metal3 13104 34104 13104 34104 0 net20
rlabel metal2 15848 35728 15848 35728 0 net21
rlabel metal2 16744 35728 16744 35728 0 net22
rlabel metal2 18872 35000 18872 35000 0 net23
rlabel metal2 19432 31920 19432 31920 0 net24
rlabel metal2 8904 6384 8904 6384 0 net25
rlabel metal2 9128 14112 9128 14112 0 net26
rlabel metal2 14056 17248 14056 17248 0 net27
rlabel metal3 14504 15960 14504 15960 0 net28
rlabel metal2 19432 16632 19432 16632 0 net29
rlabel metal2 28616 12656 28616 12656 0 net3
rlabel metal2 19432 15736 19432 15736 0 net30
rlabel metal2 10584 16520 10584 16520 0 net31
rlabel metal2 18200 20720 18200 20720 0 net32
rlabel metal2 20440 21280 20440 21280 0 net33
rlabel metal2 20552 22232 20552 22232 0 net34
rlabel metal2 21728 23128 21728 23128 0 net35
rlabel metal2 26936 9352 26936 9352 0 net36
rlabel metal2 29176 7056 29176 7056 0 net37
rlabel metal2 32256 7224 32256 7224 0 net38
rlabel metal2 30632 14448 30632 14448 0 net39
rlabel metal2 44184 24528 44184 24528 0 net4
rlabel metal2 32648 11312 32648 11312 0 net40
rlabel metal2 24528 18424 24528 18424 0 net41
rlabel metal2 23576 29848 23576 29848 0 net42
rlabel metal2 24416 28392 24416 28392 0 net43
rlabel metal2 24808 29176 24808 29176 0 net44
rlabel metal2 33376 20552 33376 20552 0 net45
rlabel metal2 29736 29568 29736 29568 0 net46
rlabel metal2 32928 30184 32928 30184 0 net47
rlabel metal2 29960 30520 29960 30520 0 net48
rlabel metal2 29624 29400 29624 29400 0 net49
rlabel metal3 43764 20104 43764 20104 0 net5
rlabel metal2 31640 34104 31640 34104 0 net50
rlabel metal2 32592 39592 32592 39592 0 net51
rlabel metal2 31640 41160 31640 41160 0 net52
rlabel metal2 31864 29624 31864 29624 0 net53
rlabel metal2 35784 30184 35784 30184 0 net54
rlabel metal2 41048 29792 41048 29792 0 net55
rlabel metal2 40936 40544 40936 40544 0 net56
rlabel metal2 41272 39312 41272 39312 0 net57
rlabel metal2 43848 36064 43848 36064 0 net58
rlabel metal2 38808 38024 38808 38024 0 net59
rlabel metal2 43792 23240 43792 23240 0 net6
rlabel metal2 40264 30016 40264 30016 0 net60
rlabel metal2 32368 33544 32368 33544 0 net61
rlabel metal2 43848 26992 43848 26992 0 net7
rlabel metal2 43848 6384 43848 6384 0 net8
rlabel metal2 44072 30240 44072 30240 0 net9
rlabel metal2 44184 6048 44184 6048 0 rst_n
rlabel metal2 35112 38332 35112 38332 0 slow_clock\[0\]
rlabel metal2 34440 38388 34440 38388 0 slow_clock\[1\]
rlabel metal2 35616 41160 35616 41160 0 slow_clock\[2\]
rlabel metal2 34664 41216 34664 41216 0 slow_clock\[3\]
rlabel metal2 30352 37912 30352 37912 0 slow_clock\[4\]
rlabel metal2 29736 40320 29736 40320 0 slow_clock\[5\]
rlabel metal2 29960 38052 29960 38052 0 slow_clock\[6\]
rlabel metal3 40432 34216 40432 34216 0 spi_dac_i_2.counter\[0\]
rlabel via2 37016 30856 37016 30856 0 spi_dac_i_2.counter\[1\]
rlabel metal3 40264 31080 40264 31080 0 spi_dac_i_2.counter\[2\]
rlabel metal2 43512 29736 43512 29736 0 spi_dac_i_2.counter\[3\]
rlabel metal3 41384 30856 41384 30856 0 spi_dac_i_2.counter\[4\]
rlabel metal3 40152 39032 40152 39032 0 spi_dac_i_2.spi_dat_buff\[0\]
rlabel metal2 35728 31864 35728 31864 0 spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal3 35952 33880 35952 33880 0 spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 40880 41272 40880 41272 0 spi_dac_i_2.spi_dat_buff\[1\]
rlabel metal2 43848 39088 43848 39088 0 spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 44184 40712 44184 40712 0 spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal3 41440 37800 41440 37800 0 spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 41160 36120 41160 36120 0 spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal3 35224 35784 35224 35784 0 spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal3 35896 34888 35896 34888 0 spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal2 36232 34776 36232 34776 0 spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal3 37184 30632 37184 30632 0 spi_dac_i_2.spi_dat_buff\[9\]
<< properties >>
string FIXED_BBOX 0 0 46000 46000
<< end >>
