* NGSPICE file created from tholin_avalonsemi_tbb1143.ext - technology: gf180mcuD

.subckt tholin_avalonsemi_tbb1143 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] rst_n vdd vss
.ends

