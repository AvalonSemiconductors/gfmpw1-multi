* NGSPICE file created from wrapped_sn76489.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

.subckt wrapped_sn76489 custom_settings[0] custom_settings[1] io_in_1[0] io_in_1[1]
+ io_in_1[2] io_in_1[3] io_in_1[4] io_in_1[5] io_in_1[6] io_in_1[7] io_in_2 io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[17] io_out[18] io_out[19] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] rst_n vdd vss wb_clk_i io_out[15] io_out[14]
+ io_out[13] io_out[3] io_out[2] io_out[1] io_out[16]
X_2106_ _0373_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2037_ _0328_ _0329_ _0331_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2084__B _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1270_ _0715_ _0716_ _0718_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_58_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2655_ _0129_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1606_ _1048_ _1049_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2586_ _0060_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1537_ _0951_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1468_ _0911_ _0916_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1399_ _0839_ _0847_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_69_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1978__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2079__B _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1666__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2672__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2440_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\] _0648_ _0646_ _0649_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1672__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2371_ _0599_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1322_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\] _0771_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_75_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2707_ _0181_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2545__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2638_ _0112_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2569_ _0043_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2695__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Left_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_76_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1887__A1 _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1940_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\] _0252_ _0255_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2568__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1871_ _0194_ _0202_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2119__A2 _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2423_ _1104_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2354_ _0587_ _0137_ _0588_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1305_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\] _0754_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2285_ tt_um_rejunity_sn76489.pwm.accumulator\[4\] net19 _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2447__B _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1577__I _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2710__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2070_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\] _0358_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
+ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1923_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\] _0238_ _0243_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1854_ _1252_ _1253_ _1254_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1785_ _1195_ _1197_ _1157_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2406_ _0614_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2337_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\] tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\]
+ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\] _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2268_ tt_um_rejunity_sn76489.pwm.accumulator\[2\] _0521_ _0522_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2276__A1 _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2199_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\] _0465_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
+ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_79_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2200__A1 _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _1006_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2606__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2122_ _0280_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2053_ _0343_ _0344_ _0330_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1906_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\] tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
+ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\] _0952_ tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
+ tt_um_rejunity_sn76489.control_noise\[0\]\[1\] _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1837_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\] _0892_ _1240_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1768_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\] _0818_ _1183_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1699_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\] _1122_ _1127_ _1128_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2249__A1 _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2629__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput20 net20 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2488__A1 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2671_ _0145_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1622_ _1063_ _1064_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1553_ _0997_ _0998_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1484_ _0909_ _0910_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2479__A1 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2105_ _0388_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2036_ _0328_ _0329_ _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2403__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2654_ _0128_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2585_ _0059_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1605_ _0960_ _0844_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1536_ _0976_ _0979_ _0981_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1467_ _0830_ _0912_ _0915_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1398_ _0840_ _0841_ _0843_ _0844_ _0846_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_49_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2019_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\] _0869_ _0316_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_45_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2526__D _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2114__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2370_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\] _0596_ _0593_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\]
+ _0597_ net22 _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1321_ _0767_ _0769_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_75_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2706_ _0180_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2637_ _0111_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2568_ _0042_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2499_ _0690_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1519_ _0963_ _0936_ _0835_ _0965_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__1812__B _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1870_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\] _1026_ _0201_ _0202_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_43_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2422_ _0634_ _0629_ _0636_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2353_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\] _0000_ _0132_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\]
+ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1304_ _0750_ _0751_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2284_ _0533_ _0535_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2055__A2 _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1999_ _0299_ _0296_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\] _0301_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2662__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2285__A2 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2535__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1922_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\] _0241_ _0242_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2685__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1853_ _1252_ _1253_ _1238_ _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1784_ _1196_ _1032_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2405_ _0622_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2336_ _0575_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\] tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\]
+ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2267_ _0824_ _0864_ _0821_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_79_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2198_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
+ _0463_ _0464_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_67_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2193__B _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2558__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2122__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2121_ _0365_ _0398_ _0401_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2052_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\] _1018_ _0344_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1905_ _0220_ _0227_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1836_ _1236_ _1237_ _1239_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1767_ _1171_ _1182_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1698_ _1126_ _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2700__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2319_ _0560_ _0563_ _0564_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_input11_I io_in_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput21 net21 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2670_ _0144_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1621_ _1046_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1552_ _0966_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1483_ _0928_ _0930_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input3_I io_in_1[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2104_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\] _0384_ _0386_ _0387_ _0377_
+ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2035_ _0209_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_80_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1819_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\] _1051_ _1224_ _1226_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1914__A1 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1905__A1 _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2653_ _0127_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2584_ _0058_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1604_ _0777_ _0815_ _0781_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_10_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1535_ _0971_ _0975_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1466_ _0913_ _0914_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1397_ _0840_ _0841_ _0845_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__2321__A1 _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2619__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2018_ _1210_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1320_ _0768_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2705_ _0179_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2636_ _0110_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2567_ _0041_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2498_ _0690_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1518_ _0964_ _0936_ _0825_ _0963_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1449_ _0867_ _0896_ _0897_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_2_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2591__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2421_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\] _0635_ _0624_ _0636_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2524__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2352_ _0820_ _0515_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1303_ tt_um_rejunity_sn76489.chan\[0\].attenuation.in _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2283_ _0224_ _0534_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_15_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1998_ _0299_ _0296_ _0300_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2619_ _0093_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2506__A1 _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1921_ _0231_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1852_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\] _1028_ _1253_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1783_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[4\] _1196_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2404_ net8 _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2335_ _0575_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\] _0576_ _0133_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2266_ _0513_ _0518_ _0519_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2197_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
+ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
+ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_46_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_26_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1728__B _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2120_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\] _0389_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
+ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_77_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2051_ _0341_ _0342_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2652__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1904_ tt_um_rejunity_sn76489.clk_counter\[6\] _0225_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1835_ _1236_ _1237_ _1238_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1766_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\] _0818_ _1181_ _1182_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_4_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2194__A2 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1697_ _1097_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2318_ tt_um_rejunity_sn76489.pwm.accumulator\[9\] net24 _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2249_ _0286_ _0492_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_23_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2185__A2 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput22 net22 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1696__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2675__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ _1045_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1551_ _0962_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1482_ _0735_ _0929_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2289__B _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1687__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2103_ _0380_ _0385_ _0381_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1439__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2034_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\] _0973_ _0329_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_80_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2548__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1818_ _1211_ _1225_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_15_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1749_ _1165_ _1167_ _1168_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2698__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2218__I _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1841__A1 _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2652_ _0126_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2583_ _0057_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1603_ _1045_ _1046_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1534_ _0980_ net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1465_ _0889_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1396_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _0754_ _0756_ _0845_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2017_ _0312_ _0313_ _0314_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2713__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2379__A2 _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1697__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2704_ _0178_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2635_ _0109_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2566_ _0040_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2497_ _0655_ _0689_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1517_ _0780_ _0833_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1448_ _0872_ _0895_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_27_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1379_ _0808_ _0810_ _0826_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_53_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2297__A1 _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2609__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2420_ _0628_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1980__I _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2351_ _0586_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1302_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _0751_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2282_ _0530_ _0532_ _0531_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_63_Left_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_72_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1997_ _0299_ _0296_ _0210_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2618_ _0092_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2549_ _0023_ clknet_4_11_0_wb_clk_i net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_3_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_64_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1920_ _0236_ _0239_ _0240_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1851_ _1247_ _1031_ _1251_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1782_ _1191_ _1193_ _1194_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_24_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2581__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2403_ _0620_ _0612_ _0621_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2334_ _0575_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\] _1077_ _0223_ _0576_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_46_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2265_ tt_um_rejunity_sn76489.pwm.accumulator\[1\] _0516_ _0519_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2196_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
+ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\] tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
+ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__1484__A2 _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2050_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\] _1015_ _0338_ _0342_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2415__A1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1903_ _0222_ _0226_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1834_ _1126_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1765_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\] _1179_ _1181_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1696_ _1102_ _1121_ _1125_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2317_ tt_um_rejunity_sn76489.pwm.accumulator\[8\] net23 _1062_ tt_um_rejunity_sn76489.pwm.accumulator\[9\]
+ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2248_ _0504_ _0506_ _1132_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2179_ _0396_ _0449_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput23 net23 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_58_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1550_ _0992_ _0995_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1481_ _0850_ _0906_ _0747_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2102_ _0380_ _0385_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2033_ _0323_ _0924_ _0327_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_76_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1817_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\] _1051_ _1224_ _1225_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1748_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\] _1014_ _1168_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1679_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\] _1112_ _1099_ _1114_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2642__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2651_ _0125_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1602_ _0953_ _0721_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2582_ _0056_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1533_ _0976_ _0979_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1464_ _0885_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1395_ _0760_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2016_ _0312_ _0313_ _0210_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2665__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2538__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1511__A1 _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2688__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2703_ _0177_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2634_ _0108_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2565_ _0039_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1516_ _0813_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2496_ _0627_ _0669_ _0679_ _0668_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1447_ _0872_ _0895_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1378_ _0808_ _0810_ _0826_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2350_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\] _0000_ _0511_ _0585_
+ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1301_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\] _0750_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_2281_ _0530_ _0531_ _0532_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_67_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1996_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\] _0299_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2617_ _0091_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2703__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2548_ _0022_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2479_ _0634_ _0672_ _0677_ _0676_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_65_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_21_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1714__A1 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1850_ _1246_ _1250_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1781_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\] _0913_ _1194_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2402_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\] _0617_ _0615_ _0621_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2333_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\] _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2264_ tt_um_rejunity_sn76489.pwm.accumulator\[1\] _0516_ _0518_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2195_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\] _0403_ _0462_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1979_ _0276_ _0277_ _0284_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_55_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2121__A1 _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2188__A1 _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1760__B _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1902_ _0224_ _0225_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2179__A1 _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1833_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\] _0892_ _1237_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1764_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\] _1179_ _1180_ _0024_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1654__C _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1695_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\] _1122_ _1115_ _1125_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2316_ _0558_ _0561_ _0562_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2247_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\] _0396_ _0505_ _0506_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2178_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\] _0444_ _0448_ _0449_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2006__B _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput24 net24 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput13 net13 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2571__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1480_ _0719_ _0927_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2101_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\] _0373_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
+ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2032_ _0322_ _0326_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1816_ _1219_ _1055_ _1223_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1665__B _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1375__A2 _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1747_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\] _1014_ _1167_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1678_ _1107_ _1111_ _1113_ _1093_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2594__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_59_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2650_ _0124_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1601_ _0797_ _0851_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2581_ _0055_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1532_ _0922_ _0977_ _0978_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1463_ _0891_ _0847_ _0885_ _0889_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1394_ _0750_ _0804_ _0842_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA_input1_I custom_settings[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2015_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\] _0869_ _0313_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2702_ _0176_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2633_ _0107_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.chan\[1\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2564_ _0038_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1515_ _0809_ _0959_ _0961_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_10_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2495_ _1104_ _0682_ _0688_ _0686_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_10_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1446_ _0882_ _0890_ _0894_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1377_ _0774_ _0778_ _0816_ _0814_ _0825_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_65_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2632__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1763__B _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1300_ _0722_ _0728_ _0743_ _0748_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_2280_ _0524_ _0525_ _0527_ _0529_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2655__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1995_ _0296_ _0298_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2616_ _0090_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2547_ _0021_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2478_ _0715_ _0673_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1429_ _0715_ _0877_ _0726_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_38_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2528__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2678__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1650__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1780_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\] _0913_ _1193_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2401_ _1108_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2332_ _0574_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2263_ _0456_ _0517_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2194_ _0833_ _0457_ _0461_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2130__A2 _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1978_ _0275_ net1 _0279_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2360__A2 _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1871__A1 _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1901_ tt_um_rejunity_sn76489.clk_counter\[5\] tt_um_rejunity_sn76489.clk_counter\[4\]
+ _0219_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_32_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1832_ _1232_ _1234_ _1235_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_4_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1763_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\] _1179_ _1157_ _1180_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1694_ _1096_ _1121_ _1124_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2315_ _0558_ _0561_ _0539_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2246_ _0281_ _0500_ _0503_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_69_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2177_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\] _0441_ _0448_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_75_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2073__I _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput25 net25 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput14 net14 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2716__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2100_ _0361_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2031_ _0323_ _0924_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1815_ _1218_ _1222_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1746_ _1142_ _1166_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1677_ net3 _1112_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2229_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\] _0355_ _0489_ _0490_ _0482_
+ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_67_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2260__A1 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2012__A1 _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1600_ _1024_ _1037_ _1021_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2580_ _0054_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1531_ _0926_ _0944_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1462_ _0909_ _0910_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1393_ tt_um_rejunity_sn76489.chan\[0\].attenuation.in _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2014_ _0307_ _0801_ _0310_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_54_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2561__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1729_ _1149_ _1151_ _1152_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2481__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2701_ _0175_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2584__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2632_ _0106_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2563_ _0037_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1514_ _0960_ _0845_ _0888_ _0809_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_10_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ _0777_ _0683_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1445_ _0830_ _0848_ _0893_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1376_ _0773_ _0767_ _0775_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_65_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Left_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1496__A2 _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2445__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2166__I _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1994_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\] _0293_ _0297_ _0298_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_41_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2615_ _0089_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2546_ _0020_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2477_ _1095_ _0672_ _0675_ _0676_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1428_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\] tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\]
+ _0717_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_50_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1359_ _0805_ _0806_ _0760_ _0807_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_33_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_12_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _1105_ _0611_ _0619_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2622__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2331_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\] _0573_ _0574_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2262_ tt_um_rejunity_sn76489.pwm.accumulator\[1\] _0513_ _0516_ _0517_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2193_ _0833_ _0457_ _0460_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1469__A2 _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2418__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ _1140_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1684__B _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2529_ _0003_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1703__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_7_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2645__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1900_ _0223_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1831_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\] _0811_ _1235_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1762_ _0779_ _0784_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1693_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\] _1122_ _1115_ _1124_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2314_ _0559_ _0560_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2245_ _0287_ _0500_ _0503_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2176_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\] _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1679__B _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2303__B _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput15 net15 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput26 net26 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_66_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2030_ _0322_ _0324_ _0325_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1814_ _1219_ _1055_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1745_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\] _1014_ _1165_ _1166_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_4_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1676_ _1110_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2228_ _0485_ _0488_ _0475_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2159_ _0428_ _0432_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2260__A2 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1530_ _0926_ _0944_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1461_ _0778_ _0834_ _0779_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1392_ _0751_ _0762_ _0752_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_54_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2013_ _0309_ _0311_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1801__I _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2706__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1728_ _1149_ _1151_ _1127_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1659_ _1097_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_36_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1621__I _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2700_ _0174_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2631_ _0105_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2562_ _0036_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1513_ _0750_ _0842_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2493_ _1101_ _0682_ _0687_ _0686_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1444_ _0891_ _0892_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1375_ _0802_ _0819_ _0823_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_73_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2551__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1993_ _1098_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_15_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2614_ _0088_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1708__A1 _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2545_ _0019_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2476_ _1092_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1427_ _0732_ _0873_ _0874_ _0742_ _0875_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1358_ _0758_ _0762_ _0752_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1289_ tt_um_rejunity_sn76489.chan\[3\].attenuation.in _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_66_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2574__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2330_ _1078_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2261_ _0802_ _0819_ _0515_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2192_ _0209_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_63_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1976_ _0220_ _0282_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2528_ _0002_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2597__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2459_ _0654_ _0661_ _0663_ _1093_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_19_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2036__B _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1830_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\] _0811_ _1234_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1785__B _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1761_ _1177_ _1175_ _1178_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1692_ _1118_ _1121_ _1123_ _1093_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_40_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2313_ _0553_ _0554_ _0556_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2244_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\] _0492_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
+ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2175_ _0446_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1695__B _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1959_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\] _0260_ _0269_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput16 net16 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput27 net27 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2612__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1813_ _1218_ _1220_ _1221_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1744_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\] _0984_ _1164_ _1165_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_40_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1675_ _1110_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2227_ _0485_ _0488_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2158_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\] _0426_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
+ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2635__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2089_ _0370_ _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_10_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1460_ _0844_ _0845_ _0761_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1391_ _0758_ _0763_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2658__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2012_ _0224_ _0310_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1727_ _1150_ _0923_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1692__C _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1658_ net12 _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1589_ _1030_ _0967_ _1033_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_48_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_47_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1680__A1 _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2630_ _0104_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2561_ _0035_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2492_ _0815_ _0683_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1512_ _0806_ _0807_ _0843_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1443_ _0847_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1374_ _0822_ _0796_ _0799_ _0800_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_58_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output19_I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1662__A1 _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1992_ _0295_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2613_ _0087_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2544_ _0018_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2475_ _0716_ _0673_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1426_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\] _0737_ _0730_ _0875_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_76_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1357_ _0750_ _0754_ _0752_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_1288_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _0737_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_TAPCELL_ROW_66_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1717__I _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2124__A2 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2260_ _0785_ _0786_ _0514_ _0749_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2191_ _0456_ _0459_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1975_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\] _0281_ _0282_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1537__I _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2527_ _0001_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2354__A2 _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2458_ _0795_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1409_ _0716_ _0723_ _0718_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2389_ _0610_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2042__A1 _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2541__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2691__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1760_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\] _1064_ _1157_ _1178_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1691_ net3 _1122_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_29_Left_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2312_ tt_um_rejunity_sn76489.pwm.accumulator\[8\] net23 _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2243_ _0498_ _0353_ _0501_ _0502_ _1141_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2174_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\] _0425_ _0443_ _0445_ _0439_
+ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_73_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1958_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\] _0263_ _0268_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1889_ _0212_ tt_um_rejunity_sn76489.clk_counter\[1\] tt_um_rejunity_sn76489.clk_counter\[2\]
+ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2564__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput17 net17 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 net28 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2047__B _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2263__A1 _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2510__B _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1829__A1 _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2587__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1812_ _1218_ _1220_ _1203_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1743_ _1161_ _1163_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1674_ _1086_ _1109_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2226_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\] _0478_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
+ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2157_ _0431_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2493__A1 _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2088_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\] _0373_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
+ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2245__A1 _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2381__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1390_ _0832_ _0835_ _0837_ _0838_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2011_ _0305_ _0308_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1726_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[4\] _1150_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1657_ _1095_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1588_ _1031_ _1032_ _0968_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2602__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2209_ _0470_ _0473_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2466__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_55_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2625__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2560_ _0034_ clknet_4_11_0_wb_clk_i net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2491_ _1095_ _0682_ _0685_ _0686_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1511_ _0951_ _0957_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1442_ _0839_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1373_ _0794_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1709_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\] _0822_ _1135_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2689_ _0163_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2648__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1991_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\] _0293_ _0295_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_27_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2612_ _0086_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2543_ _0017_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2474_ _0654_ _0672_ _0674_ _0665_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1425_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _0731_ _0874_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1356_ _0803_ _0804_ _0763_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1287_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\] _0736_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_66_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1643__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2190_ _0453_ _0458_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1974_ _0280_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2526_ _0000_ clknet_4_14_0_wb_clk_i net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2457_ _0660_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1408_ _0712_ _0724_ _0713_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2388_ _0610_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1339_ _0722_ _0728_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_78_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1690_ _1120_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2311_ tt_um_rejunity_sn76489.pwm.accumulator\[9\] net24 _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2242_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\] _0499_ _0495_ _0502_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2173_ _0289_ _0444_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2709__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1957_ _0266_ _0267_ _0262_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1548__I _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1888_ _1140_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput18 net18 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2509_ _1085_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2254__A2 _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1811_ _1219_ _1055_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_25_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1742_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\] _0984_ _1163_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1673_ _1081_ _1108_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2225_ _0487_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2156_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\] _0425_ _0428_ _0430_ _0419_
+ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1296__A3 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2087_ _0358_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2531__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2681__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2236__A2 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_57_Left_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_66_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1651__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2010_ _0305_ _0308_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2554__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_75_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1725_ _1145_ _1147_ _1148_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1656_ _1094_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1587_ _0910_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2208_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\] _0465_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
+ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2139_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\] _0413_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
+ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2392__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2577__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2490_ _0223_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1510_ _0727_ _0955_ _0956_ _0861_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1441_ _0885_ _0889_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1372_ _0749_ _0791_ _0820_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_65_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2688_ _0162_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1708_ _1132_ _1134_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1639_ _1079_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_69_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1990_ _0293_ _0294_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2611_ _0085_ clknet_4_11_0_wb_clk_i net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2542_ _0016_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2473_ _0723_ _0673_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1424_ _0850_ _0741_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1355_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _0804_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1286_ _0732_ _0733_ _0734_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_66_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2615__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2348__A1 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2520__A1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2490__I _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1973_ _0275_ net1 _0278_ _0279_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_7_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2525_ _0706_ _0703_ _0707_ _0695_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2456_ _0660_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1407_ _0715_ _0718_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2387_ _0606_ _0607_ _0608_ _0609_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__2511__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2638__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1338_ _0785_ _0786_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1269_ _0717_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2508__C _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2243__C _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2310_ _0541_ _0557_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2241_ _0396_ _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2172_ _0437_ _0442_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1956_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\] _0260_ _0267_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_31_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1887_ _0194_ _0214_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 net19 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2508_ _1104_ _0691_ _0697_ _0695_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2439_ _0642_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2519__B _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1810_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[8\] _1219_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_25_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1741_ _1142_ _1162_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1672_ net7 _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2224_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\] _0468_ _0485_ _0486_ _0482_
+ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2155_ _0422_ _0427_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2086_ _0372_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1939_ _0253_ _0254_ _0251_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2181__A2 _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1683__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1724_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\] _0901_ _1148_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1655_ net4 _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1586_ _0909_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2207_ _0472_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2138_ _0410_ _0415_ _0213_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2069_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
+ _0356_ _0357_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_14_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1752__I _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1701__B _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1440_ _0803_ _0886_ _0887_ _0888_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_1371_ _0802_ _0819_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2671__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2687_ _0161_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1707_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\] _0822_ _1133_ _1134_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_41_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1638_ _1076_ _1078_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1569_ _1004_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_69_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2544__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2127__A2 _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2694__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1657__I _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2610_ _0084_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2541_ _0015_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2472_ _0671_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1423_ _0868_ _0863_ _0871_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1354_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\] _0803_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1877__A1 _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1285_ _0729_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_66_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2567__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1972_ tt_um_rejunity_sn76489.clk_counter\[0\] tt_um_rejunity_sn76489.clk_counter\[1\]
+ tt_um_rejunity_sn76489.clk_counter\[3\] tt_um_rejunity_sn76489.clk_counter\[2\]
+ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_71_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2524_ net5 _0703_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2455_ _0655_ _0659_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2386_ tt_um_rejunity_sn76489.latch_control_reg\[2\] _1084_ _0609_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1406_ _0849_ _0850_ _0851_ _0852_ _0854_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1337_ _0761_ _0766_ _0779_ _0784_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1268_ _0708_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2240_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\] _0495_ _0499_ _0500_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2171_ _0437_ _0442_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1955_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\] _0263_ _0266_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_31_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1886_ _0212_ tt_um_rejunity_sn76489.clk_counter\[1\] _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_3_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2605__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2507_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _0692_ _0697_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2438_ _0632_ _0643_ _0647_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2369_ _0598_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_39_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1462__A2 _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2628__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1740_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\] _0984_ _1161_ _1162_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1671_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\] _1107_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input8_I io_in_1[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2223_ _0480_ _0484_ _0475_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2154_ _0288_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2085_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\] _0362_ _0370_ _0371_ _0297_
+ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_36_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1938_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\] _0249_ _0254_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1869_ _0197_ _0199_ _0200_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2090__B _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1380__A1 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1723_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\] _0901_ _1147_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1654_ _1080_ _1088_ _1090_ _1093_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1585_ _1028_ _1029_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2206_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\] _0468_ _0470_ _0471_ _0439_
+ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2137_ _0355_ _0414_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2068_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
+ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
+ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1370_ _0811_ _0818_ _0785_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_65_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2686_ _0160_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1706_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\] _0788_ _1133_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1637_ net12 _1077_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1568_ _1011_ _1012_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1499_ _0946_ net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_69_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2540_ _0014_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2471_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1422_ _0869_ _0870_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1353_ _0794_ _0801_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1284_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _0733_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_66_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2669_ _0143_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1668__I _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1971_ _0276_ _0277_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2523_ tt_um_rejunity_sn76489.control_noise\[0\]\[2\] _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2454_ _0656_ _0657_ _0658_ _0609_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2385_ net11 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1405_ _0849_ _0850_ _0853_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1336_ _0761_ _0766_ _0779_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
Xinput1 custom_settings[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1267_ _0711_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2534__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2684__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2202__I _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2170_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\] _0441_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
+ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2557__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1954_ _0264_ _0265_ _0262_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1885_ _0212_ _0213_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2506_ _1101_ _0691_ _0696_ _0695_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2437_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\] _0644_ _0646_ _0647_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1861__I _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2368_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\] _0596_ _0593_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\]
+ _0597_ net21 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1319_ tt_um_rejunity_sn76489.chan\[1\].attenuation.in _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2299_ tt_um_rejunity_sn76489.pwm.accumulator\[6\] _0980_ _0543_ _0544_ _0548_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_39_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2184__A1 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1670_ _1105_ _1088_ _1106_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1681__I _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2222_ _0480_ _0484_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2153_ _0422_ _0427_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2084_ _0364_ _0369_ _0366_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1937_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\] _0252_ _0253_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1868_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\] _0994_ _0200_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1799_ _1207_ _1208_ _1209_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_26_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_35_Left_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_33_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1722_ _1142_ _1146_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1653_ _1092_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_44_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1584_ _0939_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1371__A2 _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2205_ _0466_ _0469_ _0429_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_53_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2136_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\] _0413_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
+ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2067_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
+ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\] tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
+ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_17_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_62_Left_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2210__I _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2618__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2085__C _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1705_ _1131_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2685_ _0159_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1636_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\] tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
+ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1592__A2 _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1567_ _0976_ _0979_ _0987_ _1009_ _0981_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_1_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1498_ _0922_ _0945_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_69_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2186__B _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2119_ _0395_ _0353_ _0399_ _0400_ _0283_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_1_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2590__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2470_ _0655_ _0670_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1421_ _0862_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1352_ _0796_ _0799_ _0800_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_1283_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\] _0732_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_66_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2668_ _0142_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1619_ _1062_ net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_6_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2599_ _0073_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2505__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1970_ _0275_ net1 _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_11_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2522_ _0632_ _0703_ _0705_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2453_ _0606_ tt_um_rejunity_sn76489.latch_control_reg\[0\] _0658_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2384_ tt_um_rejunity_sn76489.latch_control_reg\[0\] _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1404_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\] _0795_ _0734_ _0853_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1335_ _0782_ _0776_ _0783_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xinput2 custom_settings[1] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1266_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\] _0715_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\] _0260_ _0265_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1884_ _1131_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2193__A2 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2505_ _0803_ _0692_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2436_ _0614_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2367_ _0581_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1318_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] _0767_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2298_ tt_um_rejunity_sn76489.pwm.accumulator\[6\] net21 _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2651__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2221_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\] _0478_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
+ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2152_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\] _0426_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
+ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2674__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2083_ _0364_ _0369_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_36_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1936_ _0231_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1867_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\] _0994_ _0199_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1798_ _1207_ _1208_ _1203_ _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2419_ _1101_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1677__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2547__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2697__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1721_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\] _0901_ _1145_ _1146_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_13_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1652_ _1091_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1583_ _0935_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2204_ _0466_ _0469_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2135_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
+ _0411_ _0412_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2066_ _0288_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_48_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1919_ _0235_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2712__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ _1130_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2684_ _0158_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1635_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\] _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1566_ _0987_ _1009_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_18_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1497_ _0926_ _0944_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_69_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2118_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\] _0397_ _0392_ _0400_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2049_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\] _1015_ _0341_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1420_ _0855_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1351_ _0733_ _0746_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1282_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\] _0730_ _0731_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2608__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2667_ _0141_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1618_ _1043_ _1061_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_6_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2598_ _0072_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1549_ _0993_ _0994_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_66_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1492__A2 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2441__A1 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2521_ tt_um_rejunity_sn76489.control_noise\[0\]\[1\] _0702_ _1092_ _0705_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2452_ net9 net10 _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2383_ tt_um_rejunity_sn76489.latch_control_reg\[1\] _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1403_ _0736_ _0733_ _0739_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1334_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\] _0768_ _0783_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1265_ _0710_ _0712_ _0713_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xinput3 io_in_1[0] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2580__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output15_I net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2390__B _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1952_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\] _0263_ _0264_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1883_ tt_um_rejunity_sn76489.clk_counter\[0\] _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2504_ _1095_ _0691_ _0694_ _0695_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2435_ _0605_ _0643_ _0645_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2459__C _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2366_ _1079_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1317_ _0753_ _0764_ _0765_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2297_ _0541_ _0546_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2404__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2220_ _0483_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2151_ _0413_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2082_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\] _0358_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
+ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1935_ _0248_ _0250_ _0251_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1866_ _0194_ _0198_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1797_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\] _0998_ _1208_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2418_ _0632_ _0629_ _0633_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2349_ _0581_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1720_ _1143_ _1144_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_53_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1651_ net12 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2641__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1582_ _0963_ _0832_ _0836_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1356__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2203_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\] _0465_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
+ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input6_I io_in_1[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2134_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
+ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
+ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2065_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\] _0353_ _0354_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1918_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\] _0238_ _0239_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1849_ _1247_ _1031_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2664__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1338__A1 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_9_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1968__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1703_ net12 _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_1_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2683_ _0157_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1634_ _1075_ net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1565_ _1010_ net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_1_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1496_ _0931_ _0943_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_69_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2537__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2117_ _0396_ _0398_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2048_ _0338_ _0339_ _0340_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2687__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1559__A1 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1350_ _0797_ _0742_ _0798_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1281_ _0729_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2666_ _0140_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1617_ _1044_ _1060_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2597_ _0071_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1548_ _0991_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1479_ _0857_ _0904_ _0727_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_69_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_59_Left_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2702__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1713__A1 _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2142__I _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2520_ _0605_ _0703_ _0704_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2451_ _1081_ _1082_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1981__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1402_ _0742_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2382_ _0604_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1333_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _0780_ _0781_ _0782_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1264_ tt_um_rejunity_sn76489.chan\[2\].attenuation.in _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput4 io_in_1[1] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2718_ _0192_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.control_noise\[0\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2649_ _0123_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1951_ _0230_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1882_ _0208_ _0206_ _0211_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2503_ _0223_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2434_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\] _0644_ _0638_ _0645_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2365_ _0595_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1316_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _0755_ _0765_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_47_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2296_ tt_um_rejunity_sn76489.pwm.accumulator\[6\] net21 _0545_ _0546_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_39_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2150_ _0361_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2081_ _0368_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2570__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1934_ _0234_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1865_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\] _0994_ _0197_ _0198_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1796_ _1205_ _1206_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2417_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\] _0630_ _0624_ _0633_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2348_ _0283_ _0582_ _0584_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2279_ tt_um_rejunity_sn76489.pwm.accumulator\[4\] _0898_ _0919_ _0531_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_79_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2593__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1650_ net3 _1089_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1581_ _1025_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2150__I _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2202_ _0361_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2133_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
+ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\] tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
+ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2064_ _0280_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1292__A1 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1917_ _0237_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1848_ _1246_ _1248_ _1249_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_31_Left_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1779_ _1171_ _1192_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_40_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_55_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1338__A2 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2682_ _0156_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1702_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\] _0788_ _1129_ _0013_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1633_ _1067_ _1069_ _1074_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1564_ _0982_ _0987_ _1009_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_1495_ _0941_ _0942_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_55_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2116_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\] _0392_ _0397_ _0398_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2047_ _0338_ _0339_ _0330_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2631__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2508__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1280_ tt_um_rejunity_sn76489.chan\[3\].attenuation.in _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2665_ _0139_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2596_ _0070_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1970__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1616_ _1047_ _1059_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1547_ _0989_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1478_ _0923_ _0924_ _0925_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2654__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2423__I _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2527__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2450_ _0608_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1401_ _0737_ _0744_ _0738_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_2381_ net3 _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1332_ _0768_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2677__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1263_ _0711_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xinput5 io_in_1[2] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2717_ _0191_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.control_noise\[0\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2648_ _0122_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2579_ _0053_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.chan\[3\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_76_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1950_ _0259_ _0261_ _0262_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1881_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\] _1052_ _0210_ _0211_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_78_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2502_ _0804_ _0692_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2433_ _0642_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2364_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\] _0589_ _0593_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\]
+ _0585_ net20 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1315_ _0758_ _0762_ _0763_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2350__A2 _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2295_ _0543_ _0544_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2080_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\] _0362_ _0364_ _0367_ _0297_
+ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2715__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1933_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\] _0249_ _0250_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1864_ _0195_ _0196_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1795_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\] _1029_ _1201_ _1206_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_12_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2416_ _1094_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2347_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\] _0575_ _0583_ _0584_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2278_ _0529_ _0527_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1580_ _0843_ _0886_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2201_ _0462_ _0467_ _1132_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2132_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\] _0403_ _0410_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _0352_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_76_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2241__A1 _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1916_ tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
+ _0229_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1847_ _1246_ _1248_ _1238_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1778_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\] _0913_ _1191_ _1192_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_55_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2663__D _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2560__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2681_ _0155_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1701_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\] _0788_ _1127_ _1129_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1632_ _1070_ _1072_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1563_ _1002_ _1008_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_1_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1494_ _0932_ _0933_ _0940_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2115_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\] _0389_ _0397_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2046_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\] _1015_ _0339_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2462__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2583__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_sn76489_40 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_39_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_14_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2664_ _0138_ clknet_4_13_0_wb_clk_i net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2595_ _0069_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1615_ _1054_ _1058_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_1_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1546_ _0989_ _0991_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1477_ _0908_ _0917_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_66_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2435__A1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2029_ _0322_ _0324_ _0210_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1477__A2 _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2426__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1400_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\] _0730_ _0849_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2380_ _0215_ _0229_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2362__C2 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1331_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] _0780_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_79_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1262_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\] _0711_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput6 io_in_1[3] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2716_ _0190_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2647_ _0121_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2621__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2578_ _0052_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[6\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1529_ _0971_ _0975_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_25_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_76_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1880_ _0209_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2501_ _0654_ _0691_ _0693_ _0686_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2644__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2432_ _0642_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2363_ _0594_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1314_ _0755_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2294_ _0542_ _0946_ _0536_ _0534_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1669__B _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2667__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1932_ _0237_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1863_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\] _0997_ _1257_ _0196_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1794_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\] _1029_ _1205_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2415_ _0605_ _0629_ _0631_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2346_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\] tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
+ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2277_ tt_um_rejunity_sn76489.pwm.accumulator\[3\] _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2074__I _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2250__A2 _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2200_ _0289_ _0466_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2131_ _0952_ _0406_ _0409_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2062_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\] _1063_ _0351_ _1228_
+ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_76_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1915_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\] _0232_ _0236_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ _1247_ _1031_ _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1777_ _1185_ _1186_ _1190_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_12_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1682__B _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2329_ _0571_ _0569_ _0572_ _0215_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input12_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2705__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1611__I _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2680_ _0154_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1700_ _1105_ _1121_ _1128_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1631_ _1073_ net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1562_ _1007_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1493_ _0932_ _0933_ _0940_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input4_I io_in_1[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2114_ _0280_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2045_ _0334_ _0336_ _0337_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_52_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1829_ _1211_ _1233_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_68_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_sn76489_30 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_6_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2663_ _0137_ clknet_4_14_0_wb_clk_i net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2594_ _0068_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1614_ _1025_ _1055_ _1057_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1545_ _0764_ _0844_ _0846_ _0990_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__2380__A1 _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1476_ _0907_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_19_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2028_ _0323_ _0924_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_37_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2550__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2123__A1 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1330_ _0770_ _0772_ _0776_ _0778_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_79_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1261_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\] _0710_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xinput7 io_in_1[4] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2573__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2715_ _0189_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2646_ _0120_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2577_ _0051_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1528_ _0931_ _0943_ _0974_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_77_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1459_ _0905_ _0907_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2077__I _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2596__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2500_ _0754_ _0692_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2431_ _0606_ _0607_ _0608_ _0627_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2362_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\] _0589_ _0593_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\]
+ _0585_ net19 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1313_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\] _0762_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2293_ _0542_ _0946_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2629_ _0103_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2326__A1 _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1704__I _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1540__A2 _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1931_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\] _0241_ _0248_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2611__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1862_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\] _0997_ _0195_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput10 io_in_1[7] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1793_ _1201_ _1202_ _1204_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2414_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\] _0630_ _0624_ _0631_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2345_ _1076_ _1077_ net16 _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2276_ _0456_ _0528_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2634__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2130_ _0952_ _0406_ _0330_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_49_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2061_ _0346_ _0350_ _0347_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1914_ _0734_ _0232_ _0233_ _0235_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_44_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1845_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[4\] _1247_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_12_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1776_ _1187_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2328_ tt_um_rejunity_sn76489.pwm.accumulator\[11\] net26 _0572_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2657__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2259_ _0722_ _0728_ _0743_ _0748_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_55_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1440__A1 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1630_ _1070_ _1072_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1561_ _1004_ _1006_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1492_ _0935_ _0939_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2113_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\] _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2044_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\] _0983_ _0337_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1670__A1 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\] _0811_ _1232_ _1233_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1973__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1693__B _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1759_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\] _1064_ _1177_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_13_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_68_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2029__B _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_sn76489_31 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_26_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2662_ _0136_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2593_ _0067_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1613_ _1034_ _1035_ _0995_ _1056_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1544_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _0759_ _0990_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1475_ _0905_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2132__A2 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1891__A1 _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2027_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[4\] _0323_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_45_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1260_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\] _0708_ _0709_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2718__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 io_in_1[5] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ _0188_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.latch_control_reg\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2645_ _0119_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2576_ _0050_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2353__A2 _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1527_ _0972_ _0973_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1458_ _0906_ _0851_ _0743_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1389_ _0812_ _0780_ _0775_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_77_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1881__B _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1900__I _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2430_ _0623_ _0630_ _0641_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_47_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2540__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2361_ _0574_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1312_ _0753_ _0757_ _0759_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_47_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2292_ tt_um_rejunity_sn76489.pwm.accumulator\[5\] _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2690__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_56_Left_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2023__A1 _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_65_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2628_ _0102_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2559_ _0033_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_74_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2563__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1930_ _0246_ _0247_ _0240_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1861_ _1210_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput11 io_in_2 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1792_ _1201_ _1202_ _1203_ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2413_ _0628_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2344_ _0581_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2275_ tt_um_rejunity_sn76489.pwm.accumulator\[3\] _0526_ _0527_ _0528_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_59_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2586__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1715__I _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2235__A1 _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2060_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\] _1063_ _0350_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2474__A1 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1913_ _0234_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1844_ _1242_ _1244_ _1245_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1775_ _1171_ _1189_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2327_ tt_um_rejunity_sn76489.pwm.accumulator\[11\] net26 _0571_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2258_ tt_um_rejunity_sn76489.pwm.accumulator\[0\] _0511_ _0513_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2189_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\] _0457_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
+ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2465__A1 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2315__B _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_3_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1560_ _0854_ _0851_ _0745_ _1005_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_39_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1491_ _0825_ _0936_ _0938_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2112_ _0394_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2119__C _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2043_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\] _0983_ _0336_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\] _1230_ _1232_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2624__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1758_ _1171_ _1176_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1689_ _1120_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2438__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_sn76489_32 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2647__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2661_ _0135_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1612_ _1025_ _1027_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2592_ _0066_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1543_ _0936_ _0988_ _0963_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1474_ _0898_ _0919_ _0921_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_66_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2026_ _0318_ _0320_ _0321_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_9_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 io_in_1[6] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_62_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2713_ _0187_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.latch_control_reg\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2644_ _0118_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.chan\[0\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2575_ _0049_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[3\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1526_ _0930_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1457_ _0853_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1388_ _0813_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1699__B _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2009_ _0307_ _0801_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2360_ _0527_ _0137_ _0592_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1311_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\] _0756_ _0760_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_2291_ _1131_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2627_ _0101_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2558_ _0032_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2489_ _0812_ _0683_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1509_ _0953_ _0904_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2053__B _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2708__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2253__A2 _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1860_ _1257_ _1258_ _0193_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput12 rst_n net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1791_ _1126_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2412_ _0628_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2343_ _1130_ _1077_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2274_ _0867_ _0896_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1821__I _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2138__B _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1989_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\] _0292_ _1228_ _0294_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1286__A3 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2530__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2680__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1641__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1912_ _1130_ tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise _0234_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1843_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\] _0914_ _1245_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1774_ _1185_ _1188_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2326_ _0541_ _0570_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2257_ tt_um_rejunity_sn76489.pwm.accumulator\[0\] _0511_ _0512_ _0119_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2188_ _0286_ _0441_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2553__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1976__A1 _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1490_ _0832_ _0937_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2111_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\] _0384_ _0391_ _0393_ _0377_
+ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__2576__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2042_ _0315_ _0335_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\] _1230_ _1231_ _0035_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1757_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\] _1064_ _1175_ _1176_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1688_ _1081_ _1082_ _1119_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_40_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2309_ _0555_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input10_I io_in_1[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_51_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2126__A1 _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2599__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_74_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_sn76489_33 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_39_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1404__A3 _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2660_ _0134_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1611_ _1027_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2591_ _0065_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1542_ _0832_ _0835_ _0782_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1473_ _0903_ _0918_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2117__A1 _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I custom_settings[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2025_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\] _0900_ _0321_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1809_ _1214_ _1216_ _1217_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2614__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2712_ _0186_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.latch_control_reg\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2643_ _0117_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2574_ _0048_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[2\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1525_ _0928_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1561__A2 _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1456_ _0904_ _0721_ _0722_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1387_ _0773_ _0812_ _0775_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2008_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[1\] _0307_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2637__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2501__A1 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1644__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1310_ _0758_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\] _0756_ _0759_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2290_ _0537_ _0538_ _0540_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2626_ _0100_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ _0031_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2488_ _0654_ _0682_ _0684_ _0676_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1508_ _0953_ _0904_ _0954_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1439_ _0803_ _0751_ _0763_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2385__I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1790_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\] _1029_ _1202_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2411_ _0626_ _0607_ _0608_ _0627_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2342_ _0573_ _0580_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2273_ _0524_ _0525_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1988_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\] _0292_ _0293_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2609_ _0083_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1691__A1 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1911_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\] _0231_ _0233_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1842_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\] _0914_ _1244_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1773_ _1186_ _1187_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2325_ tt_um_rejunity_sn76489.pwm.accumulator\[11\] net26 _0569_ _0570_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2256_ tt_um_rejunity_sn76489.pwm.accumulator\[0\] _0511_ _0460_ _0512_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2187_ _1131_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2506__C _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2110_ _0289_ _0392_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2041_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\] _0983_ _0334_ _0335_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_9_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1825_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\] _1230_ _1203_ _1231_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1756_ _1169_ _1173_ _1174_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1687_ net9 _1085_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1894__A1 _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2308_ tt_um_rejunity_sn76489.pwm.accumulator\[8\] _1013_ _1039_ _0556_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2239_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\] _0492_ _0499_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2670__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2071__A1 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1637__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_sn76489_34 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_14_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1610_ _1050_ _1053_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2590_ _0064_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2543__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1541_ _0985_ _0986_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1472_ _0920_ net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2693__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2024_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\] _0900_ _0320_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_65_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1808_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\] _0993_ _1217_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1739_ _1159_ _1160_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2072__B _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2566__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_79_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2283__A1 _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_70_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2711_ _0185_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2642_ _0116_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2573_ _0047_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[1\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1524_ _0958_ _0970_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1455_ _0858_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1386_ _0773_ _0833_ _0834_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2007_ _0305_ _0306_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2589__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2514__C _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1660__I _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_25_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2625_ _0099_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_34_Left_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2556_ _0030_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2487_ _0767_ _0683_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1507_ _0953_ _0709_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1438_ _0804_ _0757_ _0765_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2495__A1 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1570__I _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1369_ _0812_ _0813_ _0817_ _0782_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XPHY_EDGE_ROW_43_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_21_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2334__C _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2604__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_61_Left_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2410_ tt_um_rejunity_sn76489.latch_control_reg\[2\] net10 _0627_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_2
X_2341_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\] _0578_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
+ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2272_ tt_um_rejunity_sn76489.pwm.accumulator\[2\] _0521_ _0520_ _0525_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2477__A1 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1987_ _0283_ _0290_ _0292_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2627__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2608_ _0082_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2539_ _0013_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2329__C _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2345__B net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2459__A1 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1910_ _0231_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1985__A3 _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1841_ _1211_ _1243_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1772_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\] _0891_ _1187_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2324_ _0565_ _0567_ _0568_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2255_ _0787_ _0790_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2186_ _0453_ _0455_ _1132_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2040_ _0328_ _0332_ _0333_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_71_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1824_ _0761_ _0766_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1755_ _1172_ _1022_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1686_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\] _1118_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2307_ _0553_ _0554_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2238_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\] _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2169_ _0426_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1885__A2 _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwrapped_sn76489_35 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_14_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1540_ _0958_ _0970_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1663__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1471_ _0898_ _0919_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2023_ _0315_ _0319_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_65_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_73_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1807_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\] _0993_ _1216_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_60_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1738_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\] _0972_ _1155_ _1160_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1669_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\] _1089_ _1099_ _1106_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1658__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2710_ _0184_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2641_ _0115_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2572_ _0046_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.clk_counter\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2660__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1546__A1 _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1523_ _0967_ _0969_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1454_ _0882_ _0899_ _0902_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1385_ _0771_ _0767_ _0769_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_2006_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\] _0789_ _0297_ _0306_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2683__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1700__A1 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1767__A1 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2624_ _0098_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2555_ _0029_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2486_ _0681_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1506_ _0710_ _0952_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1437_ _0760_ _0841_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1368_ _0814_ _0816_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2556__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1299_ _0745_ _0740_ _0747_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2247__A2 _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1758__A1 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2183__A1 _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2525__C _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2410__A2 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2340_ _0573_ _0579_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2579__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2271_ tt_um_rejunity_sn76489.pwm.accumulator\[2\] _0521_ _0524_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2229__A2 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1986_ _0291_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2607_ _0081_ clknet_4_14_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2538_ _0012_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1912__A1 _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2469_ _0657_ _0668_ _0669_ _0609_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_78_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2080__C _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1840_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\] _0914_ _1242_ _1243_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_4_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2395__A1 _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1771_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\] _0891_ _1186_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_69_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2323_ tt_um_rejunity_sn76489.pwm.accumulator\[10\] _1073_ _0568_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2254_ _0842_ _0507_ _0510_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2185_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\] _0403_ _0454_ _0455_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1969_ tt_um_rejunity_sn76489.clk_counter\[5\] tt_um_rejunity_sn76489.clk_counter\[4\]
+ tt_um_rejunity_sn76489.clk_counter\[6\] _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_43_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2310__A1 _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2129__A1 _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2617__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1823_ _1226_ _1229_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1754_ _1172_ _1022_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1685_ _1105_ _1111_ _1117_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2306_ _0550_ _1010_ _0547_ _0548_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2237_ _0497_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_68_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2168_ _0440_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2099_ _0383_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xwrapped_sn76489_36 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_14_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1470_ _0903_ _0918_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2522__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2022_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\] _0900_ _0318_ _0319_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_65_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_73_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1806_ _1211_ _1215_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1737_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\] _0972_ _1159_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1668_ _1104_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1599_ _1011_ _1012_ _1041_ _1042_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_68_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2504__A1 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1713__B _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2640_ _0114_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2571_ _0045_ clknet_4_11_0_wb_clk_i net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1522_ _0968_ _0941_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1546__A2 _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1453_ _0900_ _0901_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1384_ tt_um_rejunity_sn76489.chan\[1\].attenuation.in _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2005_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\] _0789_ _0305_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_77_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1584__I _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1528__A2 _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2623_ _0097_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2554_ _0028_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1505_ _0713_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2485_ _0681_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1436_ _0836_ _0883_ _0884_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1367_ _0777_ _0815_ _0781_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1298_ _0746_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1694__A1 _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2650__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2270_ _0520_ _0522_ _0523_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2269__B _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1685__A1 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1985_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\] tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
+ _0285_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2606_ _0080_ clknet_4_11_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2537_ _0011_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2468_ _0626_ tt_um_rejunity_sn76489.latch_control_reg\[0\] _0669_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1419_ _0830_ _0848_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2399_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\] _0617_ _0615_ _0619_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2673__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1770_ _1181_ _1183_ _1184_ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_71_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2546__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2322_ tt_um_rejunity_sn76489.pwm.accumulator\[10\] net25 _0567_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2696__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1370__A3 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2253_ _0842_ _0507_ _0460_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2184_ _0281_ _0449_ _0452_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2018__I _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2181__C _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1968_ net2 _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_55_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1899_ _1091_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1897__A1 _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_49_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2569__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1822_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\] _1051_ _1228_ _1229_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1753_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\] _1172_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1684_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\] _1112_ _1115_ _1117_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2305_ _0550_ _1010_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2236_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\] _0355_ _0494_ _0496_ _0482_
+ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_68_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2167_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\] _0425_ _0437_ _0438_ _0439_
+ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2098_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\] _0362_ _0380_ _0382_ _0377_
+ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_0_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2711__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1587__I _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2359__A2 _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_sn76489_37 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_39_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2021_ _0312_ _0316_ _0317_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_65_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1805_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\] _0993_ _1214_ _1215_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1736_ _1155_ _1156_ _1158_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1667_ net6 _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1598_ _1017_ _1038_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2219_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\] _0468_ _0480_ _0481_ _0482_
+ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_48_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2607__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2570_ _0044_ clknet_4_10_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1521_ _0935_ _0939_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1452_ _0881_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1383_ _0831_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2004_ _0220_ _0304_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2699_ _0173_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1719_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\] _0870_ _1137_ _1144_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_24_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2422__A1 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2622_ _0096_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[2\].attenuation.in
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2553_ _0027_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1504_ _0747_ _0949_ _0950_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_50_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2484_ _0655_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1435_ _0778_ _0838_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1366_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _0815_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1297_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] _0730_ _0746_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_30_Left_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1719__B _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1984_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\] _0289_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
+ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_43_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2605_ _0079_ clknet_4_9_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2536_ _0010_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2467_ _0622_ _1082_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1418_ _0821_ _0865_ _0866_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2398_ _1102_ _0611_ _0618_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1349_ _0737_ _0795_ _0738_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_78_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2321_ _0541_ _0566_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2252_ _0456_ _0509_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2183_ _0365_ _0449_ _0452_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_47_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _0232_ _0273_ _0274_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1898_ tt_um_rejunity_sn76489.clk_counter\[4\] _0219_ tt_um_rejunity_sn76489.clk_counter\[5\]
+ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2640__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2519_ tt_um_rejunity_sn76489.control_noise\[0\]\[0\] _0702_ _0652_ _0704_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1822__B _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2065__A2 _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1821_ _1227_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1752_ _1141_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2663__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1683_ _1102_ _1111_ _1116_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2304_ _0549_ _0551_ _0552_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2235_ _0366_ _0495_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2166_ _1227_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2097_ _0375_ _0379_ _0381_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2056__A2 _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2536__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_sn76489_38 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2686__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2020_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\] _0869_ _0317_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_65_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1804_ _1212_ _1213_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_25_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1735_ _1155_ _1156_ _1157_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_68_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1666_ _1102_ _1088_ _1103_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1597_ _1017_ _1038_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_5_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2559__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2218_ _1098_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2149_ _0424_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_77_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1779__A1 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1520_ _0962_ _0966_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1451_ _0876_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1382_ _0771_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\] _0769_ _0831_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2701__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2003_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\] _0302_ _0304_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_77_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2698_ _0172_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1718_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\] _0870_ _1143_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1649_ _1087_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2110__A1 _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_59_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2621_ _0095_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2552_ _0026_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1503_ _0947_ _0906_ _0747_ _0875_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_50_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2483_ _0627_ _0658_ _0679_ _0656_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1434_ _0815_ _0783_ _0831_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1365_ _0771_ _0780_ _0781_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_37_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1296_ _0732_ _0744_ _0734_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_38_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1825__B _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1735__B _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2398__A1 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1983_ _0288_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_43_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2604_ _0078_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2535_ _0009_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2466_ _0637_ _0661_ _0667_ _0665_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1417_ _0824_ _0864_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2397_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\] _0617_ _0615_ _0618_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1348_ _0736_ _0738_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1279_ _0725_ _0714_ _0727_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_64_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_40_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2320_ tt_um_rejunity_sn76489.pwm.accumulator\[10\] net25 _0565_ _0566_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2251_ _0504_ _0508_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2182_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\] _0441_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
+ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2592__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1966_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\] _0232_ _0235_ _0274_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1897_ _0220_ _0221_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2518_ _0702_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2449_ _0604_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ _1091_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1974__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1751_ _1142_ _1170_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1576__A2 _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1682_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\] _1112_ _1115_ _1116_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2303_ _0549_ _0551_ _0539_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2234_ _0489_ _0493_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2165_ _0433_ _0436_ _0429_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2096_ _0288_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1949_ _0234_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2516__A1 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_sn76489_39 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_65_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2630__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1803_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\] _0998_ _1207_ _1213_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1734_ _1126_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1665_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\] _1089_ _1099_ _1103_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1596_ _1040_ net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2217_ _0474_ _0479_ _0475_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2148_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\] _0384_ _0422_ _0423_ _0419_
+ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1879__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2079_ _0359_ _0363_ _0366_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2503__I _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2653__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1450_ _0890_ _0894_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1381_ _0829_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_78_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2002_ _0301_ _0303_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2195__A2 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2697_ _0171_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1717_ _1141_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2526__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1648_ _1087_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1579_ _1021_ _1023_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2676__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2620_ _0094_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__2549__CLK clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1982__I _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2551_ _0025_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2482_ _1083_ net10 _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2699__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1502_ _0947_ _0906_ _0948_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1433_ _0876_ _0881_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_10_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1364_ _0783_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1295_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\] _0744_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_38_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1603__A1 _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1982_ _0287_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_43_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2603_ _0077_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2534_ _0008_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2465_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] _0662_ _0667_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2396_ _0610_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1416_ _0824_ _0864_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1661__B _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1347_ _0736_ _0795_ _0739_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_48_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1278_ _0726_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2714__CLK clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_40_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__A1 _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2250_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\] _0507_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
+ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_0_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2181_ _0447_ _0353_ _0450_ _0451_ _1141_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_48_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1965_ _0739_ _0272_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_55_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1896_ tt_um_rejunity_sn76489.clk_counter\[4\] _0219_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_11_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2517_ _1109_ _1119_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2448_ _0623_ _0644_ _0653_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2379_ _1075_ _0137_ _0603_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2059__A1 _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1806__A1 _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2416__I _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1750_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\] _1022_ _1169_ _1170_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_80_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1681_ _1098_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2302_ _0550_ _1010_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input9_I io_in_1[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2233_ _0489_ _0493_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2164_ _0433_ _0436_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_68_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2095_ _0375_ _0379_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_51_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1948_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\] _0260_ _0261_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1879_ _1097_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2452__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_sn76489_29 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_47_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2582__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2443__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1802_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\] _0998_ _1212_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1733_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\] _0972_ _1156_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1664_ _1101_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1595_ _1013_ _1039_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2216_ _0474_ _0479_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2147_ _0417_ _0421_ _0381_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2078_ _0365_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1895__I _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1380_ _0785_ _0827_ _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2001_ _0224_ _0302_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2696_ _0170_ clknet_4_3_0_wb_clk_i tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1716_ _1140_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1647_ _1081_ _1082_ _1086_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1578_ _1019_ _1022_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2620__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2550_ _0024_ clknet_4_8_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2481_ _0637_ _0672_ _0678_ _0676_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1501_ _0947_ _0744_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1432_ _0860_ _0878_ _0880_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1363_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\] _0812_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1294_ _0731_ _0735_ _0740_ _0742_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_TAPCELL_ROW_38_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1612__A2 _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2643__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2679_ _0153_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1603__A2 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2419__I _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1981_ _0286_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2666__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1993__I _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2602_ _0076_ clknet_4_12_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2533_ _0007_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2464_ _0634_ _0661_ _0666_ _0665_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2395_ _1096_ _0611_ _0616_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1415_ _0830_ _0848_ _0863_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1346_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\] _0795_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1277_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] _0717_ _0726_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2064__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2539__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2689__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2180_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\] _0448_ _0444_ _0451_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_48_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ tt_um_rejunity_sn76489.control_noise\[0\]\[2\] tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
+ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1895_ _1210_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2516_ _0283_ _1109_ _1119_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2447_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\] _0648_ _0652_ _0653_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2378_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\] _0589_ _0132_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\]
+ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1329_ _0777_ _0768_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XTAP_TAPCELL_ROW_54_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1680_ _1096_ _1111_ _1114_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2704__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2301_ tt_um_rejunity_sn76489.pwm.accumulator\[7\] _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2232_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\] _0492_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
+ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2163_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\] _0426_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
+ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2094_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\] _0373_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
+ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_51_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1947_ _0237_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1878_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\] _1052_ _0208_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2452__A2 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2201__B _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1801_ _1210_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_13_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1732_ _1150_ _0923_ _1154_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1663_ net5 _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_80_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1594_ _1017_ _1038_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_5_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_37_Left_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2215_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\] _0478_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
+ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2146_ _0417_ _0421_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2077_ _0286_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_55_Left_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_64_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_73_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2000_ tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\] _0299_ _0295_ _0302_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_18_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1715_ _1130_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2695_ _0169_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1646_ _1083_ _1085_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1577_ _1020_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2129_ _0315_ _0408_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2572__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2016__B _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2343__A1 _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2480_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] _0673_ _0678_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1500_ _0732_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1431_ _0720_ _0879_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1362_ _0808_ _0810_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2595__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1293_ _0741_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_38_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2678_ _0152_ clknet_4_6_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1629_ _1043_ _1061_ _1071_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1980_ _0285_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2601_ _0075_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2532_ _0006_ clknet_4_4_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2463_ _0947_ _0662_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2394_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\] _0612_ _0615_ _0616_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1414_ _0855_ _0862_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1345_ _0725_ _0714_ _0792_ _0793_ _0716_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_64_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1276_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\] _0724_ _0717_ _0725_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_78_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2610__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__1521__A2 _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1963_ _0270_ _0271_ _0235_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_50_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1894_ _0215_ _0218_ _0219_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_70_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2515_ _0701_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2446_ _1091_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2377_ _0602_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1328_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\] _0777_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1259_ tt_um_rejunity_sn76489.chan\[2\].attenuation.in _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_38_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2656__CLK clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2300_ _0547_ _0548_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2231_ _0478_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2162_ _0435_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2093_ _0378_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1946_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\] _0252_ _0259_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2529__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1877_ _0194_ _0207_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2679__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2429_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\] _0635_ _0638_ _0641_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_67_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ _1140_ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_13_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1731_ _1149_ _1153_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1662_ _1096_ _1088_ _1100_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1593_ _1024_ _1037_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2214_ _0465_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2145_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\] _0413_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
+ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2131__A2 _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2076_ _0359_ _0363_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1929_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\] _0238_ _0247_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2189__A2 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1607__I _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1714_ _1137_ _1138_ _1139_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2694_ _0168_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1645_ net11 _1084_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_67_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1576_ _1019_ _1020_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_67_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2717__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2128_ _0402_ _0407_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2059_ _0315_ _0349_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_24_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1606__A1 _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1430_ _0711_ _0709_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1361_ _0751_ _0806_ _0809_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1292_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] _0729_ _0741_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_53_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2677_ _0151_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1628_ _1044_ _1060_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1559_ tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] _0735_ _1005_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2078__I _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1620__I _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2252__A1 _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2004__A1 _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ _0074_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2531_ _0005_ clknet_4_5_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2562__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2462_ _0632_ _0661_ _0664_ _0665_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_48_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2393_ _0614_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1413_ _0856_ _0857_ _0859_ _0861_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1344_ _0720_ _0725_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1275_ _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1818__A1 _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2491__A1 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output16_I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2585__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1962_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\] _0237_ _0271_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1893_ tt_um_rejunity_sn76489.clk_counter\[3\] _0217_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_70_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2514_ tt_um_rejunity_sn76489.latch_control_reg\[2\] _0698_ _1086_ _1228_ _0701_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2445_ _0620_ _0644_ _0651_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2130__B _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2376_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\] _1079_ _0590_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\]
+ _0581_ net25 _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1327_ _0773_ _0774_ _0775_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2464__A1 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2091__I _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2230_ _0491_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2600__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2161_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\] _0425_ _0433_ _0434_ _0419_
+ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2092_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\] _0362_ _0375_ _0376_ _0377_
+ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_61_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2125__B _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1945_ _0257_ _0258_ _0251_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1876_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\] _1052_ _0206_ _0207_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_71_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2428_ _0620_ _0630_ _0640_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2359_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\] _0000_ _0132_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\]
+ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2623__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2428__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1730_ _1150_ _0923_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1661_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\] _1089_ _1099_ _1100_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1592_ _1026_ _1027_ _1036_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2213_ _0477_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input7_I io_in_1[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2144_ _0420_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2075_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\] _0358_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
+ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_64_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1678__C _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1928_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\] _0241_ _0246_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2646__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1859_ _1257_ _1258_ _1238_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1633__A2 _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2669__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1713_ _1137_ _1138_ _1127_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2693_ _0167_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1644_ net10 _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1575_ _0877_ _0727_ _0860_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_67_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2127_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\] _0406_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
+ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2058_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\] _1063_ _0348_ _0349_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_24_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1360_ _0765_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1291_ _0736_ _0737_ _0739_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_46_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2676_ _0150_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1627_ _1067_ _1069_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1558_ _0859_ _0793_ _1003_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1489_ _0813_ _0834_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_37_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2261__A2 _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2707__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2530_ _0004_ clknet_4_1_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2461_ _1092_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1792__B _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1412_ _0721_ _0860_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2392_ _1097_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1343_ _0710_ _0723_ _0718_ _0720_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XPHY_EDGE_ROW_79_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1274_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\] _0723_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2243__A2 _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2659_ _0133_ clknet_4_13_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2482__A2 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1961_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\] _0263_ _0270_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ tt_um_rejunity_sn76489.clk_counter\[3\] _0217_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2513_ _0623_ _0698_ _0700_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2444_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\] _0648_ _0646_ _0651_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2375_ _0601_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1326_ tt_um_rejunity_sn76489.chan\[1\].attenuation.in _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_75_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1451__I _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2552__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2391__A1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2160_ _0428_ _0432_ _0429_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2091_ _1227_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1944_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\] _0249_ _0258_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1875_ _0201_ _0204_ _0205_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_3_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2427_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\] _0635_ _0638_ _0640_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2358_ _0591_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1309_ tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\] _0758_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2575__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2289_ _0537_ _0538_ _0539_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_67_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ _1098_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1591_ _1034_ _1035_ _0995_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2598__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2212_ tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\] _0468_ _0474_ _0476_ _0439_
+ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2143_ tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\] _0384_ _0417_ _0418_ _0419_
+ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2074_ _0361_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_64_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ _0244_ _0245_ _0240_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1858_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\] _0997_ _1258_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1789_ _1196_ _1032_ _1200_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_24_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Left_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_42_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_78_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2692_ _0166_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1712_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\] _0870_ _1138_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1643_ net9 _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1574_ _1018_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_60_Left_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2126_ _0287_ _0389_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_76_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2057_ _0346_ _0347_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2613__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1290_ _0738_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2636__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2675_ _0149_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1626_ _1053_ _1068_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1557_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] _0719_ _1003_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1488_ _0772_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1297__A1 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2109_ _0386_ _0390_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1524__A2 _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2659__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2460_ _0733_ _0662_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1411_ _0710_ _0711_ _0713_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2391_ _0605_ _0611_ _0613_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1342_ _0787_ _0790_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1273_ _0709_ _0714_ _0719_ _0721_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_78_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2658_ _0132_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2589_ _0063_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1609_ _1051_ _1052_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1960_ _0268_ _0269_ _0262_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1891_ _0215_ _0216_ _0217_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1433__A1 _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1984__A2 _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2512_ _0606_ _1085_ _0652_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2443_ _0637_ _0643_ _0650_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2374_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\] _0596_ _0590_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\]
+ _0597_ net24 _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1325_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\] _0774_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_75_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1975__A2 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2512__B _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1642__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2090_ _0370_ _0374_ _0366_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__1798__B _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1943_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\] _0252_ _0257_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1874_ _0203_ _1026_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2426_ _0637_ _0629_ _0639_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2357_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\] _0589_ _0521_ _0585_
+ _0590_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\] _0591_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_2288_ _0209_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1308_ _0754_ _0756_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_67_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1645__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1590_ _0999_ _0992_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2211_ _0470_ _0473_ _0475_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2142_ _1227_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2073_ _0287_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1926_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\] _0238_ _0245_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1857_ _1255_ _1256_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1547__I _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1788_ _1195_ _1199_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2542__CLK clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2409_ tt_um_rejunity_sn76489.latch_control_reg\[1\] _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2692__CLK clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1866__A1 _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2691_ _0165_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1711_ _1133_ _1135_ _1136_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1642_ net7 _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2565__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1573_ _0852_ _0873_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_67_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2125_ _0402_ _0405_ _0213_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2056_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\] _1018_ _0343_ _0347_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1909_ _0230_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2588__CLK clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2504__C _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2674_ _0148_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1625_ _1050_ _1058_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1556_ _0996_ _1001_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1487_ _0759_ _0806_ _0934_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2108_ _0386_ _0390_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2246__A1 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2039_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\] _0973_ _0333_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_80_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_64_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1410_ _0856_ _0857_ _0858_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2390_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\] _0612_ _0539_ _0613_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2603__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1341_ _0788_ _0789_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1272_ _0720_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2400__A1 _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2657_ _0131_ clknet_4_15_0_wb_clk_i net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1608_ _1049_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2588_ _0062_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1539_ _0983_ _0984_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2626__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_48_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1890_ _0212_ tt_um_rejunity_sn76489.clk_counter\[1\] tt_um_rejunity_sn76489.clk_counter\[2\]
+ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_55_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2511_ _0620_ _0698_ _0699_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2442_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\] _0648_ _0646_ _0650_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2373_ _0600_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1324_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _0773_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_75_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1994__B _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2649__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2709_ _0183_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_42_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1942_ _0255_ _0256_ _0251_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1873_ _0203_ _1026_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2425_ tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\] _0635_ _0638_ _0639_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2356_ _0574_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1307_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2287_ tt_um_rejunity_sn76489.pwm.accumulator\[5\] net20 _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1989__B _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2210_ _0365_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2141_ _0414_ _0416_ _0381_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2072_ _0354_ _0360_ _0213_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1627__A2 _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1925_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\] _0241_ _0244_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2052__A2 _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1856_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\] _1028_ _1252_ _1256_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1787_ _1196_ _1032_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2408_ _0623_ _0612_ _0625_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2339_ tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\] _0578_ _0579_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2062__C _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2253__B _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2690_ _0164_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1710_ tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\] _0822_ _1136_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1641_ net8 _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1572_ _1002_ _1008_ _1016_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input5_I io_in_1[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2124_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\] _0403_ _0404_ _0405_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2055_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\] _1018_ _0346_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1908_ tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
+ _0229_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_32_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1839_ _1240_ _1241_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1775__A1 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2248__B _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2532__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2682__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2673_ _0147_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1624_ _1065_ _1066_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1555_ _0967_ _0969_ _1000_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2191__A1 _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1486_ _0809_ _0841_ _0845_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2107_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\] _0389_ tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
+ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_37_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1997__B _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2038_ tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\] _0973_ _0332_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_80_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_20_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2555__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_39_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2173__A1 _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1340_ _0743_ _0748_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1271_ tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\] _0708_ _0720_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_80_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1987__A1 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2656_ _0130_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.pwm.accumulator\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1607_ _1048_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2587_ _0061_ clknet_4_7_0_wb_clk_i tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1538_ _0957_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2578__CLK clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1469_ _0908_ _0917_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1902__A1 _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__I _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2510_ _0607_ _0698_ _0652_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2441_ _0634_ _0643_ _0649_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2372_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\] _0596_ _0590_ tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\]
+ _0597_ net23 _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1323_ tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\] _0771_ _0769_ _0772_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_75_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2708_ _0182_ clknet_4_2_0_wb_clk_i tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2137__A1 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2639_ _0113_ clknet_4_0_0_wb_clk_i tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_2_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2100__I _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2256__B _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1941_ tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\] _0249_ _0256_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1872_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\] _0203_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_71_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2424_ _0614_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2355_ _1079_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1306_ tt_um_rejunity_sn76489.chan\[0\].attenuation.in _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2286_ _0536_ _0534_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2616__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2639__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _0414_ _0416_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2071_ _0355_ _0359_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1924_ _0242_ _0243_ _0240_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1855_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\] _1028_ _1255_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1786_ _1195_ _1197_ _1198_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2407_ tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\] _0617_ _0624_ _0625_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2338_ _0573_ _0577_ _0578_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2269_ _0520_ _0522_ _0460_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1640_ tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\] _1080_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1571_ _1014_ _1015_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1664__I _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2123_ _0281_ _0398_ _0401_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_49_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2054_ _0343_ _0344_ _0345_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1907_ _0228_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1838_ tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\] _0892_ _1236_ _1241_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1769_ tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\] _0818_ _1184_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1574__I _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1659__I _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2672_ _0146_ clknet_4_15_0_wb_clk_i tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1623_ _1047_ _1059_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1554_ _0999_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1485_ _0829_ _0912_ _0911_ _0915_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
.ends

