magic
tech gf180mcuD
magscale 1 5
timestamp 1699038623
<< obsm1 >>
rect 672 1471 59304 58673
<< metal2 >>
rect 2464 59600 2520 60000
rect 3024 59600 3080 60000
rect 3584 59600 3640 60000
rect 4144 59600 4200 60000
rect 4704 59600 4760 60000
rect 5264 59600 5320 60000
rect 5824 59600 5880 60000
rect 6384 59600 6440 60000
rect 6944 59600 7000 60000
rect 7504 59600 7560 60000
rect 8064 59600 8120 60000
rect 8624 59600 8680 60000
rect 9184 59600 9240 60000
rect 9744 59600 9800 60000
rect 10304 59600 10360 60000
rect 10864 59600 10920 60000
rect 11424 59600 11480 60000
rect 11984 59600 12040 60000
rect 12544 59600 12600 60000
rect 13104 59600 13160 60000
rect 13664 59600 13720 60000
rect 14224 59600 14280 60000
rect 14784 59600 14840 60000
rect 15344 59600 15400 60000
rect 15904 59600 15960 60000
rect 16464 59600 16520 60000
rect 17024 59600 17080 60000
rect 17584 59600 17640 60000
rect 18144 59600 18200 60000
rect 18704 59600 18760 60000
rect 19264 59600 19320 60000
rect 19824 59600 19880 60000
rect 20384 59600 20440 60000
rect 20944 59600 21000 60000
rect 21504 59600 21560 60000
rect 22064 59600 22120 60000
rect 22624 59600 22680 60000
rect 23184 59600 23240 60000
rect 23744 59600 23800 60000
rect 24304 59600 24360 60000
rect 24864 59600 24920 60000
rect 25424 59600 25480 60000
rect 25984 59600 26040 60000
rect 26544 59600 26600 60000
rect 27104 59600 27160 60000
rect 27664 59600 27720 60000
rect 28224 59600 28280 60000
rect 28784 59600 28840 60000
rect 29344 59600 29400 60000
rect 29904 59600 29960 60000
rect 30464 59600 30520 60000
rect 31024 59600 31080 60000
rect 31584 59600 31640 60000
rect 32144 59600 32200 60000
rect 32704 59600 32760 60000
rect 33264 59600 33320 60000
rect 33824 59600 33880 60000
rect 34384 59600 34440 60000
rect 34944 59600 35000 60000
rect 35504 59600 35560 60000
rect 36064 59600 36120 60000
rect 36624 59600 36680 60000
rect 37184 59600 37240 60000
rect 37744 59600 37800 60000
rect 38304 59600 38360 60000
rect 38864 59600 38920 60000
rect 39424 59600 39480 60000
rect 39984 59600 40040 60000
rect 40544 59600 40600 60000
rect 41104 59600 41160 60000
rect 41664 59600 41720 60000
rect 42224 59600 42280 60000
rect 42784 59600 42840 60000
rect 43344 59600 43400 60000
rect 43904 59600 43960 60000
rect 44464 59600 44520 60000
rect 45024 59600 45080 60000
rect 45584 59600 45640 60000
rect 46144 59600 46200 60000
rect 46704 59600 46760 60000
rect 47264 59600 47320 60000
rect 47824 59600 47880 60000
rect 48384 59600 48440 60000
rect 48944 59600 49000 60000
rect 49504 59600 49560 60000
rect 50064 59600 50120 60000
rect 50624 59600 50680 60000
rect 51184 59600 51240 60000
rect 51744 59600 51800 60000
rect 52304 59600 52360 60000
rect 52864 59600 52920 60000
rect 53424 59600 53480 60000
rect 53984 59600 54040 60000
rect 54544 59600 54600 60000
rect 55104 59600 55160 60000
rect 55664 59600 55720 60000
rect 56224 59600 56280 60000
rect 56784 59600 56840 60000
rect 57344 59600 57400 60000
rect 112 0 168 400
rect 560 0 616 400
rect 1008 0 1064 400
rect 1456 0 1512 400
rect 1904 0 1960 400
rect 2352 0 2408 400
rect 2800 0 2856 400
rect 3248 0 3304 400
rect 3696 0 3752 400
rect 4144 0 4200 400
rect 4592 0 4648 400
rect 5040 0 5096 400
rect 5488 0 5544 400
rect 5936 0 5992 400
rect 6384 0 6440 400
rect 6832 0 6888 400
rect 7280 0 7336 400
rect 7728 0 7784 400
rect 8176 0 8232 400
rect 8624 0 8680 400
rect 9072 0 9128 400
rect 9520 0 9576 400
rect 9968 0 10024 400
rect 10416 0 10472 400
rect 10864 0 10920 400
rect 11312 0 11368 400
rect 11760 0 11816 400
rect 12208 0 12264 400
rect 12656 0 12712 400
rect 13104 0 13160 400
rect 13552 0 13608 400
rect 14000 0 14056 400
rect 14448 0 14504 400
rect 14896 0 14952 400
rect 15344 0 15400 400
rect 15792 0 15848 400
rect 16240 0 16296 400
rect 16688 0 16744 400
rect 17136 0 17192 400
rect 17584 0 17640 400
rect 18032 0 18088 400
rect 18480 0 18536 400
rect 18928 0 18984 400
rect 19376 0 19432 400
rect 19824 0 19880 400
rect 20272 0 20328 400
rect 20720 0 20776 400
rect 21168 0 21224 400
rect 21616 0 21672 400
rect 22064 0 22120 400
rect 22512 0 22568 400
rect 22960 0 23016 400
rect 23408 0 23464 400
rect 23856 0 23912 400
rect 24304 0 24360 400
rect 24752 0 24808 400
rect 25200 0 25256 400
rect 25648 0 25704 400
rect 26096 0 26152 400
rect 26544 0 26600 400
rect 26992 0 27048 400
rect 27440 0 27496 400
rect 27888 0 27944 400
rect 28336 0 28392 400
rect 28784 0 28840 400
rect 29232 0 29288 400
rect 29680 0 29736 400
rect 30128 0 30184 400
rect 30576 0 30632 400
rect 31024 0 31080 400
rect 31472 0 31528 400
rect 31920 0 31976 400
rect 32368 0 32424 400
rect 32816 0 32872 400
rect 33264 0 33320 400
rect 33712 0 33768 400
rect 34160 0 34216 400
rect 34608 0 34664 400
rect 35056 0 35112 400
rect 35504 0 35560 400
rect 35952 0 36008 400
rect 36400 0 36456 400
rect 36848 0 36904 400
rect 37296 0 37352 400
rect 37744 0 37800 400
rect 38192 0 38248 400
rect 38640 0 38696 400
rect 39088 0 39144 400
rect 39536 0 39592 400
rect 39984 0 40040 400
rect 40432 0 40488 400
rect 40880 0 40936 400
rect 41328 0 41384 400
rect 41776 0 41832 400
rect 42224 0 42280 400
rect 42672 0 42728 400
rect 43120 0 43176 400
rect 43568 0 43624 400
rect 44016 0 44072 400
rect 44464 0 44520 400
rect 44912 0 44968 400
rect 45360 0 45416 400
rect 45808 0 45864 400
rect 46256 0 46312 400
rect 46704 0 46760 400
rect 47152 0 47208 400
rect 47600 0 47656 400
rect 48048 0 48104 400
rect 48496 0 48552 400
rect 48944 0 49000 400
rect 49392 0 49448 400
rect 49840 0 49896 400
rect 50288 0 50344 400
rect 50736 0 50792 400
rect 51184 0 51240 400
rect 51632 0 51688 400
rect 52080 0 52136 400
rect 52528 0 52584 400
rect 52976 0 53032 400
rect 53424 0 53480 400
rect 53872 0 53928 400
rect 54320 0 54376 400
rect 54768 0 54824 400
rect 55216 0 55272 400
rect 55664 0 55720 400
rect 56112 0 56168 400
rect 56560 0 56616 400
rect 57008 0 57064 400
rect 57456 0 57512 400
rect 57904 0 57960 400
rect 58352 0 58408 400
rect 58800 0 58856 400
rect 59248 0 59304 400
rect 59696 0 59752 400
<< obsm2 >>
rect 126 59570 2434 59682
rect 2550 59570 2994 59682
rect 3110 59570 3554 59682
rect 3670 59570 4114 59682
rect 4230 59570 4674 59682
rect 4790 59570 5234 59682
rect 5350 59570 5794 59682
rect 5910 59570 6354 59682
rect 6470 59570 6914 59682
rect 7030 59570 7474 59682
rect 7590 59570 8034 59682
rect 8150 59570 8594 59682
rect 8710 59570 9154 59682
rect 9270 59570 9714 59682
rect 9830 59570 10274 59682
rect 10390 59570 10834 59682
rect 10950 59570 11394 59682
rect 11510 59570 11954 59682
rect 12070 59570 12514 59682
rect 12630 59570 13074 59682
rect 13190 59570 13634 59682
rect 13750 59570 14194 59682
rect 14310 59570 14754 59682
rect 14870 59570 15314 59682
rect 15430 59570 15874 59682
rect 15990 59570 16434 59682
rect 16550 59570 16994 59682
rect 17110 59570 17554 59682
rect 17670 59570 18114 59682
rect 18230 59570 18674 59682
rect 18790 59570 19234 59682
rect 19350 59570 19794 59682
rect 19910 59570 20354 59682
rect 20470 59570 20914 59682
rect 21030 59570 21474 59682
rect 21590 59570 22034 59682
rect 22150 59570 22594 59682
rect 22710 59570 23154 59682
rect 23270 59570 23714 59682
rect 23830 59570 24274 59682
rect 24390 59570 24834 59682
rect 24950 59570 25394 59682
rect 25510 59570 25954 59682
rect 26070 59570 26514 59682
rect 26630 59570 27074 59682
rect 27190 59570 27634 59682
rect 27750 59570 28194 59682
rect 28310 59570 28754 59682
rect 28870 59570 29314 59682
rect 29430 59570 29874 59682
rect 29990 59570 30434 59682
rect 30550 59570 30994 59682
rect 31110 59570 31554 59682
rect 31670 59570 32114 59682
rect 32230 59570 32674 59682
rect 32790 59570 33234 59682
rect 33350 59570 33794 59682
rect 33910 59570 34354 59682
rect 34470 59570 34914 59682
rect 35030 59570 35474 59682
rect 35590 59570 36034 59682
rect 36150 59570 36594 59682
rect 36710 59570 37154 59682
rect 37270 59570 37714 59682
rect 37830 59570 38274 59682
rect 38390 59570 38834 59682
rect 38950 59570 39394 59682
rect 39510 59570 39954 59682
rect 40070 59570 40514 59682
rect 40630 59570 41074 59682
rect 41190 59570 41634 59682
rect 41750 59570 42194 59682
rect 42310 59570 42754 59682
rect 42870 59570 43314 59682
rect 43430 59570 43874 59682
rect 43990 59570 44434 59682
rect 44550 59570 44994 59682
rect 45110 59570 45554 59682
rect 45670 59570 46114 59682
rect 46230 59570 46674 59682
rect 46790 59570 47234 59682
rect 47350 59570 47794 59682
rect 47910 59570 48354 59682
rect 48470 59570 48914 59682
rect 49030 59570 49474 59682
rect 49590 59570 50034 59682
rect 50150 59570 50594 59682
rect 50710 59570 51154 59682
rect 51270 59570 51714 59682
rect 51830 59570 52274 59682
rect 52390 59570 52834 59682
rect 52950 59570 53394 59682
rect 53510 59570 53954 59682
rect 54070 59570 54514 59682
rect 54630 59570 55074 59682
rect 55190 59570 55634 59682
rect 55750 59570 56194 59682
rect 56310 59570 56754 59682
rect 56870 59570 57314 59682
rect 57430 59570 59738 59682
rect 126 430 59738 59570
rect 198 350 530 430
rect 646 350 978 430
rect 1094 350 1426 430
rect 1542 350 1874 430
rect 1990 350 2322 430
rect 2438 350 2770 430
rect 2886 350 3218 430
rect 3334 350 3666 430
rect 3782 350 4114 430
rect 4230 350 4562 430
rect 4678 350 5010 430
rect 5126 350 5458 430
rect 5574 350 5906 430
rect 6022 350 6354 430
rect 6470 350 6802 430
rect 6918 350 7250 430
rect 7366 350 7698 430
rect 7814 350 8146 430
rect 8262 350 8594 430
rect 8710 350 9042 430
rect 9158 350 9490 430
rect 9606 350 9938 430
rect 10054 350 10386 430
rect 10502 350 10834 430
rect 10950 350 11282 430
rect 11398 350 11730 430
rect 11846 350 12178 430
rect 12294 350 12626 430
rect 12742 350 13074 430
rect 13190 350 13522 430
rect 13638 350 13970 430
rect 14086 350 14418 430
rect 14534 350 14866 430
rect 14982 350 15314 430
rect 15430 350 15762 430
rect 15878 350 16210 430
rect 16326 350 16658 430
rect 16774 350 17106 430
rect 17222 350 17554 430
rect 17670 350 18002 430
rect 18118 350 18450 430
rect 18566 350 18898 430
rect 19014 350 19346 430
rect 19462 350 19794 430
rect 19910 350 20242 430
rect 20358 350 20690 430
rect 20806 350 21138 430
rect 21254 350 21586 430
rect 21702 350 22034 430
rect 22150 350 22482 430
rect 22598 350 22930 430
rect 23046 350 23378 430
rect 23494 350 23826 430
rect 23942 350 24274 430
rect 24390 350 24722 430
rect 24838 350 25170 430
rect 25286 350 25618 430
rect 25734 350 26066 430
rect 26182 350 26514 430
rect 26630 350 26962 430
rect 27078 350 27410 430
rect 27526 350 27858 430
rect 27974 350 28306 430
rect 28422 350 28754 430
rect 28870 350 29202 430
rect 29318 350 29650 430
rect 29766 350 30098 430
rect 30214 350 30546 430
rect 30662 350 30994 430
rect 31110 350 31442 430
rect 31558 350 31890 430
rect 32006 350 32338 430
rect 32454 350 32786 430
rect 32902 350 33234 430
rect 33350 350 33682 430
rect 33798 350 34130 430
rect 34246 350 34578 430
rect 34694 350 35026 430
rect 35142 350 35474 430
rect 35590 350 35922 430
rect 36038 350 36370 430
rect 36486 350 36818 430
rect 36934 350 37266 430
rect 37382 350 37714 430
rect 37830 350 38162 430
rect 38278 350 38610 430
rect 38726 350 39058 430
rect 39174 350 39506 430
rect 39622 350 39954 430
rect 40070 350 40402 430
rect 40518 350 40850 430
rect 40966 350 41298 430
rect 41414 350 41746 430
rect 41862 350 42194 430
rect 42310 350 42642 430
rect 42758 350 43090 430
rect 43206 350 43538 430
rect 43654 350 43986 430
rect 44102 350 44434 430
rect 44550 350 44882 430
rect 44998 350 45330 430
rect 45446 350 45778 430
rect 45894 350 46226 430
rect 46342 350 46674 430
rect 46790 350 47122 430
rect 47238 350 47570 430
rect 47686 350 48018 430
rect 48134 350 48466 430
rect 48582 350 48914 430
rect 49030 350 49362 430
rect 49478 350 49810 430
rect 49926 350 50258 430
rect 50374 350 50706 430
rect 50822 350 51154 430
rect 51270 350 51602 430
rect 51718 350 52050 430
rect 52166 350 52498 430
rect 52614 350 52946 430
rect 53062 350 53394 430
rect 53510 350 53842 430
rect 53958 350 54290 430
rect 54406 350 54738 430
rect 54854 350 55186 430
rect 55302 350 55634 430
rect 55750 350 56082 430
rect 56198 350 56530 430
rect 56646 350 56978 430
rect 57094 350 57426 430
rect 57542 350 57874 430
rect 57990 350 58322 430
rect 58438 350 58770 430
rect 58886 350 59218 430
rect 59334 350 59666 430
<< metal3 >>
rect 0 56000 400 56056
rect 59600 55888 60000 55944
rect 0 55440 400 55496
rect 59600 55440 60000 55496
rect 59600 54992 60000 55048
rect 0 54880 400 54936
rect 59600 54544 60000 54600
rect 0 54320 400 54376
rect 59600 54096 60000 54152
rect 0 53760 400 53816
rect 59600 53648 60000 53704
rect 0 53200 400 53256
rect 59600 53200 60000 53256
rect 59600 52752 60000 52808
rect 0 52640 400 52696
rect 59600 52304 60000 52360
rect 0 52080 400 52136
rect 59600 51856 60000 51912
rect 0 51520 400 51576
rect 59600 51408 60000 51464
rect 0 50960 400 51016
rect 59600 50960 60000 51016
rect 59600 50512 60000 50568
rect 0 50400 400 50456
rect 59600 50064 60000 50120
rect 0 49840 400 49896
rect 59600 49616 60000 49672
rect 0 49280 400 49336
rect 59600 49168 60000 49224
rect 0 48720 400 48776
rect 59600 48720 60000 48776
rect 59600 48272 60000 48328
rect 0 48160 400 48216
rect 59600 47824 60000 47880
rect 0 47600 400 47656
rect 59600 47376 60000 47432
rect 0 47040 400 47096
rect 59600 46928 60000 46984
rect 0 46480 400 46536
rect 59600 46480 60000 46536
rect 59600 46032 60000 46088
rect 0 45920 400 45976
rect 59600 45584 60000 45640
rect 0 45360 400 45416
rect 59600 45136 60000 45192
rect 0 44800 400 44856
rect 59600 44688 60000 44744
rect 0 44240 400 44296
rect 59600 44240 60000 44296
rect 59600 43792 60000 43848
rect 0 43680 400 43736
rect 59600 43344 60000 43400
rect 0 43120 400 43176
rect 59600 42896 60000 42952
rect 0 42560 400 42616
rect 59600 42448 60000 42504
rect 0 42000 400 42056
rect 59600 42000 60000 42056
rect 59600 41552 60000 41608
rect 0 41440 400 41496
rect 59600 41104 60000 41160
rect 0 40880 400 40936
rect 59600 40656 60000 40712
rect 0 40320 400 40376
rect 59600 40208 60000 40264
rect 0 39760 400 39816
rect 59600 39760 60000 39816
rect 59600 39312 60000 39368
rect 0 39200 400 39256
rect 59600 38864 60000 38920
rect 0 38640 400 38696
rect 59600 38416 60000 38472
rect 0 38080 400 38136
rect 59600 37968 60000 38024
rect 0 37520 400 37576
rect 59600 37520 60000 37576
rect 59600 37072 60000 37128
rect 0 36960 400 37016
rect 59600 36624 60000 36680
rect 0 36400 400 36456
rect 59600 36176 60000 36232
rect 0 35840 400 35896
rect 59600 35728 60000 35784
rect 0 35280 400 35336
rect 59600 35280 60000 35336
rect 59600 34832 60000 34888
rect 0 34720 400 34776
rect 59600 34384 60000 34440
rect 0 34160 400 34216
rect 59600 33936 60000 33992
rect 0 33600 400 33656
rect 59600 33488 60000 33544
rect 0 33040 400 33096
rect 59600 33040 60000 33096
rect 59600 32592 60000 32648
rect 0 32480 400 32536
rect 59600 32144 60000 32200
rect 0 31920 400 31976
rect 59600 31696 60000 31752
rect 0 31360 400 31416
rect 59600 31248 60000 31304
rect 0 30800 400 30856
rect 59600 30800 60000 30856
rect 59600 30352 60000 30408
rect 0 30240 400 30296
rect 59600 29904 60000 29960
rect 0 29680 400 29736
rect 59600 29456 60000 29512
rect 0 29120 400 29176
rect 59600 29008 60000 29064
rect 0 28560 400 28616
rect 59600 28560 60000 28616
rect 59600 28112 60000 28168
rect 0 28000 400 28056
rect 59600 27664 60000 27720
rect 0 27440 400 27496
rect 59600 27216 60000 27272
rect 0 26880 400 26936
rect 59600 26768 60000 26824
rect 0 26320 400 26376
rect 59600 26320 60000 26376
rect 59600 25872 60000 25928
rect 0 25760 400 25816
rect 59600 25424 60000 25480
rect 0 25200 400 25256
rect 59600 24976 60000 25032
rect 0 24640 400 24696
rect 59600 24528 60000 24584
rect 0 24080 400 24136
rect 59600 24080 60000 24136
rect 59600 23632 60000 23688
rect 0 23520 400 23576
rect 59600 23184 60000 23240
rect 0 22960 400 23016
rect 59600 22736 60000 22792
rect 0 22400 400 22456
rect 59600 22288 60000 22344
rect 0 21840 400 21896
rect 59600 21840 60000 21896
rect 59600 21392 60000 21448
rect 0 21280 400 21336
rect 59600 20944 60000 21000
rect 0 20720 400 20776
rect 59600 20496 60000 20552
rect 0 20160 400 20216
rect 59600 20048 60000 20104
rect 0 19600 400 19656
rect 59600 19600 60000 19656
rect 59600 19152 60000 19208
rect 0 19040 400 19096
rect 59600 18704 60000 18760
rect 0 18480 400 18536
rect 59600 18256 60000 18312
rect 0 17920 400 17976
rect 59600 17808 60000 17864
rect 0 17360 400 17416
rect 59600 17360 60000 17416
rect 59600 16912 60000 16968
rect 0 16800 400 16856
rect 59600 16464 60000 16520
rect 0 16240 400 16296
rect 59600 16016 60000 16072
rect 0 15680 400 15736
rect 59600 15568 60000 15624
rect 0 15120 400 15176
rect 59600 15120 60000 15176
rect 59600 14672 60000 14728
rect 0 14560 400 14616
rect 59600 14224 60000 14280
rect 0 14000 400 14056
rect 59600 13776 60000 13832
rect 0 13440 400 13496
rect 59600 13328 60000 13384
rect 0 12880 400 12936
rect 59600 12880 60000 12936
rect 59600 12432 60000 12488
rect 0 12320 400 12376
rect 59600 11984 60000 12040
rect 0 11760 400 11816
rect 59600 11536 60000 11592
rect 0 11200 400 11256
rect 59600 11088 60000 11144
rect 0 10640 400 10696
rect 59600 10640 60000 10696
rect 59600 10192 60000 10248
rect 0 10080 400 10136
rect 59600 9744 60000 9800
rect 0 9520 400 9576
rect 59600 9296 60000 9352
rect 0 8960 400 9016
rect 59600 8848 60000 8904
rect 0 8400 400 8456
rect 59600 8400 60000 8456
rect 59600 7952 60000 8008
rect 0 7840 400 7896
rect 59600 7504 60000 7560
rect 0 7280 400 7336
rect 59600 7056 60000 7112
rect 0 6720 400 6776
rect 59600 6608 60000 6664
rect 0 6160 400 6216
rect 59600 6160 60000 6216
rect 59600 5712 60000 5768
rect 0 5600 400 5656
rect 59600 5264 60000 5320
rect 0 5040 400 5096
rect 59600 4816 60000 4872
rect 0 4480 400 4536
rect 59600 4368 60000 4424
rect 0 3920 400 3976
rect 59600 3920 60000 3976
<< obsm3 >>
rect 121 56086 59743 58786
rect 430 55974 59743 56086
rect 430 55970 59570 55974
rect 121 55858 59570 55970
rect 121 55526 59743 55858
rect 430 55410 59570 55526
rect 121 55078 59743 55410
rect 121 54966 59570 55078
rect 430 54962 59570 54966
rect 430 54850 59743 54962
rect 121 54630 59743 54850
rect 121 54514 59570 54630
rect 121 54406 59743 54514
rect 430 54290 59743 54406
rect 121 54182 59743 54290
rect 121 54066 59570 54182
rect 121 53846 59743 54066
rect 430 53734 59743 53846
rect 430 53730 59570 53734
rect 121 53618 59570 53730
rect 121 53286 59743 53618
rect 430 53170 59570 53286
rect 121 52838 59743 53170
rect 121 52726 59570 52838
rect 430 52722 59570 52726
rect 430 52610 59743 52722
rect 121 52390 59743 52610
rect 121 52274 59570 52390
rect 121 52166 59743 52274
rect 430 52050 59743 52166
rect 121 51942 59743 52050
rect 121 51826 59570 51942
rect 121 51606 59743 51826
rect 430 51494 59743 51606
rect 430 51490 59570 51494
rect 121 51378 59570 51490
rect 121 51046 59743 51378
rect 430 50930 59570 51046
rect 121 50598 59743 50930
rect 121 50486 59570 50598
rect 430 50482 59570 50486
rect 430 50370 59743 50482
rect 121 50150 59743 50370
rect 121 50034 59570 50150
rect 121 49926 59743 50034
rect 430 49810 59743 49926
rect 121 49702 59743 49810
rect 121 49586 59570 49702
rect 121 49366 59743 49586
rect 430 49254 59743 49366
rect 430 49250 59570 49254
rect 121 49138 59570 49250
rect 121 48806 59743 49138
rect 430 48690 59570 48806
rect 121 48358 59743 48690
rect 121 48246 59570 48358
rect 430 48242 59570 48246
rect 430 48130 59743 48242
rect 121 47910 59743 48130
rect 121 47794 59570 47910
rect 121 47686 59743 47794
rect 430 47570 59743 47686
rect 121 47462 59743 47570
rect 121 47346 59570 47462
rect 121 47126 59743 47346
rect 430 47014 59743 47126
rect 430 47010 59570 47014
rect 121 46898 59570 47010
rect 121 46566 59743 46898
rect 430 46450 59570 46566
rect 121 46118 59743 46450
rect 121 46006 59570 46118
rect 430 46002 59570 46006
rect 430 45890 59743 46002
rect 121 45670 59743 45890
rect 121 45554 59570 45670
rect 121 45446 59743 45554
rect 430 45330 59743 45446
rect 121 45222 59743 45330
rect 121 45106 59570 45222
rect 121 44886 59743 45106
rect 430 44774 59743 44886
rect 430 44770 59570 44774
rect 121 44658 59570 44770
rect 121 44326 59743 44658
rect 430 44210 59570 44326
rect 121 43878 59743 44210
rect 121 43766 59570 43878
rect 430 43762 59570 43766
rect 430 43650 59743 43762
rect 121 43430 59743 43650
rect 121 43314 59570 43430
rect 121 43206 59743 43314
rect 430 43090 59743 43206
rect 121 42982 59743 43090
rect 121 42866 59570 42982
rect 121 42646 59743 42866
rect 430 42534 59743 42646
rect 430 42530 59570 42534
rect 121 42418 59570 42530
rect 121 42086 59743 42418
rect 430 41970 59570 42086
rect 121 41638 59743 41970
rect 121 41526 59570 41638
rect 430 41522 59570 41526
rect 430 41410 59743 41522
rect 121 41190 59743 41410
rect 121 41074 59570 41190
rect 121 40966 59743 41074
rect 430 40850 59743 40966
rect 121 40742 59743 40850
rect 121 40626 59570 40742
rect 121 40406 59743 40626
rect 430 40294 59743 40406
rect 430 40290 59570 40294
rect 121 40178 59570 40290
rect 121 39846 59743 40178
rect 430 39730 59570 39846
rect 121 39398 59743 39730
rect 121 39286 59570 39398
rect 430 39282 59570 39286
rect 430 39170 59743 39282
rect 121 38950 59743 39170
rect 121 38834 59570 38950
rect 121 38726 59743 38834
rect 430 38610 59743 38726
rect 121 38502 59743 38610
rect 121 38386 59570 38502
rect 121 38166 59743 38386
rect 430 38054 59743 38166
rect 430 38050 59570 38054
rect 121 37938 59570 38050
rect 121 37606 59743 37938
rect 430 37490 59570 37606
rect 121 37158 59743 37490
rect 121 37046 59570 37158
rect 430 37042 59570 37046
rect 430 36930 59743 37042
rect 121 36710 59743 36930
rect 121 36594 59570 36710
rect 121 36486 59743 36594
rect 430 36370 59743 36486
rect 121 36262 59743 36370
rect 121 36146 59570 36262
rect 121 35926 59743 36146
rect 430 35814 59743 35926
rect 430 35810 59570 35814
rect 121 35698 59570 35810
rect 121 35366 59743 35698
rect 430 35250 59570 35366
rect 121 34918 59743 35250
rect 121 34806 59570 34918
rect 430 34802 59570 34806
rect 430 34690 59743 34802
rect 121 34470 59743 34690
rect 121 34354 59570 34470
rect 121 34246 59743 34354
rect 430 34130 59743 34246
rect 121 34022 59743 34130
rect 121 33906 59570 34022
rect 121 33686 59743 33906
rect 430 33574 59743 33686
rect 430 33570 59570 33574
rect 121 33458 59570 33570
rect 121 33126 59743 33458
rect 430 33010 59570 33126
rect 121 32678 59743 33010
rect 121 32566 59570 32678
rect 430 32562 59570 32566
rect 430 32450 59743 32562
rect 121 32230 59743 32450
rect 121 32114 59570 32230
rect 121 32006 59743 32114
rect 430 31890 59743 32006
rect 121 31782 59743 31890
rect 121 31666 59570 31782
rect 121 31446 59743 31666
rect 430 31334 59743 31446
rect 430 31330 59570 31334
rect 121 31218 59570 31330
rect 121 30886 59743 31218
rect 430 30770 59570 30886
rect 121 30438 59743 30770
rect 121 30326 59570 30438
rect 430 30322 59570 30326
rect 430 30210 59743 30322
rect 121 29990 59743 30210
rect 121 29874 59570 29990
rect 121 29766 59743 29874
rect 430 29650 59743 29766
rect 121 29542 59743 29650
rect 121 29426 59570 29542
rect 121 29206 59743 29426
rect 430 29094 59743 29206
rect 430 29090 59570 29094
rect 121 28978 59570 29090
rect 121 28646 59743 28978
rect 430 28530 59570 28646
rect 121 28198 59743 28530
rect 121 28086 59570 28198
rect 430 28082 59570 28086
rect 430 27970 59743 28082
rect 121 27750 59743 27970
rect 121 27634 59570 27750
rect 121 27526 59743 27634
rect 430 27410 59743 27526
rect 121 27302 59743 27410
rect 121 27186 59570 27302
rect 121 26966 59743 27186
rect 430 26854 59743 26966
rect 430 26850 59570 26854
rect 121 26738 59570 26850
rect 121 26406 59743 26738
rect 430 26290 59570 26406
rect 121 25958 59743 26290
rect 121 25846 59570 25958
rect 430 25842 59570 25846
rect 430 25730 59743 25842
rect 121 25510 59743 25730
rect 121 25394 59570 25510
rect 121 25286 59743 25394
rect 430 25170 59743 25286
rect 121 25062 59743 25170
rect 121 24946 59570 25062
rect 121 24726 59743 24946
rect 430 24614 59743 24726
rect 430 24610 59570 24614
rect 121 24498 59570 24610
rect 121 24166 59743 24498
rect 430 24050 59570 24166
rect 121 23718 59743 24050
rect 121 23606 59570 23718
rect 430 23602 59570 23606
rect 430 23490 59743 23602
rect 121 23270 59743 23490
rect 121 23154 59570 23270
rect 121 23046 59743 23154
rect 430 22930 59743 23046
rect 121 22822 59743 22930
rect 121 22706 59570 22822
rect 121 22486 59743 22706
rect 430 22374 59743 22486
rect 430 22370 59570 22374
rect 121 22258 59570 22370
rect 121 21926 59743 22258
rect 430 21810 59570 21926
rect 121 21478 59743 21810
rect 121 21366 59570 21478
rect 430 21362 59570 21366
rect 430 21250 59743 21362
rect 121 21030 59743 21250
rect 121 20914 59570 21030
rect 121 20806 59743 20914
rect 430 20690 59743 20806
rect 121 20582 59743 20690
rect 121 20466 59570 20582
rect 121 20246 59743 20466
rect 430 20134 59743 20246
rect 430 20130 59570 20134
rect 121 20018 59570 20130
rect 121 19686 59743 20018
rect 430 19570 59570 19686
rect 121 19238 59743 19570
rect 121 19126 59570 19238
rect 430 19122 59570 19126
rect 430 19010 59743 19122
rect 121 18790 59743 19010
rect 121 18674 59570 18790
rect 121 18566 59743 18674
rect 430 18450 59743 18566
rect 121 18342 59743 18450
rect 121 18226 59570 18342
rect 121 18006 59743 18226
rect 430 17894 59743 18006
rect 430 17890 59570 17894
rect 121 17778 59570 17890
rect 121 17446 59743 17778
rect 430 17330 59570 17446
rect 121 16998 59743 17330
rect 121 16886 59570 16998
rect 430 16882 59570 16886
rect 430 16770 59743 16882
rect 121 16550 59743 16770
rect 121 16434 59570 16550
rect 121 16326 59743 16434
rect 430 16210 59743 16326
rect 121 16102 59743 16210
rect 121 15986 59570 16102
rect 121 15766 59743 15986
rect 430 15654 59743 15766
rect 430 15650 59570 15654
rect 121 15538 59570 15650
rect 121 15206 59743 15538
rect 430 15090 59570 15206
rect 121 14758 59743 15090
rect 121 14646 59570 14758
rect 430 14642 59570 14646
rect 430 14530 59743 14642
rect 121 14310 59743 14530
rect 121 14194 59570 14310
rect 121 14086 59743 14194
rect 430 13970 59743 14086
rect 121 13862 59743 13970
rect 121 13746 59570 13862
rect 121 13526 59743 13746
rect 430 13414 59743 13526
rect 430 13410 59570 13414
rect 121 13298 59570 13410
rect 121 12966 59743 13298
rect 430 12850 59570 12966
rect 121 12518 59743 12850
rect 121 12406 59570 12518
rect 430 12402 59570 12406
rect 430 12290 59743 12402
rect 121 12070 59743 12290
rect 121 11954 59570 12070
rect 121 11846 59743 11954
rect 430 11730 59743 11846
rect 121 11622 59743 11730
rect 121 11506 59570 11622
rect 121 11286 59743 11506
rect 430 11174 59743 11286
rect 430 11170 59570 11174
rect 121 11058 59570 11170
rect 121 10726 59743 11058
rect 430 10610 59570 10726
rect 121 10278 59743 10610
rect 121 10166 59570 10278
rect 430 10162 59570 10166
rect 430 10050 59743 10162
rect 121 9830 59743 10050
rect 121 9714 59570 9830
rect 121 9606 59743 9714
rect 430 9490 59743 9606
rect 121 9382 59743 9490
rect 121 9266 59570 9382
rect 121 9046 59743 9266
rect 430 8934 59743 9046
rect 430 8930 59570 8934
rect 121 8818 59570 8930
rect 121 8486 59743 8818
rect 430 8370 59570 8486
rect 121 8038 59743 8370
rect 121 7926 59570 8038
rect 430 7922 59570 7926
rect 430 7810 59743 7922
rect 121 7590 59743 7810
rect 121 7474 59570 7590
rect 121 7366 59743 7474
rect 430 7250 59743 7366
rect 121 7142 59743 7250
rect 121 7026 59570 7142
rect 121 6806 59743 7026
rect 430 6694 59743 6806
rect 430 6690 59570 6694
rect 121 6578 59570 6690
rect 121 6246 59743 6578
rect 430 6130 59570 6246
rect 121 5798 59743 6130
rect 121 5686 59570 5798
rect 430 5682 59570 5686
rect 430 5570 59743 5682
rect 121 5350 59743 5570
rect 121 5234 59570 5350
rect 121 5126 59743 5234
rect 430 5010 59743 5126
rect 121 4902 59743 5010
rect 121 4786 59570 4902
rect 121 4566 59743 4786
rect 430 4454 59743 4566
rect 430 4450 59570 4454
rect 121 4338 59570 4450
rect 121 4006 59743 4338
rect 430 3890 59570 4006
rect 121 1358 59743 3890
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
<< obsm4 >>
rect 1022 1508 2194 57783
rect 2414 1508 9874 57783
rect 10094 1508 17554 57783
rect 17774 1508 25234 57783
rect 25454 1508 32914 57783
rect 33134 1508 40594 57783
rect 40814 1508 48274 57783
rect 48494 1508 55954 57783
rect 56174 1508 58954 57783
rect 1022 1409 58954 1508
<< labels >>
rlabel metal2 s 47264 59600 47320 60000 6 blinker_do[0]
port 1 nsew signal input
rlabel metal2 s 47824 59600 47880 60000 6 blinker_do[1]
port 2 nsew signal input
rlabel metal2 s 48384 59600 48440 60000 6 blinker_do[2]
port 3 nsew signal input
rlabel metal3 s 59600 20048 60000 20104 6 custom_settings[0]
port 4 nsew signal output
rlabel metal3 s 59600 24528 60000 24584 6 custom_settings[10]
port 5 nsew signal output
rlabel metal3 s 59600 24976 60000 25032 6 custom_settings[11]
port 6 nsew signal output
rlabel metal3 s 59600 25424 60000 25480 6 custom_settings[12]
port 7 nsew signal output
rlabel metal3 s 59600 25872 60000 25928 6 custom_settings[13]
port 8 nsew signal output
rlabel metal3 s 59600 26320 60000 26376 6 custom_settings[14]
port 9 nsew signal output
rlabel metal3 s 59600 26768 60000 26824 6 custom_settings[15]
port 10 nsew signal output
rlabel metal3 s 59600 27216 60000 27272 6 custom_settings[16]
port 11 nsew signal output
rlabel metal3 s 59600 27664 60000 27720 6 custom_settings[17]
port 12 nsew signal output
rlabel metal3 s 59600 28112 60000 28168 6 custom_settings[18]
port 13 nsew signal output
rlabel metal3 s 59600 28560 60000 28616 6 custom_settings[19]
port 14 nsew signal output
rlabel metal3 s 59600 20496 60000 20552 6 custom_settings[1]
port 15 nsew signal output
rlabel metal3 s 59600 29008 60000 29064 6 custom_settings[20]
port 16 nsew signal output
rlabel metal3 s 59600 29456 60000 29512 6 custom_settings[21]
port 17 nsew signal output
rlabel metal3 s 59600 29904 60000 29960 6 custom_settings[22]
port 18 nsew signal output
rlabel metal3 s 59600 30352 60000 30408 6 custom_settings[23]
port 19 nsew signal output
rlabel metal3 s 59600 30800 60000 30856 6 custom_settings[24]
port 20 nsew signal output
rlabel metal3 s 59600 31248 60000 31304 6 custom_settings[25]
port 21 nsew signal output
rlabel metal3 s 59600 31696 60000 31752 6 custom_settings[26]
port 22 nsew signal output
rlabel metal3 s 59600 32144 60000 32200 6 custom_settings[27]
port 23 nsew signal output
rlabel metal3 s 59600 32592 60000 32648 6 custom_settings[28]
port 24 nsew signal output
rlabel metal3 s 59600 33040 60000 33096 6 custom_settings[29]
port 25 nsew signal output
rlabel metal3 s 59600 20944 60000 21000 6 custom_settings[2]
port 26 nsew signal output
rlabel metal3 s 59600 33488 60000 33544 6 custom_settings[30]
port 27 nsew signal output
rlabel metal3 s 59600 33936 60000 33992 6 custom_settings[31]
port 28 nsew signal output
rlabel metal3 s 59600 21392 60000 21448 6 custom_settings[3]
port 29 nsew signal output
rlabel metal3 s 59600 21840 60000 21896 6 custom_settings[4]
port 30 nsew signal output
rlabel metal3 s 59600 22288 60000 22344 6 custom_settings[5]
port 31 nsew signal output
rlabel metal3 s 59600 22736 60000 22792 6 custom_settings[6]
port 32 nsew signal output
rlabel metal3 s 59600 23184 60000 23240 6 custom_settings[7]
port 33 nsew signal output
rlabel metal3 s 59600 23632 60000 23688 6 custom_settings[8]
port 34 nsew signal output
rlabel metal3 s 59600 24080 60000 24136 6 custom_settings[9]
port 35 nsew signal output
rlabel metal2 s 2464 59600 2520 60000 6 io_in[0]
port 36 nsew signal input
rlabel metal2 s 8064 59600 8120 60000 6 io_in[10]
port 37 nsew signal input
rlabel metal2 s 8624 59600 8680 60000 6 io_in[11]
port 38 nsew signal input
rlabel metal2 s 9184 59600 9240 60000 6 io_in[12]
port 39 nsew signal input
rlabel metal2 s 9744 59600 9800 60000 6 io_in[13]
port 40 nsew signal input
rlabel metal2 s 10304 59600 10360 60000 6 io_in[14]
port 41 nsew signal input
rlabel metal2 s 10864 59600 10920 60000 6 io_in[15]
port 42 nsew signal input
rlabel metal2 s 11424 59600 11480 60000 6 io_in[16]
port 43 nsew signal input
rlabel metal2 s 11984 59600 12040 60000 6 io_in[17]
port 44 nsew signal input
rlabel metal2 s 12544 59600 12600 60000 6 io_in[18]
port 45 nsew signal input
rlabel metal2 s 13104 59600 13160 60000 6 io_in[19]
port 46 nsew signal input
rlabel metal2 s 3024 59600 3080 60000 6 io_in[1]
port 47 nsew signal input
rlabel metal2 s 13664 59600 13720 60000 6 io_in[20]
port 48 nsew signal input
rlabel metal2 s 14224 59600 14280 60000 6 io_in[21]
port 49 nsew signal input
rlabel metal2 s 14784 59600 14840 60000 6 io_in[22]
port 50 nsew signal input
rlabel metal2 s 15344 59600 15400 60000 6 io_in[23]
port 51 nsew signal input
rlabel metal2 s 15904 59600 15960 60000 6 io_in[24]
port 52 nsew signal input
rlabel metal2 s 16464 59600 16520 60000 6 io_in[25]
port 53 nsew signal input
rlabel metal2 s 17024 59600 17080 60000 6 io_in[26]
port 54 nsew signal input
rlabel metal2 s 17584 59600 17640 60000 6 io_in[27]
port 55 nsew signal input
rlabel metal2 s 18144 59600 18200 60000 6 io_in[28]
port 56 nsew signal input
rlabel metal2 s 18704 59600 18760 60000 6 io_in[29]
port 57 nsew signal input
rlabel metal2 s 3584 59600 3640 60000 6 io_in[2]
port 58 nsew signal input
rlabel metal2 s 19264 59600 19320 60000 6 io_in[30]
port 59 nsew signal input
rlabel metal2 s 19824 59600 19880 60000 6 io_in[31]
port 60 nsew signal input
rlabel metal2 s 20384 59600 20440 60000 6 io_in[32]
port 61 nsew signal input
rlabel metal2 s 20944 59600 21000 60000 6 io_in[33]
port 62 nsew signal input
rlabel metal2 s 21504 59600 21560 60000 6 io_in[34]
port 63 nsew signal input
rlabel metal2 s 22064 59600 22120 60000 6 io_in[35]
port 64 nsew signal input
rlabel metal2 s 22624 59600 22680 60000 6 io_in[36]
port 65 nsew signal input
rlabel metal2 s 23184 59600 23240 60000 6 io_in[37]
port 66 nsew signal input
rlabel metal2 s 4144 59600 4200 60000 6 io_in[3]
port 67 nsew signal input
rlabel metal2 s 4704 59600 4760 60000 6 io_in[4]
port 68 nsew signal input
rlabel metal2 s 5264 59600 5320 60000 6 io_in[5]
port 69 nsew signal input
rlabel metal2 s 5824 59600 5880 60000 6 io_in[6]
port 70 nsew signal input
rlabel metal2 s 6384 59600 6440 60000 6 io_in[7]
port 71 nsew signal input
rlabel metal2 s 6944 59600 7000 60000 6 io_in[8]
port 72 nsew signal input
rlabel metal2 s 7504 59600 7560 60000 6 io_in[9]
port 73 nsew signal input
rlabel metal3 s 0 3920 400 3976 6 io_oeb[0]
port 74 nsew signal output
rlabel metal3 s 0 9520 400 9576 6 io_oeb[10]
port 75 nsew signal output
rlabel metal3 s 0 10080 400 10136 6 io_oeb[11]
port 76 nsew signal output
rlabel metal3 s 0 10640 400 10696 6 io_oeb[12]
port 77 nsew signal output
rlabel metal3 s 0 11200 400 11256 6 io_oeb[13]
port 78 nsew signal output
rlabel metal3 s 0 11760 400 11816 6 io_oeb[14]
port 79 nsew signal output
rlabel metal3 s 0 12320 400 12376 6 io_oeb[15]
port 80 nsew signal output
rlabel metal3 s 0 12880 400 12936 6 io_oeb[16]
port 81 nsew signal output
rlabel metal3 s 0 13440 400 13496 6 io_oeb[17]
port 82 nsew signal output
rlabel metal3 s 0 14000 400 14056 6 io_oeb[18]
port 83 nsew signal output
rlabel metal3 s 0 14560 400 14616 6 io_oeb[19]
port 84 nsew signal output
rlabel metal3 s 0 4480 400 4536 6 io_oeb[1]
port 85 nsew signal output
rlabel metal3 s 0 15120 400 15176 6 io_oeb[20]
port 86 nsew signal output
rlabel metal3 s 0 15680 400 15736 6 io_oeb[21]
port 87 nsew signal output
rlabel metal3 s 0 16240 400 16296 6 io_oeb[22]
port 88 nsew signal output
rlabel metal3 s 0 16800 400 16856 6 io_oeb[23]
port 89 nsew signal output
rlabel metal3 s 0 17360 400 17416 6 io_oeb[24]
port 90 nsew signal output
rlabel metal3 s 0 17920 400 17976 6 io_oeb[25]
port 91 nsew signal output
rlabel metal3 s 0 18480 400 18536 6 io_oeb[26]
port 92 nsew signal output
rlabel metal3 s 0 19040 400 19096 6 io_oeb[27]
port 93 nsew signal output
rlabel metal3 s 0 19600 400 19656 6 io_oeb[28]
port 94 nsew signal output
rlabel metal3 s 0 20160 400 20216 6 io_oeb[29]
port 95 nsew signal output
rlabel metal3 s 0 5040 400 5096 6 io_oeb[2]
port 96 nsew signal output
rlabel metal3 s 0 20720 400 20776 6 io_oeb[30]
port 97 nsew signal output
rlabel metal3 s 0 21280 400 21336 6 io_oeb[31]
port 98 nsew signal output
rlabel metal3 s 0 21840 400 21896 6 io_oeb[32]
port 99 nsew signal output
rlabel metal3 s 0 22400 400 22456 6 io_oeb[33]
port 100 nsew signal output
rlabel metal3 s 0 22960 400 23016 6 io_oeb[34]
port 101 nsew signal output
rlabel metal3 s 0 23520 400 23576 6 io_oeb[35]
port 102 nsew signal output
rlabel metal3 s 0 24080 400 24136 6 io_oeb[36]
port 103 nsew signal output
rlabel metal3 s 0 24640 400 24696 6 io_oeb[37]
port 104 nsew signal output
rlabel metal3 s 0 5600 400 5656 6 io_oeb[3]
port 105 nsew signal output
rlabel metal3 s 0 6160 400 6216 6 io_oeb[4]
port 106 nsew signal output
rlabel metal3 s 0 6720 400 6776 6 io_oeb[5]
port 107 nsew signal output
rlabel metal3 s 0 7280 400 7336 6 io_oeb[6]
port 108 nsew signal output
rlabel metal3 s 0 7840 400 7896 6 io_oeb[7]
port 109 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 io_oeb[8]
port 110 nsew signal output
rlabel metal3 s 0 8960 400 9016 6 io_oeb[9]
port 111 nsew signal output
rlabel metal2 s 23744 59600 23800 60000 6 io_out[0]
port 112 nsew signal output
rlabel metal2 s 29344 59600 29400 60000 6 io_out[10]
port 113 nsew signal output
rlabel metal2 s 29904 59600 29960 60000 6 io_out[11]
port 114 nsew signal output
rlabel metal2 s 30464 59600 30520 60000 6 io_out[12]
port 115 nsew signal output
rlabel metal2 s 31024 59600 31080 60000 6 io_out[13]
port 116 nsew signal output
rlabel metal2 s 31584 59600 31640 60000 6 io_out[14]
port 117 nsew signal output
rlabel metal2 s 32144 59600 32200 60000 6 io_out[15]
port 118 nsew signal output
rlabel metal2 s 32704 59600 32760 60000 6 io_out[16]
port 119 nsew signal output
rlabel metal2 s 33264 59600 33320 60000 6 io_out[17]
port 120 nsew signal output
rlabel metal2 s 33824 59600 33880 60000 6 io_out[18]
port 121 nsew signal output
rlabel metal2 s 34384 59600 34440 60000 6 io_out[19]
port 122 nsew signal output
rlabel metal2 s 24304 59600 24360 60000 6 io_out[1]
port 123 nsew signal output
rlabel metal2 s 34944 59600 35000 60000 6 io_out[20]
port 124 nsew signal output
rlabel metal2 s 35504 59600 35560 60000 6 io_out[21]
port 125 nsew signal output
rlabel metal2 s 36064 59600 36120 60000 6 io_out[22]
port 126 nsew signal output
rlabel metal2 s 36624 59600 36680 60000 6 io_out[23]
port 127 nsew signal output
rlabel metal2 s 37184 59600 37240 60000 6 io_out[24]
port 128 nsew signal output
rlabel metal2 s 37744 59600 37800 60000 6 io_out[25]
port 129 nsew signal output
rlabel metal2 s 38304 59600 38360 60000 6 io_out[26]
port 130 nsew signal output
rlabel metal2 s 38864 59600 38920 60000 6 io_out[27]
port 131 nsew signal output
rlabel metal2 s 39424 59600 39480 60000 6 io_out[28]
port 132 nsew signal output
rlabel metal2 s 39984 59600 40040 60000 6 io_out[29]
port 133 nsew signal output
rlabel metal2 s 24864 59600 24920 60000 6 io_out[2]
port 134 nsew signal output
rlabel metal2 s 40544 59600 40600 60000 6 io_out[30]
port 135 nsew signal output
rlabel metal2 s 41104 59600 41160 60000 6 io_out[31]
port 136 nsew signal output
rlabel metal2 s 41664 59600 41720 60000 6 io_out[32]
port 137 nsew signal output
rlabel metal2 s 42224 59600 42280 60000 6 io_out[33]
port 138 nsew signal output
rlabel metal2 s 42784 59600 42840 60000 6 io_out[34]
port 139 nsew signal output
rlabel metal2 s 43344 59600 43400 60000 6 io_out[35]
port 140 nsew signal output
rlabel metal2 s 43904 59600 43960 60000 6 io_out[36]
port 141 nsew signal output
rlabel metal2 s 44464 59600 44520 60000 6 io_out[37]
port 142 nsew signal output
rlabel metal2 s 25424 59600 25480 60000 6 io_out[3]
port 143 nsew signal output
rlabel metal2 s 25984 59600 26040 60000 6 io_out[4]
port 144 nsew signal output
rlabel metal2 s 26544 59600 26600 60000 6 io_out[5]
port 145 nsew signal output
rlabel metal2 s 27104 59600 27160 60000 6 io_out[6]
port 146 nsew signal output
rlabel metal2 s 27664 59600 27720 60000 6 io_out[7]
port 147 nsew signal output
rlabel metal2 s 28224 59600 28280 60000 6 io_out[8]
port 148 nsew signal output
rlabel metal2 s 28784 59600 28840 60000 6 io_out[9]
port 149 nsew signal output
rlabel metal2 s 45024 59600 45080 60000 6 irq[0]
port 150 nsew signal output
rlabel metal2 s 45584 59600 45640 60000 6 irq[1]
port 151 nsew signal output
rlabel metal2 s 46144 59600 46200 60000 6 irq[2]
port 152 nsew signal output
rlabel metal3 s 0 39200 400 39256 6 mc14500_do[0]
port 153 nsew signal input
rlabel metal3 s 0 44800 400 44856 6 mc14500_do[10]
port 154 nsew signal input
rlabel metal3 s 0 45360 400 45416 6 mc14500_do[11]
port 155 nsew signal input
rlabel metal3 s 0 45920 400 45976 6 mc14500_do[12]
port 156 nsew signal input
rlabel metal3 s 0 46480 400 46536 6 mc14500_do[13]
port 157 nsew signal input
rlabel metal3 s 0 47040 400 47096 6 mc14500_do[14]
port 158 nsew signal input
rlabel metal3 s 0 47600 400 47656 6 mc14500_do[15]
port 159 nsew signal input
rlabel metal3 s 0 48160 400 48216 6 mc14500_do[16]
port 160 nsew signal input
rlabel metal3 s 0 48720 400 48776 6 mc14500_do[17]
port 161 nsew signal input
rlabel metal3 s 0 49280 400 49336 6 mc14500_do[18]
port 162 nsew signal input
rlabel metal3 s 0 49840 400 49896 6 mc14500_do[19]
port 163 nsew signal input
rlabel metal3 s 0 39760 400 39816 6 mc14500_do[1]
port 164 nsew signal input
rlabel metal3 s 0 50400 400 50456 6 mc14500_do[20]
port 165 nsew signal input
rlabel metal3 s 0 50960 400 51016 6 mc14500_do[21]
port 166 nsew signal input
rlabel metal3 s 0 51520 400 51576 6 mc14500_do[22]
port 167 nsew signal input
rlabel metal3 s 0 52080 400 52136 6 mc14500_do[23]
port 168 nsew signal input
rlabel metal3 s 0 52640 400 52696 6 mc14500_do[24]
port 169 nsew signal input
rlabel metal3 s 0 53200 400 53256 6 mc14500_do[25]
port 170 nsew signal input
rlabel metal3 s 0 53760 400 53816 6 mc14500_do[26]
port 171 nsew signal input
rlabel metal3 s 0 54320 400 54376 6 mc14500_do[27]
port 172 nsew signal input
rlabel metal3 s 0 54880 400 54936 6 mc14500_do[28]
port 173 nsew signal input
rlabel metal3 s 0 55440 400 55496 6 mc14500_do[29]
port 174 nsew signal input
rlabel metal3 s 0 40320 400 40376 6 mc14500_do[2]
port 175 nsew signal input
rlabel metal3 s 0 56000 400 56056 6 mc14500_do[30]
port 176 nsew signal input
rlabel metal3 s 0 40880 400 40936 6 mc14500_do[3]
port 177 nsew signal input
rlabel metal3 s 0 41440 400 41496 6 mc14500_do[4]
port 178 nsew signal input
rlabel metal3 s 0 42000 400 42056 6 mc14500_do[5]
port 179 nsew signal input
rlabel metal3 s 0 42560 400 42616 6 mc14500_do[6]
port 180 nsew signal input
rlabel metal3 s 0 43120 400 43176 6 mc14500_do[7]
port 181 nsew signal input
rlabel metal3 s 0 43680 400 43736 6 mc14500_do[8]
port 182 nsew signal input
rlabel metal3 s 0 44240 400 44296 6 mc14500_do[9]
port 183 nsew signal input
rlabel metal2 s 49504 59600 49560 60000 6 mc14500_sram_addr[0]
port 184 nsew signal input
rlabel metal2 s 50064 59600 50120 60000 6 mc14500_sram_addr[1]
port 185 nsew signal input
rlabel metal2 s 50624 59600 50680 60000 6 mc14500_sram_addr[2]
port 186 nsew signal input
rlabel metal2 s 51184 59600 51240 60000 6 mc14500_sram_addr[3]
port 187 nsew signal input
rlabel metal2 s 51744 59600 51800 60000 6 mc14500_sram_addr[4]
port 188 nsew signal input
rlabel metal2 s 52304 59600 52360 60000 6 mc14500_sram_addr[5]
port 189 nsew signal input
rlabel metal2 s 57344 59600 57400 60000 6 mc14500_sram_gwe
port 190 nsew signal input
rlabel metal2 s 52864 59600 52920 60000 6 mc14500_sram_in[0]
port 191 nsew signal input
rlabel metal2 s 53424 59600 53480 60000 6 mc14500_sram_in[1]
port 192 nsew signal input
rlabel metal2 s 53984 59600 54040 60000 6 mc14500_sram_in[2]
port 193 nsew signal input
rlabel metal2 s 54544 59600 54600 60000 6 mc14500_sram_in[3]
port 194 nsew signal input
rlabel metal2 s 55104 59600 55160 60000 6 mc14500_sram_in[4]
port 195 nsew signal input
rlabel metal2 s 55664 59600 55720 60000 6 mc14500_sram_in[5]
port 196 nsew signal input
rlabel metal2 s 56224 59600 56280 60000 6 mc14500_sram_in[6]
port 197 nsew signal input
rlabel metal2 s 56784 59600 56840 60000 6 mc14500_sram_in[7]
port 198 nsew signal input
rlabel metal2 s 42224 0 42280 400 6 qcpu_do[0]
port 199 nsew signal input
rlabel metal2 s 46704 0 46760 400 6 qcpu_do[10]
port 200 nsew signal input
rlabel metal2 s 47152 0 47208 400 6 qcpu_do[11]
port 201 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 qcpu_do[12]
port 202 nsew signal input
rlabel metal2 s 48048 0 48104 400 6 qcpu_do[13]
port 203 nsew signal input
rlabel metal2 s 48496 0 48552 400 6 qcpu_do[14]
port 204 nsew signal input
rlabel metal2 s 48944 0 49000 400 6 qcpu_do[15]
port 205 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 qcpu_do[16]
port 206 nsew signal input
rlabel metal2 s 49840 0 49896 400 6 qcpu_do[17]
port 207 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 qcpu_do[18]
port 208 nsew signal input
rlabel metal2 s 50736 0 50792 400 6 qcpu_do[19]
port 209 nsew signal input
rlabel metal2 s 42672 0 42728 400 6 qcpu_do[1]
port 210 nsew signal input
rlabel metal2 s 51184 0 51240 400 6 qcpu_do[20]
port 211 nsew signal input
rlabel metal2 s 51632 0 51688 400 6 qcpu_do[21]
port 212 nsew signal input
rlabel metal2 s 52080 0 52136 400 6 qcpu_do[22]
port 213 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 qcpu_do[23]
port 214 nsew signal input
rlabel metal2 s 52976 0 53032 400 6 qcpu_do[24]
port 215 nsew signal input
rlabel metal2 s 53424 0 53480 400 6 qcpu_do[25]
port 216 nsew signal input
rlabel metal2 s 53872 0 53928 400 6 qcpu_do[26]
port 217 nsew signal input
rlabel metal2 s 54320 0 54376 400 6 qcpu_do[27]
port 218 nsew signal input
rlabel metal2 s 54768 0 54824 400 6 qcpu_do[28]
port 219 nsew signal input
rlabel metal2 s 55216 0 55272 400 6 qcpu_do[29]
port 220 nsew signal input
rlabel metal2 s 43120 0 43176 400 6 qcpu_do[2]
port 221 nsew signal input
rlabel metal2 s 55664 0 55720 400 6 qcpu_do[30]
port 222 nsew signal input
rlabel metal2 s 56112 0 56168 400 6 qcpu_do[31]
port 223 nsew signal input
rlabel metal2 s 56560 0 56616 400 6 qcpu_do[32]
port 224 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 qcpu_do[3]
port 225 nsew signal input
rlabel metal2 s 44016 0 44072 400 6 qcpu_do[4]
port 226 nsew signal input
rlabel metal2 s 44464 0 44520 400 6 qcpu_do[5]
port 227 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 qcpu_do[6]
port 228 nsew signal input
rlabel metal2 s 45360 0 45416 400 6 qcpu_do[7]
port 229 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 qcpu_do[8]
port 230 nsew signal input
rlabel metal2 s 46256 0 46312 400 6 qcpu_do[9]
port 231 nsew signal input
rlabel metal3 s 59600 34384 60000 34440 6 qcpu_oeb[0]
port 232 nsew signal input
rlabel metal3 s 59600 38864 60000 38920 6 qcpu_oeb[10]
port 233 nsew signal input
rlabel metal3 s 59600 39312 60000 39368 6 qcpu_oeb[11]
port 234 nsew signal input
rlabel metal3 s 59600 39760 60000 39816 6 qcpu_oeb[12]
port 235 nsew signal input
rlabel metal3 s 59600 40208 60000 40264 6 qcpu_oeb[13]
port 236 nsew signal input
rlabel metal3 s 59600 40656 60000 40712 6 qcpu_oeb[14]
port 237 nsew signal input
rlabel metal3 s 59600 41104 60000 41160 6 qcpu_oeb[15]
port 238 nsew signal input
rlabel metal3 s 59600 41552 60000 41608 6 qcpu_oeb[16]
port 239 nsew signal input
rlabel metal3 s 59600 42000 60000 42056 6 qcpu_oeb[17]
port 240 nsew signal input
rlabel metal3 s 59600 42448 60000 42504 6 qcpu_oeb[18]
port 241 nsew signal input
rlabel metal3 s 59600 42896 60000 42952 6 qcpu_oeb[19]
port 242 nsew signal input
rlabel metal3 s 59600 34832 60000 34888 6 qcpu_oeb[1]
port 243 nsew signal input
rlabel metal3 s 59600 43344 60000 43400 6 qcpu_oeb[20]
port 244 nsew signal input
rlabel metal3 s 59600 43792 60000 43848 6 qcpu_oeb[21]
port 245 nsew signal input
rlabel metal3 s 59600 44240 60000 44296 6 qcpu_oeb[22]
port 246 nsew signal input
rlabel metal3 s 59600 44688 60000 44744 6 qcpu_oeb[23]
port 247 nsew signal input
rlabel metal3 s 59600 45136 60000 45192 6 qcpu_oeb[24]
port 248 nsew signal input
rlabel metal3 s 59600 45584 60000 45640 6 qcpu_oeb[25]
port 249 nsew signal input
rlabel metal3 s 59600 46032 60000 46088 6 qcpu_oeb[26]
port 250 nsew signal input
rlabel metal3 s 59600 46480 60000 46536 6 qcpu_oeb[27]
port 251 nsew signal input
rlabel metal3 s 59600 46928 60000 46984 6 qcpu_oeb[28]
port 252 nsew signal input
rlabel metal3 s 59600 47376 60000 47432 6 qcpu_oeb[29]
port 253 nsew signal input
rlabel metal3 s 59600 35280 60000 35336 6 qcpu_oeb[2]
port 254 nsew signal input
rlabel metal3 s 59600 47824 60000 47880 6 qcpu_oeb[30]
port 255 nsew signal input
rlabel metal3 s 59600 48272 60000 48328 6 qcpu_oeb[31]
port 256 nsew signal input
rlabel metal3 s 59600 48720 60000 48776 6 qcpu_oeb[32]
port 257 nsew signal input
rlabel metal3 s 59600 35728 60000 35784 6 qcpu_oeb[3]
port 258 nsew signal input
rlabel metal3 s 59600 36176 60000 36232 6 qcpu_oeb[4]
port 259 nsew signal input
rlabel metal3 s 59600 36624 60000 36680 6 qcpu_oeb[5]
port 260 nsew signal input
rlabel metal3 s 59600 37072 60000 37128 6 qcpu_oeb[6]
port 261 nsew signal input
rlabel metal3 s 59600 37520 60000 37576 6 qcpu_oeb[7]
port 262 nsew signal input
rlabel metal3 s 59600 37968 60000 38024 6 qcpu_oeb[8]
port 263 nsew signal input
rlabel metal3 s 59600 38416 60000 38472 6 qcpu_oeb[9]
port 264 nsew signal input
rlabel metal2 s 57008 0 57064 400 6 qcpu_sram_addr[0]
port 265 nsew signal input
rlabel metal2 s 57456 0 57512 400 6 qcpu_sram_addr[1]
port 266 nsew signal input
rlabel metal2 s 57904 0 57960 400 6 qcpu_sram_addr[2]
port 267 nsew signal input
rlabel metal2 s 58352 0 58408 400 6 qcpu_sram_addr[3]
port 268 nsew signal input
rlabel metal2 s 58800 0 58856 400 6 qcpu_sram_addr[4]
port 269 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 qcpu_sram_addr[5]
port 270 nsew signal input
rlabel metal2 s 59696 0 59752 400 6 qcpu_sram_gwe
port 271 nsew signal input
rlabel metal3 s 59600 49168 60000 49224 6 qcpu_sram_in[0]
port 272 nsew signal input
rlabel metal3 s 59600 49616 60000 49672 6 qcpu_sram_in[1]
port 273 nsew signal input
rlabel metal3 s 59600 50064 60000 50120 6 qcpu_sram_in[2]
port 274 nsew signal input
rlabel metal3 s 59600 50512 60000 50568 6 qcpu_sram_in[3]
port 275 nsew signal input
rlabel metal3 s 59600 50960 60000 51016 6 qcpu_sram_in[4]
port 276 nsew signal input
rlabel metal3 s 59600 51408 60000 51464 6 qcpu_sram_in[5]
port 277 nsew signal input
rlabel metal3 s 59600 51856 60000 51912 6 qcpu_sram_in[6]
port 278 nsew signal input
rlabel metal3 s 59600 52304 60000 52360 6 qcpu_sram_in[7]
port 279 nsew signal input
rlabel metal3 s 59600 52752 60000 52808 6 qcpu_sram_out[0]
port 280 nsew signal output
rlabel metal3 s 59600 53200 60000 53256 6 qcpu_sram_out[1]
port 281 nsew signal output
rlabel metal3 s 59600 53648 60000 53704 6 qcpu_sram_out[2]
port 282 nsew signal output
rlabel metal3 s 59600 54096 60000 54152 6 qcpu_sram_out[3]
port 283 nsew signal output
rlabel metal3 s 59600 54544 60000 54600 6 qcpu_sram_out[4]
port 284 nsew signal output
rlabel metal3 s 59600 54992 60000 55048 6 qcpu_sram_out[5]
port 285 nsew signal output
rlabel metal3 s 59600 55440 60000 55496 6 qcpu_sram_out[6]
port 286 nsew signal output
rlabel metal3 s 59600 55888 60000 55944 6 qcpu_sram_out[7]
port 287 nsew signal output
rlabel metal2 s 46704 59600 46760 60000 6 rst_blinker
port 288 nsew signal output
rlabel metal3 s 0 38640 400 38696 6 rst_mc14500
port 289 nsew signal output
rlabel metal3 s 0 38080 400 38136 6 rst_qcpu
port 290 nsew signal output
rlabel metal3 s 0 25200 400 25256 6 rst_sid
port 291 nsew signal output
rlabel metal2 s 48944 59600 49000 60000 6 rst_sn76489
port 292 nsew signal output
rlabel metal3 s 0 25760 400 25816 6 sid_do[0]
port 293 nsew signal input
rlabel metal3 s 0 31360 400 31416 6 sid_do[10]
port 294 nsew signal input
rlabel metal3 s 0 31920 400 31976 6 sid_do[11]
port 295 nsew signal input
rlabel metal3 s 0 32480 400 32536 6 sid_do[12]
port 296 nsew signal input
rlabel metal3 s 0 33040 400 33096 6 sid_do[13]
port 297 nsew signal input
rlabel metal3 s 0 33600 400 33656 6 sid_do[14]
port 298 nsew signal input
rlabel metal3 s 0 34160 400 34216 6 sid_do[15]
port 299 nsew signal input
rlabel metal3 s 0 34720 400 34776 6 sid_do[16]
port 300 nsew signal input
rlabel metal3 s 0 35280 400 35336 6 sid_do[17]
port 301 nsew signal input
rlabel metal3 s 0 35840 400 35896 6 sid_do[18]
port 302 nsew signal input
rlabel metal3 s 0 36400 400 36456 6 sid_do[19]
port 303 nsew signal input
rlabel metal3 s 0 26320 400 26376 6 sid_do[1]
port 304 nsew signal input
rlabel metal3 s 0 36960 400 37016 6 sid_do[20]
port 305 nsew signal input
rlabel metal3 s 0 26880 400 26936 6 sid_do[2]
port 306 nsew signal input
rlabel metal3 s 0 27440 400 27496 6 sid_do[3]
port 307 nsew signal input
rlabel metal3 s 0 28000 400 28056 6 sid_do[4]
port 308 nsew signal input
rlabel metal3 s 0 28560 400 28616 6 sid_do[5]
port 309 nsew signal input
rlabel metal3 s 0 29120 400 29176 6 sid_do[6]
port 310 nsew signal input
rlabel metal3 s 0 29680 400 29736 6 sid_do[7]
port 311 nsew signal input
rlabel metal3 s 0 30240 400 30296 6 sid_do[8]
port 312 nsew signal input
rlabel metal3 s 0 30800 400 30856 6 sid_do[9]
port 313 nsew signal input
rlabel metal3 s 0 37520 400 37576 6 sid_oeb
port 314 nsew signal input
rlabel metal2 s 29680 0 29736 400 6 sn76489_do[0]
port 315 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 sn76489_do[10]
port 316 nsew signal input
rlabel metal2 s 34608 0 34664 400 6 sn76489_do[11]
port 317 nsew signal input
rlabel metal2 s 35056 0 35112 400 6 sn76489_do[12]
port 318 nsew signal input
rlabel metal2 s 35504 0 35560 400 6 sn76489_do[13]
port 319 nsew signal input
rlabel metal2 s 35952 0 36008 400 6 sn76489_do[14]
port 320 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 sn76489_do[15]
port 321 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 sn76489_do[16]
port 322 nsew signal input
rlabel metal2 s 37296 0 37352 400 6 sn76489_do[17]
port 323 nsew signal input
rlabel metal2 s 37744 0 37800 400 6 sn76489_do[18]
port 324 nsew signal input
rlabel metal2 s 38192 0 38248 400 6 sn76489_do[19]
port 325 nsew signal input
rlabel metal2 s 30128 0 30184 400 6 sn76489_do[1]
port 326 nsew signal input
rlabel metal2 s 38640 0 38696 400 6 sn76489_do[20]
port 327 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 sn76489_do[21]
port 328 nsew signal input
rlabel metal2 s 39536 0 39592 400 6 sn76489_do[22]
port 329 nsew signal input
rlabel metal2 s 39984 0 40040 400 6 sn76489_do[23]
port 330 nsew signal input
rlabel metal2 s 40432 0 40488 400 6 sn76489_do[24]
port 331 nsew signal input
rlabel metal2 s 40880 0 40936 400 6 sn76489_do[25]
port 332 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 sn76489_do[26]
port 333 nsew signal input
rlabel metal2 s 41776 0 41832 400 6 sn76489_do[27]
port 334 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 sn76489_do[2]
port 335 nsew signal input
rlabel metal2 s 31024 0 31080 400 6 sn76489_do[3]
port 336 nsew signal input
rlabel metal2 s 31472 0 31528 400 6 sn76489_do[4]
port 337 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 sn76489_do[5]
port 338 nsew signal input
rlabel metal2 s 32368 0 32424 400 6 sn76489_do[6]
port 339 nsew signal input
rlabel metal2 s 32816 0 32872 400 6 sn76489_do[7]
port 340 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 sn76489_do[8]
port 341 nsew signal input
rlabel metal2 s 33712 0 33768 400 6 sn76489_do[9]
port 342 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 343 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 343 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 343 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 343 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 344 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 344 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 344 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 344 nsew ground bidirectional
rlabel metal2 s 112 0 168 400 6 wb_clk_i
port 345 nsew signal input
rlabel metal2 s 560 0 616 400 6 wb_rst_i
port 346 nsew signal input
rlabel metal3 s 59600 19600 60000 19656 6 wbs_ack_o
port 347 nsew signal output
rlabel metal2 s 1008 0 1064 400 6 wbs_adr_i[0]
port 348 nsew signal input
rlabel metal2 s 5488 0 5544 400 6 wbs_adr_i[10]
port 349 nsew signal input
rlabel metal2 s 5936 0 5992 400 6 wbs_adr_i[11]
port 350 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 wbs_adr_i[12]
port 351 nsew signal input
rlabel metal2 s 6832 0 6888 400 6 wbs_adr_i[13]
port 352 nsew signal input
rlabel metal2 s 7280 0 7336 400 6 wbs_adr_i[14]
port 353 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 wbs_adr_i[15]
port 354 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wbs_adr_i[16]
port 355 nsew signal input
rlabel metal2 s 8624 0 8680 400 6 wbs_adr_i[17]
port 356 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 wbs_adr_i[18]
port 357 nsew signal input
rlabel metal2 s 9520 0 9576 400 6 wbs_adr_i[19]
port 358 nsew signal input
rlabel metal2 s 1456 0 1512 400 6 wbs_adr_i[1]
port 359 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 wbs_adr_i[20]
port 360 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 wbs_adr_i[21]
port 361 nsew signal input
rlabel metal2 s 10864 0 10920 400 6 wbs_adr_i[22]
port 362 nsew signal input
rlabel metal2 s 11312 0 11368 400 6 wbs_adr_i[23]
port 363 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 wbs_adr_i[24]
port 364 nsew signal input
rlabel metal2 s 12208 0 12264 400 6 wbs_adr_i[25]
port 365 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 wbs_adr_i[26]
port 366 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 wbs_adr_i[27]
port 367 nsew signal input
rlabel metal2 s 13552 0 13608 400 6 wbs_adr_i[28]
port 368 nsew signal input
rlabel metal2 s 14000 0 14056 400 6 wbs_adr_i[29]
port 369 nsew signal input
rlabel metal2 s 1904 0 1960 400 6 wbs_adr_i[2]
port 370 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 wbs_adr_i[30]
port 371 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 wbs_adr_i[31]
port 372 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 wbs_adr_i[3]
port 373 nsew signal input
rlabel metal2 s 2800 0 2856 400 6 wbs_adr_i[4]
port 374 nsew signal input
rlabel metal2 s 3248 0 3304 400 6 wbs_adr_i[5]
port 375 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 wbs_adr_i[6]
port 376 nsew signal input
rlabel metal2 s 4144 0 4200 400 6 wbs_adr_i[7]
port 377 nsew signal input
rlabel metal2 s 4592 0 4648 400 6 wbs_adr_i[8]
port 378 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 wbs_adr_i[9]
port 379 nsew signal input
rlabel metal3 s 59600 18704 60000 18760 6 wbs_cyc_i
port 380 nsew signal input
rlabel metal2 s 15344 0 15400 400 6 wbs_dat_i[0]
port 381 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 wbs_dat_i[10]
port 382 nsew signal input
rlabel metal2 s 20272 0 20328 400 6 wbs_dat_i[11]
port 383 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_dat_i[12]
port 384 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 wbs_dat_i[13]
port 385 nsew signal input
rlabel metal2 s 21616 0 21672 400 6 wbs_dat_i[14]
port 386 nsew signal input
rlabel metal2 s 22064 0 22120 400 6 wbs_dat_i[15]
port 387 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 wbs_dat_i[16]
port 388 nsew signal input
rlabel metal2 s 22960 0 23016 400 6 wbs_dat_i[17]
port 389 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 wbs_dat_i[18]
port 390 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 wbs_dat_i[19]
port 391 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 wbs_dat_i[1]
port 392 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 wbs_dat_i[20]
port 393 nsew signal input
rlabel metal2 s 24752 0 24808 400 6 wbs_dat_i[21]
port 394 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 wbs_dat_i[22]
port 395 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 wbs_dat_i[23]
port 396 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 wbs_dat_i[24]
port 397 nsew signal input
rlabel metal2 s 26544 0 26600 400 6 wbs_dat_i[25]
port 398 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 wbs_dat_i[26]
port 399 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 wbs_dat_i[27]
port 400 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 wbs_dat_i[28]
port 401 nsew signal input
rlabel metal2 s 28336 0 28392 400 6 wbs_dat_i[29]
port 402 nsew signal input
rlabel metal2 s 16240 0 16296 400 6 wbs_dat_i[2]
port 403 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 wbs_dat_i[30]
port 404 nsew signal input
rlabel metal2 s 29232 0 29288 400 6 wbs_dat_i[31]
port 405 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 wbs_dat_i[3]
port 406 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 wbs_dat_i[4]
port 407 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 wbs_dat_i[5]
port 408 nsew signal input
rlabel metal2 s 18032 0 18088 400 6 wbs_dat_i[6]
port 409 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 wbs_dat_i[7]
port 410 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 wbs_dat_i[8]
port 411 nsew signal input
rlabel metal2 s 19376 0 19432 400 6 wbs_dat_i[9]
port 412 nsew signal input
rlabel metal3 s 59600 3920 60000 3976 6 wbs_dat_o[0]
port 413 nsew signal output
rlabel metal3 s 59600 8400 60000 8456 6 wbs_dat_o[10]
port 414 nsew signal output
rlabel metal3 s 59600 8848 60000 8904 6 wbs_dat_o[11]
port 415 nsew signal output
rlabel metal3 s 59600 9296 60000 9352 6 wbs_dat_o[12]
port 416 nsew signal output
rlabel metal3 s 59600 9744 60000 9800 6 wbs_dat_o[13]
port 417 nsew signal output
rlabel metal3 s 59600 10192 60000 10248 6 wbs_dat_o[14]
port 418 nsew signal output
rlabel metal3 s 59600 10640 60000 10696 6 wbs_dat_o[15]
port 419 nsew signal output
rlabel metal3 s 59600 11088 60000 11144 6 wbs_dat_o[16]
port 420 nsew signal output
rlabel metal3 s 59600 11536 60000 11592 6 wbs_dat_o[17]
port 421 nsew signal output
rlabel metal3 s 59600 11984 60000 12040 6 wbs_dat_o[18]
port 422 nsew signal output
rlabel metal3 s 59600 12432 60000 12488 6 wbs_dat_o[19]
port 423 nsew signal output
rlabel metal3 s 59600 4368 60000 4424 6 wbs_dat_o[1]
port 424 nsew signal output
rlabel metal3 s 59600 12880 60000 12936 6 wbs_dat_o[20]
port 425 nsew signal output
rlabel metal3 s 59600 13328 60000 13384 6 wbs_dat_o[21]
port 426 nsew signal output
rlabel metal3 s 59600 13776 60000 13832 6 wbs_dat_o[22]
port 427 nsew signal output
rlabel metal3 s 59600 14224 60000 14280 6 wbs_dat_o[23]
port 428 nsew signal output
rlabel metal3 s 59600 14672 60000 14728 6 wbs_dat_o[24]
port 429 nsew signal output
rlabel metal3 s 59600 15120 60000 15176 6 wbs_dat_o[25]
port 430 nsew signal output
rlabel metal3 s 59600 15568 60000 15624 6 wbs_dat_o[26]
port 431 nsew signal output
rlabel metal3 s 59600 16016 60000 16072 6 wbs_dat_o[27]
port 432 nsew signal output
rlabel metal3 s 59600 16464 60000 16520 6 wbs_dat_o[28]
port 433 nsew signal output
rlabel metal3 s 59600 16912 60000 16968 6 wbs_dat_o[29]
port 434 nsew signal output
rlabel metal3 s 59600 4816 60000 4872 6 wbs_dat_o[2]
port 435 nsew signal output
rlabel metal3 s 59600 17360 60000 17416 6 wbs_dat_o[30]
port 436 nsew signal output
rlabel metal3 s 59600 17808 60000 17864 6 wbs_dat_o[31]
port 437 nsew signal output
rlabel metal3 s 59600 5264 60000 5320 6 wbs_dat_o[3]
port 438 nsew signal output
rlabel metal3 s 59600 5712 60000 5768 6 wbs_dat_o[4]
port 439 nsew signal output
rlabel metal3 s 59600 6160 60000 6216 6 wbs_dat_o[5]
port 440 nsew signal output
rlabel metal3 s 59600 6608 60000 6664 6 wbs_dat_o[6]
port 441 nsew signal output
rlabel metal3 s 59600 7056 60000 7112 6 wbs_dat_o[7]
port 442 nsew signal output
rlabel metal3 s 59600 7504 60000 7560 6 wbs_dat_o[8]
port 443 nsew signal output
rlabel metal3 s 59600 7952 60000 8008 6 wbs_dat_o[9]
port 444 nsew signal output
rlabel metal3 s 59600 19152 60000 19208 6 wbs_stb_i
port 445 nsew signal input
rlabel metal3 s 59600 18256 60000 18312 6 wbs_we_i
port 446 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8594574
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/Multiplexer/runs/23_11_03_20_02/results/signoff/multiplexer.magic.gds
string GDS_START 344468
<< end >>

