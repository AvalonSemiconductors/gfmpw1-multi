* NGSPICE file created from blinker.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

.subckt blinker io_out[0] io_out[1] io_out[2] rst_n vdd vss wb_clk_i
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_3_3__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_501_ _127_ _142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_432_ PC\[1\] _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_13_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_895_ _038_ clknet_3_2__leaf_wb_clk_i LFSR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__780__C _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_878_ _021_ clknet_3_7__leaf_wb_clk_i counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_680_ _279_ _286_ _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_801_ _388_ _299_ _389_ _053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_732_ _298_ _333_ _334_ _335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_3_7__f_wb_clk_i clknet_0_wb_clk_i clknet_3_7__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_594_ counter\[15\] _223_ counter\[17\] counter\[16\] _224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_663_ _230_ _272_ _273_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_715_ _307_ _311_ _319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_646_ _260_ _261_ _262_ _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_577_ _111_ _142_ _204_ _072_ _209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_500_ _137_ _140_ _124_ _141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_431_ PC\[2\] _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_629_ _250_ _251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_894_ _037_ clknet_3_2__leaf_wb_clk_i LFSR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_6__f_wb_clk_i clknet_0_wb_clk_i clknet_3_6__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_877_ _020_ clknet_3_5__leaf_wb_clk_i counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_800_ clock_div\[8\] _357_ _365_ _389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_731_ _301_ LFSR\[3\] _334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_662_ counter\[17\] counter\[19\] counter\[18\] _267_ _273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_16_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_593_ counter\[14\] _223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_26_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_714_ _287_ _318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_576_ _126_ _199_ _200_ _208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_645_ _218_ _258_ counter\[13\] _262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_430_ PC\[3\] _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_628_ _229_ _250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_3_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_559_ _185_ _122_ _193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_5__f_wb_clk_i clknet_0_wb_clk_i clknet_3_5__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_893_ _036_ clknet_3_3__leaf_wb_clk_i OP_reg vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_28_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__890__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Left_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_876_ _019_ clknet_3_5__leaf_wb_clk_i counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_730_ _330_ _332_ _293_ _333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_661_ counter\[18\] _269_ counter\[19\] _272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_592_ counter\[6\] _219_ _221_ _222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_859_ _002_ clknet_3_0__leaf_wb_clk_i tune_ROM\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_713_ _299_ _314_ _317_ _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_575_ _201_ _203_ _207_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_644_ counter\[11\] counter\[13\] counter\[12\] _255_ _261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_15_Left_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_558_ _127_ _192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_627_ _246_ _247_ _249_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_489_ PC\[0\] _112_ _130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_4__f_wb_clk_i clknet_0_wb_clk_i clknet_3_4__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_0_Left_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_892_ _035_ clknet_3_6__leaf_wb_clk_i just_inc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Left_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_875_ _018_ clknet_3_5__leaf_wb_clk_i counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_660_ _231_ _271_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_591_ counter\[5\] _220_ counter\[7\] _221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_32_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_927_ _070_ clknet_3_2__leaf_wb_clk_i master_clk_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_789_ clock_div\[5\] _381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_858_ _001_ clknet_3_1__leaf_wb_clk_i tune_ROM\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_712_ LFSR\[0\] _316_ _296_ _317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3__f_wb_clk_i clknet_0_wb_clk_i clknet_3_3__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_643_ _229_ _260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_3_0__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_574_ _204_ _205_ _206_ _167_ _207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_5_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_557_ _157_ _189_ _190_ _191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_488_ _109_ _123_ _125_ _074_ _128_ _129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_626_ _248_ _249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_609_ net5 _234_ _237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_891_ _034_ clknet_3_0__leaf_wb_clk_i PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_874_ _017_ clknet_3_5__leaf_wb_clk_i counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__837__A1 _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_590_ counter\[4\] _220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_926_ _069_ clknet_3_2__leaf_wb_clk_i master_clk_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_788_ _379_ _380_ _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_3_2__f_wb_clk_i clknet_0_wb_clk_i clknet_3_2__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_12_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_857_ _000_ clknet_3_1__leaf_wb_clk_i tune_ROM\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__581__I _211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_711_ _315_ _316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_26_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_573_ _145_ _204_ _206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_642_ _218_ _258_ _259_ _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_909_ _052_ clknet_3_6__leaf_wb_clk_i clock_div\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_625_ counter\[7\] _245_ _248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_487_ _127_ _128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_556_ _185_ _182_ _188_ _190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_20_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_608_ net5 _234_ _236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_539_ _105_ _176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_890_ _033_ clknet_3_0__leaf_wb_clk_i PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_1__f_wb_clk_i clknet_0_wb_clk_i clknet_3_1__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_873_ _016_ clknet_3_5__leaf_wb_clk_i counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_925_ _068_ clknet_3_2__leaf_wb_clk_i master_clk_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_856_ _416_ _427_ _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_787_ clock_div\[4\] _375_ _376_ _380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_710_ _280_ _315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_641_ _218_ _258_ _251_ _259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_572_ _192_ _160_ _188_ _032_ _205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_27_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_908_ _051_ clknet_3_7__leaf_wb_clk_i clock_div\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_839_ _414_ _416_ _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__767__I _212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_486_ _071_ _126_ _127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_624_ counter\[7\] _245_ _247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_555_ _109_ _182_ _188_ _189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_20_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_538_ _134_ _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_607_ _230_ _235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_469_ PC\[1\] _100_ _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xclkbuf_3_0__f_wb_clk_i clknet_0_wb_clk_i clknet_3_0__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__860__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_872_ _015_ clknet_3_5__leaf_wb_clk_i counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__470__A1 _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_855_ master_clk_div\[6\] _426_ _427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_29_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_786_ _378_ _379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_924_ _067_ clknet_3_2__leaf_wb_clk_i master_clk_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_7_Left_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_571_ _114_ _119_ _148_ _139_ _204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_640_ _246_ _257_ _258_ _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_769_ _364_ _299_ _366_ _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_907_ _050_ clknet_3_6__leaf_wb_clk_i clock_div\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_838_ _415_ _416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_485_ PC\[4\] _096_ _126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_623_ _230_ _246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_554_ _118_ _124_ _188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_9_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_468_ net1 _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_606_ _233_ _216_ _234_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_537_ _031_ _173_ _174_ _175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_871_ _014_ clknet_3_5__leaf_wb_clk_i counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_23_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_854_ master_clk_div\[5\] _424_ _426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_923_ _066_ clknet_3_2__leaf_wb_clk_i master_clk_div\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_785_ clock_div\[4\] _375_ _378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__452__A2 _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_570_ _192_ _202_ _034_ _203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_768_ prev_clk_div _357_ _365_ _366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_906_ _049_ clknet_3_7__leaf_wb_clk_i clock_div\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_837_ _120_ _315_ _415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_699_ tune_ROM\[4\] _303_ _304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_484_ _124_ _125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_622_ _235_ _244_ _245_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_553_ _177_ _181_ _187_ _033_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_9_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_536_ _153_ _151_ _174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_467_ _108_ _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_605_ counter\[0\] counter\[1\] _234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_5_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_519_ _034_ _144_ _158_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_870_ _013_ clknet_3_5__leaf_wb_clk_i counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_853_ _416_ _425_ _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_784_ _375_ _377_ _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_922_ _065_ clknet_3_2__leaf_wb_clk_i master_clk_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_905_ _048_ clknet_3_7__leaf_wb_clk_i clock_div\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_836_ master_clk_div\[0\] _414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_767_ _212_ _365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_698_ tune_ROM\[3\] _303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_14_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_552_ _109_ _183_ _184_ _167_ _186_ _187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_483_ _106_ _110_ _113_ _124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_621_ counter\[5\] counter\[4\] counter\[6\] _239_ _245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_7_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_819_ rhythm_LFSR\[1\] rhythm_LFSR\[0\] _404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_604_ _232_ _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_535_ _172_ _173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_466_ net1 _101_ _107_ _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_33_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_5__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_449_ tempo_LFSR\[2\] tempo_LFSR\[1\] tempo_LFSR\[0\] _092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_518_ _150_ _156_ _157_ _158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_852_ _083_ _424_ _425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_783_ clock_div\[3\] _374_ _376_ _377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_921_ _064_ clknet_3_2__leaf_wb_clk_i master_clk_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_904_ _047_ clknet_3_6__leaf_wb_clk_i clock_div\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_766_ clock_div\[8\] _364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_697_ _292_ _302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__830__A1 _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_835_ _233_ _413_ _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_620_ counter\[6\] _242_ _244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_551_ _167_ _185_ _122_ _152_ _186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_749_ LFSR\[4\] _316_ _349_ _342_ _350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_818_ _403_ _056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_482_ _114_ _031_ _122_ _123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_603_ _120_ _232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_534_ _110_ _111_ _130_ _172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_465_ _074_ _106_ _095_ _073_ _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_33_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_517_ _105_ _157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_448_ tempo_LFSR\[3\] _091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_851_ _415_ _423_ _424_ _068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_782_ _295_ _376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_920_ _063_ clknet_3_4__leaf_wb_clk_i net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_27_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Left_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_765_ _318_ _362_ _363_ _043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_696_ _300_ _301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_903_ _046_ clknet_3_6__leaf_wb_clk_i clock_div\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_17_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_834_ net2 _228_ _413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_817_ rhythm_LFSR\[2\] _390_ _402_ _342_ _403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_13_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_550_ _108_ _185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_481_ _099_ _120_ _121_ _122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_748_ just_rst _288_ _287_ _348_ _349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_679_ just_inc _283_ _285_ _286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__567__A1 PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_14_Left_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_533_ _168_ _171_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_602_ counter\[0\] _231_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_464_ _075_ _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_447_ _088_ rhythm_LFSR\[2\] _089_ _080_ _090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_0_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_516_ _146_ _154_ _155_ _142_ _156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_36_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_850_ master_clk_div\[4\] _421_ _424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_781_ clock_div\[3\] _374_ _375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_28_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_764_ LFSR\[6\] _357_ _296_ _363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_25_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_902_ _045_ clknet_3_3__leaf_wb_clk_i clock_div\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_833_ _301_ _299_ _328_ _062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_695_ _081_ _300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__889__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_480_ _106_ _100_ _121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_747_ _292_ _347_ _348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_816_ _394_ _401_ _402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_678_ _284_ _285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_601_ _230_ _231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_463_ _105_ _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_10_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_532_ _157_ _169_ _170_ _171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_33_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_446_ rhythm_LFSR\[1\] rhythm_LFSR\[0\] _089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_0_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_515_ _146_ _140_ _119_ _155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__458__A1 PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_429_ PC\[4\] _072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_780_ _372_ _373_ _374_ _233_ _047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xinput1 rst_n net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_901_ _044_ clknet_3_3__leaf_wb_clk_i prev_clk_div vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_763_ _302_ _359_ _361_ _362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_694_ _298_ _299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_832_ _091_ _283_ _285_ _412_ _232_ _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_6_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_746_ _308_ _345_ _346_ _347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_815_ just_rst rhythm_LFSR\[3\] tune_ROM\[0\] _400_ _401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_13_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_677_ _093_ _282_ _284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_2__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_600_ _229_ _230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_462_ _104_ _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_531_ _072_ _159_ _136_ _170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_4_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_729_ _331_ _332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_514_ _132_ _147_ _152_ _030_ _154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_445_ rhythm_LFSR\[3\] _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__724__I _212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_428_ net1 _071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_900_ _043_ clknet_3_3__leaf_wb_clk_i LFSR\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_693_ _280_ _298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_762_ _351_ _337_ _360_ _302_ _361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_831_ _409_ tempo_LFSR\[0\] _412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_745_ _320_ _306_ _322_ _346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_814_ _391_ _400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_676_ _282_ _283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_13_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_461_ _071_ _097_ _103_ _104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_530_ _109_ _147_ _142_ _125_ _169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_728_ _307_ _303_ _320_ tune_ROM\[2\] _331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_18_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_659_ counter\[18\] _269_ _271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_444_ _086_ _087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_513_ _153_ _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_761_ _351_ _306_ _360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_830_ _233_ _411_ _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_692_ OP_reg _294_ _297_ _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_6_Left_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_32_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_744_ _304_ _344_ _345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_813_ _399_ _055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_675_ _281_ _090_ _282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_460_ _098_ _101_ _102_ _103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_727_ _304_ _306_ _308_ _330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_658_ _260_ _269_ _270_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_14_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_589_ counter\[10\] _217_ counter\[13\] _218_ _219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XPHY_EDGE_ROW_35_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_443_ master_clk_div\[1\] master_clk_div\[0\] _084_ _085_ _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_512_ _138_ _153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__606__A1 _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__859__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_760_ LFSR\[1\] LFSR\[0\] _359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_691_ OP_reg _294_ _296_ _297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_889_ _032_ clknet_3_0__leaf_wb_clk_i PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_674_ _082_ _280_ _281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_743_ _321_ _312_ _344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_812_ rhythm_LFSR\[1\] _390_ _398_ _342_ _399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_36_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_726_ _329_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_657_ counter\[17\] _267_ _270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_588_ counter\[12\] _218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_442_ master_clk_div\[3\] master_clk_div\[2\] _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_511_ _151_ _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_709_ _301_ LFSR\[1\] _302_ _313_ _314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_690_ _295_ _296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_888_ _031_ clknet_3_1__leaf_wb_clk_i PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_811_ _394_ _397_ _398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_742_ _343_ _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_673_ _087_ _280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_725_ LFSR\[1\] _318_ _327_ _328_ _329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_656_ counter\[17\] _267_ _269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_587_ counter\[11\] _217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_441_ master_clk_div\[4\] _083_ master_clk_div\[6\] _084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_510_ _115_ _116_ _113_ _117_ _151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_708_ _304_ _306_ _309_ _312_ _313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_639_ counter\[11\] _255_ _258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__439__B _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_887_ _030_ clknet_3_1__leaf_wb_clk_i PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_22_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_741_ LFSR\[3\] _316_ _341_ _342_ _343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_810_ _300_ rhythm_LFSR\[2\] _391_ _396_ _397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_672_ _232_ _279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_724_ _212_ _328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_655_ _267_ _268_ _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_586_ counter\[0\] counter\[1\] _216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_4_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_440_ master_clk_div\[5\] _083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_707_ _310_ _311_ _312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_638_ counter\[11\] _255_ _257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_569_ _132_ _160_ _152_ _140_ _202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_7__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_886_ _029_ clknet_3_1__leaf_wb_clk_i PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_26_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_10_Left_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_740_ _295_ _342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_671_ _231_ _278_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_869_ _012_ clknet_3_5__leaf_wb_clk_i counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_723_ _298_ _325_ _326_ _327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_654_ counter\[16\] _265_ _251_ _268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_585_ counter\[8\] counter\[9\] _215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_4_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Left_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_706_ tune_ROM\[2\] _303_ _311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_637_ _246_ _255_ _256_ _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__689__I _212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_568_ _174_ _199_ _200_ _145_ _201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_10_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_499_ _139_ _140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_885_ _028_ clknet_3_7__leaf_wb_clk_i counter\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_670_ counter\[22\] _277_ _278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_799_ _078_ _079_ _388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_21_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_868_ _011_ clknet_3_5__leaf_wb_clk_i counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__862__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_722_ _301_ LFSR\[2\] _326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_653_ counter\[15\] counter\[14\] counter\[16\] _261_ _267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_584_ counter\[3\] net5 _213_ _214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_4_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__490__A1 _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_705_ tune_ROM\[2\] tune_ROM\[3\] _310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_567_ PC\[3\] _174_ _200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_498_ _138_ _139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_636_ counter\[10\] _254_ _256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_619_ _235_ _242_ _243_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_22_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_884_ _027_ clknet_3_7__leaf_wb_clk_i counter\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_798_ _279_ _387_ _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_867_ _010_ clknet_3_4__leaf_wb_clk_i counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_721_ _293_ _324_ _325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_652_ _260_ _265_ _266_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_11_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_583_ counter\[19\] counter\[18\] _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_10_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_919_ _062_ clknet_3_3__leaf_wb_clk_i just_rst vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_4_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_704_ _307_ _308_ _309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_497_ _071_ _111_ _138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__481__A2 _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_635_ counter\[7\] counter\[10\] _215_ _245_ _255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_566_ _132_ _147_ _185_ _199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_618_ _220_ _240_ counter\[5\] _243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_549_ _030_ _031_ _114_ _184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_883_ _026_ clknet_3_7__leaf_wb_clk_i counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_866_ _009_ clknet_3_4__leaf_wb_clk_i counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_797_ clock_div\[7\] _385_ _387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_35_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_720_ _308_ _310_ _319_ _323_ _324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_651_ counter\[15\] _264_ _266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_582_ _071_ _212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_849_ master_clk_div\[4\] _421_ _423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_918_ _061_ clknet_3_4__leaf_wb_clk_i tempo_LFSR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_703_ tune_ROM\[5\] _308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_565_ _191_ _196_ _198_ _192_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_634_ _246_ _253_ _254_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_496_ _099_ _137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_17_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_4__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_617_ counter\[5\] _220_ _240_ _242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_479_ _115_ _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_548_ _176_ _182_ _183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Left_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_882_ _025_ clknet_3_4__leaf_wb_clk_i counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__430__I PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_5_Left_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_796_ _383_ _384_ _386_ _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_865_ _008_ clknet_3_4__leaf_wb_clk_i net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_31_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_650_ counter\[15\] _264_ _265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_848_ _415_ _421_ _422_ _067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_779_ clock_div\[2\] clock_div\[1\] _367_ _087_ _374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_917_ _060_ clknet_3_4__leaf_wb_clk_i tempo_LFSR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_581_ _211_ net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_702_ tune_ROM\[4\] _307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_495_ _134_ _135_ _136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_633_ _215_ _248_ _254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_564_ _176_ _122_ _197_ _180_ _173_ _198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_478_ _119_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_547_ _137_ _153_ _118_ _172_ _182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_616_ _231_ _241_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_881_ _024_ clknet_3_4__leaf_wb_clk_i counter\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_795_ _376_ _385_ _386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_864_ _007_ clknet_3_4__leaf_wb_clk_i counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_580_ OP_reg just_inc _211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_916_ _059_ clknet_3_6__leaf_wb_clk_i tempo_LFSR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_847_ master_clk_div\[3\] _419_ _422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_778_ clock_div\[1\] _367_ _298_ _373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_701_ _305_ tune_ROM\[2\] _306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_632_ counter\[8\] _249_ counter\[9\] _253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_563_ _146_ _188_ _164_ _197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__457__A2 _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_494_ _116_ _117_ _135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_477_ _118_ _119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_615_ _220_ _240_ _241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_546_ _179_ _180_ _033_ _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__444__I _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_529_ _161_ _162_ _166_ _145_ _167_ _168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_18_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_880_ _023_ clknet_3_5__leaf_wb_clk_i counter\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_794_ clock_div\[6\] _381_ _378_ _385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_21_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_863_ _006_ clknet_3_4__leaf_wb_clk_i counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_11_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_846_ master_clk_div\[3\] _419_ _421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_777_ clock_div\[2\] _372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_915_ _058_ clknet_3_4__leaf_wb_clk_i tempo_LFSR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_700_ tune_ROM\[4\] _305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__457__A3 _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_829_ tempo_LFSR\[2\] _282_ _284_ tempo_LFSR\[3\] _411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_562_ _192_ _195_ _196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_493_ _133_ _134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_631_ counter\[8\] _249_ _252_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_545_ _128_ _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_614_ _235_ _238_ _240_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_476_ _115_ _116_ _117_ _118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_9_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_459_ PC\[5\] _102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_528_ _104_ _167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_793_ _381_ _379_ _384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_862_ _005_ clknet_3_0__leaf_wb_clk_i tune_ROM\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_9_Left_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_845_ _416_ _419_ _420_ _066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_776_ _279_ _371_ _046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_914_ _057_ clknet_3_6__leaf_wb_clk_i rhythm_LFSR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_492_ _108_ _133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_630_ counter\[8\] _249_ _251_ _252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_561_ _174_ _193_ _194_ _176_ _195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_759_ _318_ _356_ _358_ _042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_828_ _279_ _410_ _059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_1__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_613_ _239_ _240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__835__A1 _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_475_ PC\[1\] _100_ _099_ _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_544_ _125_ _136_ _105_ _180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_527_ _163_ _164_ _165_ _166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_458_ PC\[3\] _099_ PC\[1\] _100_ _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_35_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_792_ clock_div\[6\] _383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_861_ _004_ clknet_3_0__leaf_wb_clk_i tune_ROM\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_25_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_844_ _417_ _414_ master_clk_div\[2\] _420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_775_ clock_div\[1\] _369_ _371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_913_ _056_ clknet_3_1__leaf_wb_clk_i rhythm_LFSR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__891__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_560_ _139_ _148_ _151_ _134_ _194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_491_ _131_ _132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_758_ LFSR\[5\] _357_ _296_ _358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_689_ _212_ _295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_827_ tempo_LFSR\[1\] _283_ _285_ tempo_LFSR\[2\] _410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__599__A1 _212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_543_ _159_ _160_ _178_ _029_ _152_ _030_ _179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_612_ counter\[0\] counter\[1\] counter\[3\] net3 _239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_474_ _074_ _106_ _095_ _116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_13_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_526_ _139_ _151_ _134_ _165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_457_ PC\[0\] _082_ _086_ _094_ _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_509_ _145_ _149_ _150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_791_ _381_ _379_ _382_ _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_860_ _003_ clknet_3_0__leaf_wb_clk_i tune_ROM\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_774_ _368_ _370_ _045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_843_ _417_ master_clk_div\[0\] master_clk_div\[2\] _419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_912_ _055_ clknet_3_0__leaf_wb_clk_i rhythm_LFSR\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_32_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_490_ _120_ _121_ _130_ _131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_3_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_757_ _315_ _357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_688_ _287_ _293_ _294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_826_ _408_ _283_ _285_ _409_ _232_ _058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_22_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_611_ counter\[3\] _236_ _238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_473_ net1 _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_542_ _148_ _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_809_ tune_ROM\[0\] tune_ROM\[1\] _396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_456_ PC\[2\] _099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_525_ _137_ _131_ _164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_439_ prev_clk_div _078_ _079_ _081_ _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_TAPCELL_ROW_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_508_ _146_ _147_ _148_ _140_ _149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_15_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_790_ _381_ _379_ _365_ _382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_842_ _417_ _414_ _418_ _065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_911_ _054_ clknet_3_3__leaf_wb_clk_i rhythm_LFSR\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_32_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_773_ _328_ _369_ _370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_756_ just_rst LFSR\[6\] _355_ _356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_687_ _292_ _293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_825_ tempo_LFSR\[1\] _409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_541_ _137_ _153_ _178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_610_ _235_ _236_ _237_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_472_ _110_ _111_ _113_ _114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_26_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_739_ _287_ _339_ _340_ _341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_808_ _390_ _393_ _395_ _054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__450__B _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_455_ _072_ _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_524_ _101_ _107_ _163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_18_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_438_ _080_ _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_507_ _110_ _113_ _148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_3_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_910_ _053_ clknet_3_3__leaf_wb_clk_i clock_div\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_29_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_772_ _367_ _315_ _369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_841_ _417_ _414_ _295_ _418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_755_ _351_ _352_ _354_ _302_ _355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_824_ tempo_LFSR\[0\] _408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_686_ _081_ _291_ _292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_540_ _159_ _165_ _175_ _032_ _176_ _177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_471_ PC\[0\] _112_ _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_738_ _300_ LFSR\[4\] _340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_807_ rhythm_LFSR\[0\] _394_ _365_ _395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_669_ counter\[21\] _274_ _277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_16_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_454_ PC\[5\] _072_ _096_ _097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_523_ _125_ _136_ _162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_18_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Left_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_437_ just_rst _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_506_ _135_ _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_6_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_771_ _367_ _316_ _368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_840_ master_clk_div\[1\] _417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__861__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Left_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_823_ _407_ _057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_685_ LFSR\[6\] _288_ _289_ _290_ _291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__695__I _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_754_ _351_ _353_ _311_ _354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_737_ _293_ _338_ _339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_806_ _281_ _394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_668_ counter\[21\] _274_ _276_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_599_ _212_ _228_ _229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_470_ _082_ _087_ _094_ _112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_13_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_522_ _159_ _160_ _128_ _161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_453_ _073_ _074_ _075_ _095_ _096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_33_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__674__A1 _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput2 net2 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_436_ clock_div\[8\] _076_ _077_ _079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_23_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_6__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_505_ _133_ _146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_770_ clock_div\[0\] _367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_899_ _042_ clknet_3_3__leaf_wb_clk_i LFSR\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_684_ LFSR\[1\] LFSR\[0\] _290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_753_ _307_ _310_ _353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_822_ rhythm_LFSR\[3\] _390_ _406_ _376_ _407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_16_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_736_ _309_ _337_ _338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_805_ rhythm_LFSR\[1\] _391_ _392_ _393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_667_ counter\[21\] _274_ _250_ _276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_598_ _214_ _215_ _216_ _227_ _228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_6_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_521_ _133_ _135_ _160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_452_ PC\[0\] _082_ _087_ _094_ _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_719_ _320_ _322_ _323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput3 net5 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_2_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_435_ _076_ _077_ clock_div\[8\] _078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_504_ _128_ _145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__912__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_898_ _041_ clknet_3_2__leaf_wb_clk_i LFSR\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_683_ LFSR\[4\] LFSR\[3\] LFSR\[2\] _289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_752_ _321_ _303_ _352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_821_ tune_ROM\[0\] _392_ _405_ _394_ _406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_735_ _321_ _310_ _337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_666_ _274_ _275_ _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_804_ tune_ROM\[1\] _391_ _392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_597_ _222_ _226_ _227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_520_ _114_ _159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_27_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_718_ _321_ _311_ _322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_649_ _260_ _263_ _264_ _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_451_ _090_ _093_ _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xoutput4 net4 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_2_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_434_ clock_div\[7\] clock_div\[6\] clock_div\[2\] clock_div\[1\] _077_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_23_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_503_ _129_ _143_ _144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_897_ _040_ clknet_3_2__leaf_wb_clk_i LFSR\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_682_ LFSR\[5\] _288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_751_ _320_ _351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_820_ _300_ _089_ _404_ _405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_8_Left_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__603__I _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout5 net3 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__686__A1 _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_734_ _336_ _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_665_ counter\[20\] _273_ _251_ _275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_596_ counter\[22\] _224_ _225_ _226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_803_ _090_ _391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_450_ _091_ _092_ _081_ _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_717_ tune_ROM\[4\] _321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_648_ counter\[14\] _261_ _264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_579_ _034_ _208_ _210_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_433_ clock_div\[5\] clock_div\[4\] clock_div\[3\] clock_div\[0\] _076_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_9_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_502_ _132_ _136_ _141_ _142_ _143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_31_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_896_ _039_ clknet_3_2__leaf_wb_clk_i LFSR\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_750_ _350_ _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_681_ _280_ _287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_879_ _022_ clknet_3_7__leaf_wb_clk_i counter\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_733_ LFSR\[2\] _318_ _335_ _328_ _336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_26_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_664_ counter\[20\] _273_ _274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_595_ counter\[21\] counter\[20\] _225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_802_ _281_ _390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_716_ tune_ROM\[5\] _320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_647_ counter\[14\] _261_ _263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_578_ _033_ _204_ _209_ _032_ _157_ _210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
.ends

