* NGSPICE file created from wrapped_ay8913.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

.subckt wrapped_ay8913 custom_settings[0] custom_settings[1] io_in_1[0] io_in_1[1]
+ io_in_1[2] io_in_1[3] io_in_1[4] io_in_1[5] io_in_1[6] io_in_1[7] io_in_2[0] io_in_2[1]
+ io_out[10] io_out[11] io_out[17] io_out[18] io_out[19] io_out[20] io_out[21] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] rst_n vdd vss wb_clk_i io_out[1] io_out[16]
+ io_out[15] io_out[0] io_out[14] io_out[13] io_out[12] io_out[22]
X_2106_ _0056_ clknet_leaf_22_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2037_ tt_um_rejunity_ay8913.pwm_A.accumulator\[6\] _0597_ _0593_ _0601_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_52_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1684__A1 _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1270_ net5 _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1606_ _0254_ _0255_ _0248_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1537_ _1003_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1468_ tt_um_rejunity_ay8913.envelope_generator.period\[8\] _0943_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1399_ _0840_ _0872_ _0883_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_28_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1322_ tt_um_rejunity_ay8913.pwm_B.accumulator\[8\] _0832_ _0833_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1253_ _0786_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1409__A1 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1184_ _0734_ _0739_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1887__A1 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1940_ tt_um_rejunity_ay8913.tone_A_generator.counter\[5\] _0536_ _0538_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1871_ _0473_ _0480_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1305_ _0819_ _0820_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1236_ _0767_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1098_ _0670_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1167_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\] _0726_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2070_ _0020_ clknet_leaf_37_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1923_ _0492_ _0525_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1854_ _0408_ _0307_ _0425_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1785_ _0371_ _0403_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2199_ _0149_ clknet_leaf_7_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.hold
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1219_ _0719_ tt_um_rejunity_ay8913.pwm_C.accumulator\[8\] _0760_ _0762_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2268_ _0218_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_14_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_14_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_13_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _0895_ tt_um_rejunity_ay8913.envelope_attack _0893_ tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
+ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2122_ _0072_ clknet_leaf_37_wb_clk_i net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2053_ _0003_ clknet_leaf_31_wb_clk_i tt_um_rejunity_ay8913.noise_generator.period\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1906_ tt_um_rejunity_ay8913.tone_A_generator.period\[5\] _0509_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1768_ _0732_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1837_ _0451_ _0452_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1699_ tt_um_rejunity_ay8913.tone_C_generator.counter\[10\] _0325_ _0326_ tt_um_rejunity_ay8913.tone_C_generator.counter\[9\]
+ _0327_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_35_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput20 net20 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1622_ _0244_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1553_ _0942_ _1011_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1484_ _0958_ _0945_ _0941_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_52_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2105_ _0055_ clknet_leaf_22_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2036_ _0599_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1536_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\] _1002_ _1003_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1605_ tt_um_rejunity_ay8913.noise_generator.lfsr\[6\] _0250_ _0255_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1467_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\] _0942_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1398_ _0671_ tt_um_rejunity_ay8913.envelope_generator.period\[12\] _0873_ _0883_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1372__A1 _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2019_ _0588_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1115__A1 _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1666__A2 _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1106__A1 _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1321_ tt_um_rejunity_ay8913.pwm_B.accumulator\[7\] _0826_ _0832_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1252_ _0630_ _0784_ _0785_ tt_um_rejunity_ay8913.tone_B_generator.period\[8\] _0786_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_24_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1183_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\] _0727_ _0736_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\]
+ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_19_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1345__A1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1519_ _0990_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1103__I _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_39_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_39_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1870_ _0415_ _0479_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1166_ _0715_ _0725_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1304_ tt_um_rejunity_ay8913.pwm_B.accumulator\[3\] _0817_ _0753_ _0820_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1235_ _0764_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1097_ net13 _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1566__A1 _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1999_ _0835_ _0571_ _0575_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1768__I _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1922_ _0524_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_44_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1853_ _0425_ _0408_ _0986_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1784_ _0323_ _0401_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_12_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2198_ _0148_ clknet_leaf_8_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1218_ tt_um_rejunity_ay8913.pwm_C.accumulator\[8\] _0760_ _0761_ _0038_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1149_ _0699_ _0712_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2267_ _0217_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1778__A1 _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2121_ _0071_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2052_ _0002_ clknet_leaf_31_wb_clk_i tt_um_rejunity_ay8913.noise_generator.period\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1905_ tt_um_rejunity_ay8913.tone_A_generator.counter\[4\] _0497_ _0504_ _0506_ _0507_
+ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_29_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1698_ _0322_ tt_um_rejunity_ay8913.tone_C_generator.period\[11\] _0327_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1767_ _0390_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1836_ _0449_ tt_um_rejunity_ay8913.tone_B_generator.period\[10\] _0452_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input11_I io_in_2[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput21 net21 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1552_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\] _1015_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1621_ _0265_ _0266_ _0259_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1483_ _0942_ _0875_ _0943_ _0944_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2104_ _0054_ clknet_leaf_22_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input3_I io_in_1[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2035_ tt_um_rejunity_ay8913.pwm_A.accumulator\[6\] _0597_ _0599_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_32_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1819_ tt_um_rejunity_ay8913.tone_B_generator.counter\[3\] _0435_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1535_ _0996_ _1001_ _1002_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1604_ tt_um_rejunity_ay8913.noise_generator.lfsr\[7\] _0245_ _0254_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1466_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\] _0880_ _0878_
+ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\] _0941_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1397_ _0675_ _0880_ _0881_ _0882_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_38_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2018_ _0778_ _0584_ _0585_ tt_um_rejunity_ay8913.envelope_generator.period\[6\]
+ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_19_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1320_ _0659_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_11_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1251_ _0732_ _0783_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1182_ _0734_ _0738_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_19_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_9_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_9_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1449_ tt_um_rejunity_ay8913.envelope_generator.period\[2\] _0924_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1518_ _0980_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1303_ tt_um_rejunity_ay8913.pwm_B.accumulator\[3\] _0817_ _0819_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1096_ _0668_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1165_ net19 _0722_ _0724_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\] _0725_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1234_ _0772_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1263__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1998_ _0686_ _0567_ _0856_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1921_ _0670_ _0523_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1852_ _0464_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1783_ _0402_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1362__C _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2266_ _0216_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1079_ _0632_ _0655_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1217_ tt_um_rejunity_ay8913.pwm_C.accumulator\[8\] _0760_ _0707_ _0761_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1148_ _0706_ _0704_ _0709_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2197_ _0147_ clknet_leaf_31_wb_clk_i tt_um_rejunity_ay8913.noise_generator.tone.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1778__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_7_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_23_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_23_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2120_ _0070_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2051_ _0001_ clknet_leaf_32_wb_clk_i tt_um_rejunity_ay8913.noise_generator.period\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1904_ _0505_ tt_um_rejunity_ay8913.tone_A_generator.period\[3\] _0507_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1835_ _0448_ tt_um_rejunity_ay8913.tone_B_generator.period\[11\] _0451_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1697_ tt_um_rejunity_ay8913.tone_C_generator.period\[9\] _0326_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1766_ _0884_ _0386_ _0388_ _0389_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2249_ _0199_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput22 net22 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_14_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1551_ _1007_ _1014_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1482_ _0955_ _0956_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1620_ tt_um_rejunity_ay8913.noise_generator.lfsr\[10\] _0261_ _0266_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2103_ _0053_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2034_ _0597_ _0598_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1818_ tt_um_rejunity_ay8913.tone_B_generator.period\[3\] _0434_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1749_ _0339_ _0372_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_8_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1534_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\] tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\]
+ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\] _0995_ _1002_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1465_ _0938_ tt_um_rejunity_ay8913.envelope_generator.period\[12\] _0939_ _0940_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1603_ _0252_ _0253_ _0248_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2017_ _0587_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1396_ _0686_ _0876_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_36_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1181_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\] _0727_ _0736_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\]
+ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_19_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1250_ _0783_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1517_ _0988_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1448_ tt_um_rejunity_ay8913.envelope_generator.period\[3\] _0923_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1379_ _0869_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1400__I _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2049__A1 _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1233_ _0648_ _0765_ _0768_ tt_um_rejunity_ay8913.tone_C_generator.period\[3\] _0772_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1302_ _0817_ _0818_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1095_ _0655_ _0667_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1164_ _0723_ _0721_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1997_ _0631_ _0571_ _0574_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1920_ _0519_ _0521_ _0522_ _0981_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_21_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1851_ _0466_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1782_ _0371_ _0400_ _0401_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_46_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1216_ _0689_ _0759_ _0760_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2196_ _0146_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2265_ _0215_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1078_ tt_um_rejunity_ay8913.latched_register\[1\] _0654_ _0655_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1147_ _0710_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_51_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2050_ _0000_ clknet_leaf_32_wb_clk_i tt_um_rejunity_ay8913.noise_generator.period\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1903_ _0505_ tt_um_rejunity_ay8913.tone_A_generator.period\[3\] tt_um_rejunity_ay8913.tone_A_generator.period\[2\]
+ _0498_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_32_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1765_ tt_um_rejunity_ay8913.tone_C_generator.counter\[5\] tt_um_rejunity_ay8913.tone_C_generator.counter\[4\]
+ _0378_ _0379_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1834_ _0448_ tt_um_rejunity_ay8913.tone_B_generator.period\[11\] tt_um_rejunity_ay8913.tone_B_generator.period\[10\]
+ _0449_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1696_ tt_um_rejunity_ay8913.tone_C_generator.period\[10\] _0325_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2179_ _0129_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2248_ _0198_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1481_ _0912_ tt_um_rejunity_ay8913.envelope_generator.period\[7\] _0956_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1550_ _1013_ _1011_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2102_ _0052_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2033_ tt_um_rejunity_ay8913.pwm_A.accumulator\[5\] _0595_ _0593_ _0598_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1817_ tt_um_rejunity_ay8913.tone_B_generator.period\[4\] _0433_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1748_ _0375_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1679_ _0313_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1127__A1 _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1602_ tt_um_rejunity_ay8913.noise_generator.lfsr\[5\] _0250_ _0253_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1533_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\] _1000_ _1001_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1464_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\] _0880_ _0939_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1395_ _0871_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2016_ net8 _0584_ _0585_ tt_um_rejunity_ay8913.envelope_generator.period\[5\] _0587_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1223__I _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1339__A1 _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1180_ _0734_ _0737_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_19_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1516_ _0899_ _0982_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1447_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\] _0922_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1378_ _0650_ _0861_ _0863_ tt_um_rejunity_ay8913.noise_disable_B _0869_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1750__A1 _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1291__C _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_17_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_17_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1232_ _0771_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1301_ tt_um_rejunity_ay8913.pwm_B.accumulator\[2\] _0623_ _0753_ _0818_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1094_ tt_um_rejunity_ay8913.latched_register\[3\] tt_um_rejunity_ay8913.latched_register\[2\]
+ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1163_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\] _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1996_ _0683_ _0568_ _0856_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1411__I _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1962__A1 _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1781_ _0352_ _0398_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1850_ _0409_ _0465_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_46_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1146_ _0706_ _0709_ _0703_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1215_ tt_um_rejunity_ay8913.pwm_C.accumulator\[6\] tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
+ _0755_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2195_ _0145_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2264_ _0214_ clknet_leaf_2_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1077_ _0653_ _0635_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1979_ _0561_ _0562_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1902_ tt_um_rejunity_ay8913.tone_A_generator.counter\[3\] _0505_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_32_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_32_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_32_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_52_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1764_ _0344_ _0387_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1833_ tt_um_rejunity_ay8913.tone_B_generator.counter\[10\] _0449_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1695_ _0322_ tt_um_rejunity_ay8913.tone_C_generator.period\[11\] tt_um_rejunity_ay8913.tone_C_generator.period\[10\]
+ _0323_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2247_ _0197_ clknet_leaf_2_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2178_ _0128_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1129_ _0695_ _0694_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1090__A1 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1480_ _0940_ _0941_ _0946_ _0954_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2032_ tt_um_rejunity_ay8913.pwm_A.accumulator\[5\] _0595_ _0597_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2101_ _0051_ clknet_leaf_24_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1816_ _0427_ _0430_ _0431_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1678_ _0699_ _0301_ _0311_ _0312_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1747_ _0371_ _0372_ _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1669__A3 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1532_ _0996_ _0999_ _1000_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1601_ tt_um_rejunity_ay8913.noise_generator.lfsr\[6\] _0245_ _0252_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I custom_settings[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1463_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\] _0938_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1394_ tt_um_rejunity_ay8913.envelope_generator.period\[11\] _0880_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_38_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2015_ _0586_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1520__A2 _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1284__A1 _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1511__A2 _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1515_ _0983_ _0987_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1446_ _0918_ tt_um_rejunity_ay8913.envelope_generator.period\[5\] tt_um_rejunity_ay8913.envelope_generator.period\[4\]
+ _0920_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1377_ _0868_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1162_ _0721_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1231_ _0646_ _0765_ _0768_ tt_um_rejunity_ay8913.tone_C_generator.period\[2\] _0771_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1300_ tt_um_rejunity_ay8913.pwm_B.accumulator\[2\] _0623_ _0817_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1093_ _0665_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1995_ _0633_ _0571_ _0573_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_30_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1429_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\] _0905_ _0907_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1848__B _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1780_ _0352_ _0398_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2263_ _0213_ clknet_leaf_17_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1145_ tt_um_rejunity_ay8913.pwm_master.accumulator\[7\] _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1214_ tt_um_rejunity_ay8913.pwm_C.accumulator\[6\] _0756_ tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
+ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2194_ _0144_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1076_ tt_um_rejunity_ay8913.latched_register\[0\] _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ tt_um_rejunity_ay8913.clk_counter\[4\] _0558_ _0559_ _0562_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_2_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1332__I _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1901_ _0498_ tt_um_rejunity_ay8913.tone_A_generator.period\[2\] _0501_ _0503_ _0504_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_16_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1832_ tt_um_rejunity_ay8913.tone_B_generator.counter\[11\] _0448_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1694_ tt_um_rejunity_ay8913.tone_C_generator.counter\[10\] _0323_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1763_ tt_um_rejunity_ay8913.tone_C_generator.counter\[4\] _0378_ _0379_ _0387_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2246_ _0196_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2177_ _0127_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1128_ _0690_ _0626_ _0627_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1059_ _0640_ _0637_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput14 net14 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2100_ _0050_ clknet_leaf_24_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2031_ _0595_ _0596_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1815_ _0423_ tt_um_rejunity_ay8913.tone_B_generator.period\[2\] _0431_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_40_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1677_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\] _0309_ _0312_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1746_ _0319_ _0373_ _0330_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2229_ _0179_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1610__I _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1531_ _0919_ _0998_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1462_ _0916_ _0936_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1057__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1600_ _0249_ _0251_ _0248_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1393_ _0675_ _0878_ _0872_ _0879_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_38_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2014_ _0650_ _0584_ _0585_ tt_um_rejunity_ay8913.envelope_generator.period\[4\]
+ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_9_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1729_ _0353_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1445_ _0919_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1514_ _0929_ _0986_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1376_ _0800_ _0862_ _0864_ tt_um_rejunity_ay8913.noise_disable_A _0868_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_2_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_2_2__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1161_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\] tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
+ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1230_ _0770_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_26_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_26_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1092_ net3 _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1994_ _0677_ _0568_ _0829_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1428_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\] _0905_ _0906_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1359_ _0857_ _0722_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2262_ _0212_ clknet_leaf_15_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1166__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1213_ tt_um_rejunity_ay8913.pwm_C.accumulator\[6\] _0756_ _0758_ _0036_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_35_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1144_ _0706_ _0704_ _0708_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2193_ _0143_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1075_ _0652_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1977_ tt_um_rejunity_ay8913.clk_counter\[4\] _0558_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1396__A1 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1900_ tt_um_rejunity_ay8913.tone_A_generator.counter\[0\] _0502_ _0500_ tt_um_rejunity_ay8913.tone_A_generator.counter\[1\]
+ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1831_ _0416_ _0442_ _0446_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1926__A3 _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1693_ tt_um_rejunity_ay8913.tone_C_generator.counter\[11\] _0322_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1762_ _0991_ _0385_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1139__A1 _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2245_ _0195_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_27_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2176_ _0126_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_11_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1127_ _0689_ _0693_ _0694_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1058_ _0639_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1378__A1 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput15 net15 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2030_ tt_um_rejunity_ay8913.pwm_A.accumulator\[4\] _0592_ _0593_ _0596_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1814_ tt_um_rejunity_ay8913.tone_B_generator.counter\[0\] _0428_ _0429_ _0430_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1745_ _0981_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_40_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1676_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\] _0309_ _0311_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2159_ _0109_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2228_ _0178_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.tone_B vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1202__B _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1771__A1 _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1530_ _0919_ _0998_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1461_ _0913_ _0917_ _0921_ _0934_ _0935_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1392_ _0683_ _0876_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1762__A1 _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2013_ _0578_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1073__I _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1957__B _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1728_ _0346_ _0349_ _0351_ _0356_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_13_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1659_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[4\] _0298_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1158__I _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1444_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\] _0919_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1375_ _0867_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1513_ _0980_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1160_ _0720_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1091_ _0664_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1993_ _0653_ _0571_ _0572_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1427_ _0903_ _0904_ _0905_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1358_ _0856_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_41_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1289_ _0808_ _0810_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_21_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2261_ _0211_ clknet_leaf_15_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1212_ tt_um_rejunity_ay8913.pwm_C.accumulator\[6\] _0756_ _0707_ _0758_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2192_ _0142_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.noise_generator.signal_edge.signal
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1143_ _0706_ _0704_ _0707_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1074_ _0651_ _0637_ _0641_ tt_um_rejunity_ay8913.noise_generator.period\[4\] _0652_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1976_ _0558_ _0560_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1830_ _0445_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1761_ _0368_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1692_ _0980_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_10_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_10_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2244_ _0194_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2175_ _0125_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1126_ tt_um_rejunity_ay8913.pwm_master.accumulator\[2\] _0624_ _0691_ _0692_ _0694_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1057_ net13 _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1959_ _0655_ _0836_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput16 net16 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_54_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1853__A3 _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1813_ tt_um_rejunity_ay8913.tone_B_generator.counter\[1\] tt_um_rejunity_ay8913.tone_B_generator.period\[1\]
+ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1744_ tt_um_rejunity_ay8913.tone_C_generator.counter\[1\] tt_um_rejunity_ay8913.tone_C_generator.counter\[0\]
+ _0990_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1675_ _0303_ _0309_ _0310_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2158_ _0108_ clknet_leaf_12_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2089_ _0039_ clknet_leaf_37_wb_clk_i net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1109_ _0679_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2227_ _0177_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1771__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1287__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1460_ _0918_ tt_um_rejunity_ay8913.envelope_generator.period\[5\] _0935_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1514__A2 _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1391_ tt_um_rejunity_ay8913.envelope_generator.period\[10\] _0878_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_38_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1762__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2012_ _0576_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1278__A1 _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1727_ _0353_ _0355_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1658_ _0289_ tt_um_rejunity_ay8913.noise_generator.period\[3\] tt_um_rejunity_ay8913.noise_generator.period\[2\]
+ _0295_ _0296_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_13_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1589_ tt_um_rejunity_ay8913.noise_generator.lfsr\[2\] _0237_ _0243_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1174__I _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1512_ _0983_ _0148_ _0985_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1443_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\] _0918_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1374_ _0798_ _0862_ _0864_ tt_um_rejunity_ay8913.tone_disable_C _0867_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1968__B _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1423__A1 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2039__B _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output19_I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1090_ _0648_ _0657_ _0660_ tt_um_rejunity_ay8913.tone_C_generator.period\[11\] _0664_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_51_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1992_ _0629_ _0568_ _0829_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_35_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_35_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1426_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\] tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\]
+ _0898_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1357_ _0670_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1288_ _0809_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2260_ _0210_ clknet_leaf_22_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2191_ _0141_ clknet_leaf_5_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[16\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1211_ _0756_ _0757_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1142_ _0680_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1073_ _0650_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1311__B _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1975_ tt_um_rejunity_ay8913.clk_counter\[3\] _0557_ _0559_ _0560_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1409_ _0884_ _0889_ _0881_ _0890_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_38_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1357__I _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1760_ _0384_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1691_ _0319_ _0986_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2174_ _0124_ clknet_leaf_6_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.invert_output
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2243_ _0193_ clknet_leaf_2_wb_clk_i tt_um_rejunity_ay8913.envelope_B vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1125_ tt_um_rejunity_ay8913.pwm_master.accumulator\[2\] _0624_ _0691_ _0692_ _0693_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1092__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1056_ _0637_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1889_ _0491_ _0321_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1958_ tt_um_rejunity_ay8913.tone_A _0523_ _0548_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1267__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput17 net17 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2006__A1 _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1812_ tt_um_rejunity_ay8913.tone_B_generator.period\[0\] _0428_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1674_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\] _0306_ _0310_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1743_ _0369_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2226_ _0176_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2157_ _0107_ clknet_leaf_7_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2088_ _0038_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1039_ _0622_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1108_ net13 _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1390_ _0675_ _0875_ _0872_ _0877_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_54_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2011_ _0583_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1588_ tt_um_rejunity_ay8913.noise_generator.lfsr\[3\] _0233_ _0242_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1726_ _0354_ _0332_ _0347_ tt_um_rejunity_ay8913.tone_C_generator.counter\[6\] _0355_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1657_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\] _0294_ _0296_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2209_ _0159_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1442_ tt_um_rejunity_ay8913.envelope_generator.period\[6\] _0917_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1511_ tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal _0982_ _0985_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_10_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1373_ _0866_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1671__A2 _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1709_ tt_um_rejunity_ay8913.tone_C_generator.counter\[3\] _0336_ _0337_ tt_um_rejunity_ay8913.tone_C_generator.counter\[4\]
+ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1111__A1 _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_5_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_5_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1788__C _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1991_ _0567_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1425_ _0892_ _0898_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\]
+ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1356_ _0855_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1341__A1 _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1287_ _0718_ _0728_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_21_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1399__A1 _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1072_ net7 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2190_ _0140_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1323__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1141_ tt_um_rejunity_ay8913.pwm_master.accumulator\[6\] _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1210_ tt_um_rejunity_ay8913.pwm_C.accumulator\[5\] _0752_ _0753_ _0757_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1974_ _0698_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1408_ net10 _0873_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1339_ _0790_ _0843_ _0845_ tt_um_rejunity_ay8913.tone_A_generator.period\[0\] _0846_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1690_ tt_um_rejunity_ay8913.tone_C_generator.counter\[0\] _0319_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2242_ _0192_ clknet_leaf_3_wb_clk_i tt_um_rejunity_ay8913.amplitude_B\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2173_ _0123_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1055_ _0632_ _0636_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1124_ _0690_ _0626_ _0627_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1957_ tt_um_rejunity_ay8913.tone_A _0523_ _0391_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1888_ tt_um_rejunity_ay8913.tone_A_generator.counter\[0\] _0491_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1992__B _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput18 net18 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1774__A1 _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1811_ _0425_ _0426_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1673_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\] _0306_ _0309_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1742_ _0320_ _0370_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2225_ _0175_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2156_ _0106_ clknet_leaf_7_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.stop
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1107_ _0675_ _0676_ _0669_ _0678_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1038_ _0619_ _0620_ _0608_ tt_um_rejunity_ay8913.envelope_B _0621_ _0622_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2087_ _0037_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2010_ _0686_ _0577_ _0579_ tt_um_rejunity_ay8913.envelope_generator.period\[3\]
+ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_29_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1986__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1098__I _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1725_ tt_um_rejunity_ay8913.tone_C_generator.counter\[7\] _0354_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1587_ _0240_ _0241_ _0239_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1753__A4 _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1656_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\] _0294_ _0295_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2139_ _0089_ clknet_leaf_3_wb_clk_i tt_um_rejunity_ay8913.tone_disable_C vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2208_ _0158_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1441_ _0915_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1510_ _0984_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1372_ _0796_ _0862_ _0864_ tt_um_rejunity_ay8913.tone_disable_B _0866_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1120__A2 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1708_ tt_um_rejunity_ay8913.tone_C_generator.period\[4\] _0337_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1639_ _0278_ _0279_ _0715_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_18_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_54_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1990_ _0568_ _0570_ _0715_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_15_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1355_ _0780_ _0850_ _0851_ tt_um_rejunity_ay8913.tone_A_generator.period\[7\] _0855_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1424_ _0902_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1286_ _0730_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1140_ _0702_ _0700_ _0705_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1071_ _0649_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1973_ tt_um_rejunity_ay8913.clk_counter\[3\] _0557_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_7_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1407_ tt_um_rejunity_ay8913.envelope_generator.period\[15\] _0889_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1338_ _0844_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1269_ _0797_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2172_ _0122_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2241_ _0191_ clknet_leaf_14_wb_clk_i tt_um_rejunity_ay8913.tone_A vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1054_ _0633_ tt_um_rejunity_ay8913.latched_register\[0\] _0635_ _0636_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1123_ _0626_ _0627_ _0690_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1956_ _0520_ _0547_ _0533_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1887_ _0857_ _0489_ _0490_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_7_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput19 net19 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_54_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1810_ tt_um_rejunity_ay8913.tone_B_generator.period\[1\] _0426_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1741_ _0369_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1672_ _0303_ _0306_ _0308_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2155_ _0105_ clknet_leaf_8_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1106_ _0677_ _0672_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2224_ _0174_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1037_ tt_um_rejunity_ay8913.amplitude_B\[0\] tt_um_rejunity_ay8913.envelope_B tt_um_rejunity_ay8913.tone_disable_B
+ tt_um_rejunity_ay8913.tone_B _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_2086_ _0036_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1939_ tt_um_rejunity_ay8913.tone_A_generator.counter\[5\] _0510_ tt_um_rejunity_ay8913.tone_A_generator.counter\[3\]
+ _0531_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_31_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1508__A2 _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1986__A2 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1724_ _0352_ _0326_ _0333_ tt_um_rejunity_ay8913.tone_C_generator.counter\[8\] _0353_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1586_ tt_um_rejunity_ay8913.noise_generator.lfsr\[1\] _0237_ _0241_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1655_ _0291_ _0293_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1998__B _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2138_ _0088_ clknet_leaf_3_wb_clk_i tt_um_rejunity_ay8913.tone_disable_B vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2069_ _0019_ clknet_leaf_37_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2207_ _0157_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1665__A1 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1440_ _0912_ tt_um_rejunity_ay8913.envelope_generator.period\[7\] tt_um_rejunity_ay8913.envelope_generator.period\[6\]
+ _0914_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1371_ _0865_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_18_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1638_ tt_um_rejunity_ay8913.noise_generator.lfsr\[15\] _0272_ _0279_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1707_ tt_um_rejunity_ay8913.tone_C_generator.period\[3\] _0336_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1569_ tt_um_rejunity_ay8913.envelope_generator.hold tt_um_rejunity_ay8913.envelope_alternate
+ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_51_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_35_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1354_ _0854_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1423_ _0658_ tt_um_rejunity_ay8913.restart_envelope _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1285_ _0807_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_46_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_13_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_13_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_18_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1070_ _0648_ _0638_ _0642_ tt_um_rejunity_ay8913.noise_generator.period\[3\] _0649_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1972_ _0689_ _0556_ _0557_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_15_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1337_ _0766_ _0842_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1406_ _0884_ _0887_ _0881_ _0888_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1268_ _0796_ _0792_ _0794_ tt_um_rejunity_ay8913.tone_B_generator.period\[1\] _0797_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1199_ _0609_ _0614_ tt_um_rejunity_ay8913.pwm_C.accumulator\[2\] _0749_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1856__A4 _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2018__A1 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2171_ _0121_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2240_ _0190_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1122_ tt_um_rejunity_ay8913.pwm_master.accumulator\[3\] _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1053_ tt_um_rejunity_ay8913.active _0634_ net11 net13 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1955_ tt_um_rejunity_ay8913.tone_A_generator.counter\[10\] _0545_ _0547_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1886_ _0373_ _0463_ tt_um_rejunity_ay8913.tone_B _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1740_ _0321_ _0368_ _0640_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1671_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\] _0307_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\]
+ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input8_I io_in_1[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2154_ _0104_ clknet_leaf_8_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1105_ net4 _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2223_ _0173_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2085_ _0035_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1036_ tt_um_rejunity_ay8913.noise_disable_B _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1938_ _0527_ _0535_ _0536_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_31_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1869_ _0467_ _0478_ _0479_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_47_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1380__A1 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1986__A3 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_38_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_38_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1723_ tt_um_rejunity_ay8913.tone_C_generator.counter\[9\] _0352_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1654_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\] _0292_ _0290_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\]
+ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1585_ tt_um_rejunity_ay8913.noise_generator.lfsr\[2\] _0233_ _0240_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2206_ _0156_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2137_ _0087_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.tone_disable_A vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2068_ _0018_ clknet_leaf_37_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1353__A1 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1370_ _0790_ _0862_ _0864_ tt_um_rejunity_ay8913.tone_disable_A _0865_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1637_ tt_um_rejunity_ay8913.noise_generator.lfsr\[16\] _0244_ _0278_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1706_ _0334_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1499_ net2 _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1568_ _0947_ _0225_ _1007_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_1_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1422_ _0892_ _0898_ _0901_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1353_ _0778_ _0850_ _0851_ tt_um_rejunity_ay8913.tone_A_generator.period\[6\] _0854_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_38_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1284_ _0780_ _0802_ _0803_ tt_um_rejunity_ay8913.tone_B_generator.period\[7\] _0807_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_46_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1583__I _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1971_ tt_um_rejunity_ay8913.clk_counter\[0\] _0554_ tt_um_rejunity_ay8913.clk_counter\[2\]
+ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_15_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1405_ net9 _0873_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput1 custom_settings[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1336_ _0842_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1267_ net4 _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1198_ tt_um_rejunity_ay8913.pwm_C.accumulator\[2\] _0609_ _0614_ _0748_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_6_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2170_ _0120_ clknet_leaf_18_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1052_ net12 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1172__B _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1121_ _0659_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1954_ _0533_ _0546_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1885_ tt_um_rejunity_ay8913.tone_B _0373_ _0463_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1319_ tt_um_rejunity_ay8913.pwm_B.accumulator\[7\] _0827_ _0830_ _0070_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1759__A1 _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1998__A1 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1670_ _0990_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2222_ _0172_ clknet_leaf_21_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1104_ tt_um_rejunity_ay8913.tone_A_generator.period\[9\] _0676_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2153_ _0103_ clknet_leaf_7_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1035_ tt_um_rejunity_ay8913.noise_generator.lfsr\[0\] _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2084_ _0034_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1937_ _0510_ tt_um_rejunity_ay8913.tone_A_generator.counter\[3\] _0532_ _0536_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_31_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1868_ tt_um_rejunity_ay8913.tone_B_generator.counter\[5\] _0418_ _0435_ _0470_ _0479_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1799_ tt_um_rejunity_ay8913.tone_B_generator.counter\[6\] _0415_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_54_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_8_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_8_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1584_ _0234_ _0238_ _0239_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1722_ _0319_ tt_um_rejunity_ay8913.tone_C_generator.period\[0\] tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
+ _0330_ _0350_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_13_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ tt_um_rejunity_ay8913.noise_generator.period\[0\] _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2205_ _0155_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2067_ _0017_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2136_ _0086_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1705_ tt_um_rejunity_ay8913.tone_C_generator.counter\[7\] _0332_ _0333_ tt_um_rejunity_ay8913.tone_C_generator.counter\[8\]
+ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1567_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\] _1023_ _0225_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1636_ _0276_ _0277_ _0270_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1498_ _0972_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2119_ _0069_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_1_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1280__A1 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1271__A1 _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1421_ _0892_ _0898_ _0900_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1352_ _0853_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_50_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1283_ _0806_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_46_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_22_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_22_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1619_ tt_um_rejunity_ay8913.noise_generator.lfsr\[11\] _0256_ _0265_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ _0553_ _0554_ tt_um_rejunity_ay8913.clk_counter\[2\] _0556_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1404_ tt_um_rejunity_ay8913.envelope_generator.period\[14\] _0887_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1335_ _0667_ _0763_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput2 custom_settings[1] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1266_ _0795_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1197_ _0743_ _0747_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1051_ tt_um_rejunity_ay8913.latched_register\[1\] _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1120_ tt_um_rejunity_ay8913.pwm_master.accumulator\[2\] net19 _0688_ _0013_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1953_ _0493_ _0545_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1884_ _0448_ _0488_ _0473_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1318_ tt_um_rejunity_ay8913.pwm_B.accumulator\[7\] _0827_ _0829_ _0830_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1249_ _0667_ _0782_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1686__A1 _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2152_ _0102_ clknet_leaf_6_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2221_ _0171_ clknet_leaf_21_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1103_ _0674_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1034_ tt_um_rejunity_ay8913.noise_generator.lfsr\[0\] _0616_ _0608_ tt_um_rejunity_ay8913.envelope_A
+ _0617_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_2083_ _0033_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1936_ tt_um_rejunity_ay8913.tone_A_generator.counter\[3\] _0532_ _0510_ _0535_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1867_ _0417_ _0477_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1798_ tt_um_rejunity_ay8913.tone_B_generator.counter\[7\] _0414_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1112__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1721_ _0339_ tt_um_rejunity_ay8913.tone_C_generator.period\[2\] _0350_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1583_ _0674_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1652_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\] _0290_ _0291_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2135_ _0085_ clknet_leaf_29_wb_clk_i net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2204_ _0154_ clknet_leaf_32_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2066_ _0016_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1919_ _0520_ tt_um_rejunity_ay8913.tone_A_generator.period\[11\] _0522_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1704_ tt_um_rejunity_ay8913.tone_C_generator.period\[8\] _0333_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1566_ _0989_ _0224_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1497_ _0926_ _0964_ _0971_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1635_ tt_um_rejunity_ay8913.noise_generator.lfsr\[14\] _0272_ _0277_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2049_ _0840_ _0606_ _0607_ _0611_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2118_ _0068_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_1_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1351_ _0776_ _0850_ _0851_ tt_um_rejunity_ay8913.tone_A_generator.period\[5\] _0853_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1420_ _0899_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1282_ _0778_ _0802_ _0803_ tt_um_rejunity_ay8913.tone_B_generator.period\[6\] _0806_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_46_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1618_ _0263_ _0264_ _0259_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1549_ _0942_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_49_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_39_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1403_ _0884_ _0885_ _0881_ _0886_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1265_ _0790_ _0792_ _0794_ tt_um_rejunity_ay8913.tone_B_generator.period\[0\] _0795_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1334_ _0840_ _0837_ _0838_ _0841_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1196_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\] _0724_ _0735_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\]
+ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput3 io_in_1[0] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1050_ tt_um_rejunity_ay8913.latched_register\[3\] _0631_ _0632_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1952_ _0525_ _0544_ _0545_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_43_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1883_ tt_um_rejunity_ay8913.tone_B_generator.counter\[10\] _0486_ _0488_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1248_ _0633_ _0654_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1317_ _0680_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_54_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1179_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\] _0727_ _0736_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\]
+ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2151_ _0101_ clknet_leaf_7_wb_clk_i tt_um_rejunity_ay8913.restart_envelope vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2220_ _0170_ clknet_leaf_21_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1102_ _0640_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2082_ _0032_ clknet_leaf_2_wb_clk_i tt_um_rejunity_ay8913.pwm_C.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1033_ tt_um_rejunity_ay8913.amplitude_A\[0\] tt_um_rejunity_ay8913.envelope_A tt_um_rejunity_ay8913.tone_disable_A
+ tt_um_rejunity_ay8913.tone_A _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1935_ _0533_ _0534_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1639__B _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1866_ _0418_ _0435_ _0471_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_26_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1797_ _0412_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1374__A1 _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1117__A1 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1720_ tt_um_rejunity_ay8913.tone_C_generator.counter\[6\] _0347_ _0348_ tt_um_rejunity_ay8913.tone_C_generator.counter\[5\]
+ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1651_ tt_um_rejunity_ay8913.noise_generator.period\[1\] _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1582_ _0619_ _0237_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2134_ _0084_ clknet_leaf_35_wb_clk_i net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2065_ _0015_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2203_ _0153_ clknet_leaf_24_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input6_I io_in_1[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_16_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_16_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_44_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1918_ _0520_ tt_um_rejunity_ay8913.tone_A_generator.period\[11\] tt_um_rejunity_ay8913.tone_A_generator.period\[10\]
+ _0493_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1849_ _0464_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1889__A2 _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1634_ tt_um_rejunity_ay8913.noise_generator.lfsr\[15\] _0267_ _0276_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1329__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1703_ tt_um_rejunity_ay8913.tone_C_generator.period\[7\] _0332_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1565_ _0948_ _1023_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1496_ _0928_ _0967_ _0955_ _0970_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_39_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1501__A1 _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2117_ _0067_ clknet_leaf_38_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2048_ _0665_ _0606_ _0607_ _0610_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_44_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1740__A1 _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1350_ _0852_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1281_ _0805_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_46_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1617_ tt_um_rejunity_ay8913.noise_generator.lfsr\[9\] _0261_ _0264_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1548_ _1006_ _1011_ _1012_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1479_ _0949_ _0950_ _0952_ _0953_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xclkbuf_leaf_31_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_31_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1789__A1 _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1402_ net8 _0876_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1264_ _0793_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1333_ tt_um_rejunity_ay8913.envelope_A _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput4 io_in_1[1] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1195_ _0743_ _0746_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1951_ tt_um_rejunity_ay8913.tone_A_generator.counter\[9\] _0543_ _0545_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1882_ _0467_ _0487_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_47_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1178_ _0735_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1316_ _0827_ _0828_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1247_ _0781_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2150_ _0100_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[15\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1101_ _0666_ _0669_ _0673_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1032_ tt_um_rejunity_ay8913.noise_disable_A _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2081_ _0031_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1934_ _0505_ _0532_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1865_ _0473_ _0476_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1796_ _0410_ tt_um_rejunity_ay8913.tone_B_generator.period\[9\] tt_um_rejunity_ay8913.tone_B_generator.period\[8\]
+ _0411_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1581_ _0236_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1650_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\] _0289_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_13_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2202_ _0152_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.envelope_continue vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2133_ _0083_ clknet_leaf_30_wb_clk_i net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2064_ _0014_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1917_ tt_um_rejunity_ay8913.tone_A_generator.counter\[11\] _0520_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1848_ _0373_ _0463_ _0670_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1779_ _0399_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1274__A1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1564_ _1006_ _1022_ _1023_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_41_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1633_ _0274_ _0275_ _0270_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1702_ _0319_ tt_um_rejunity_ay8913.tone_C_generator.period\[0\] tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
+ _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1495_ _0915_ _0968_ _0956_ _0969_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1501__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1265__A1 _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2116_ _0066_ clknet_leaf_39_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2047_ _0811_ _0606_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1256__A1 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_1_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_1_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_23_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1280_ _0776_ _0802_ _0803_ tt_um_rejunity_ay8913.tone_B_generator.period\[5\] _0805_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1547_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\] _1004_ _0944_ _1012_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1616_ tt_um_rejunity_ay8913.noise_generator.lfsr\[10\] _0256_ _0263_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1478_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\] _0889_ _0943_
+ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\] _0953_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_37_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1789__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1401_ tt_um_rejunity_ay8913.envelope_generator.period\[13\] _0885_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1332_ _0650_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_36_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1263_ _0766_ _0791_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1194_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\] _0740_ _0741_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\]
+ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput5 io_in_1[2] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1950_ tt_um_rejunity_ay8913.tone_A_generator.counter\[9\] _0543_ _0544_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1881_ _0449_ _0486_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1315_ tt_um_rejunity_ay8913.pwm_B.accumulator\[6\] _0824_ _0822_ _0828_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1177_ _0730_ _0722_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1246_ _0780_ _0773_ _0774_ tt_um_rejunity_ay8913.tone_C_generator.period\[7\] _0781_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_output20_I net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1052__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1100_ _0671_ tt_um_rejunity_ay8913.tone_A_generator.period\[8\] _0672_ _0673_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2080_ _0030_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1031_ _0609_ _0614_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1933_ _0524_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2020__A1 _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1864_ _0418_ _0475_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1795_ tt_um_rejunity_ay8913.tone_B_generator.counter\[8\] _0411_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1229_ _0644_ _0765_ _0768_ tt_um_rejunity_ay8913.tone_C_generator.period\[1\] _0770_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2002__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1580_ _0235_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_13_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2132_ _0082_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2201_ _0151_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.envelope_attack vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1047__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2063_ _0013_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.pwm_master.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1916_ _0493_ tt_um_rejunity_ay8913.tone_A_generator.period\[10\] _0495_ _0517_ _0518_
+ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1847_ _0456_ _0457_ _0462_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1778_ _0391_ _0386_ _0397_ _0398_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_12_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_25_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_25_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1420__I _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_3__f_wb_clk_i clknet_0_wb_clk_i clknet_2_3__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1701_ tt_um_rejunity_ay8913.tone_C_generator.counter\[1\] _0330_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_14_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1563_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\] tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\]
+ _1020_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1494_ _0925_ _0924_ tt_um_rejunity_ay8913.envelope_generator.period\[0\] _0929_
+ _0935_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_39_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1632_ tt_um_rejunity_ay8913.noise_generator.lfsr\[13\] _0272_ _0275_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2115_ _0065_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.pwm_B.accumulator\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1505__I _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2046_ _0636_ _0836_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1546_ _1009_ _1010_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1477_ _0951_ tt_um_rejunity_ay8913.envelope_generator.period\[13\] tt_um_rejunity_ay8913.envelope_generator.period\[12\]
+ _0938_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1615_ _0260_ _0262_ _0259_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1235__I _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2029_ tt_um_rejunity_ay8913.pwm_A.accumulator\[4\] _0592_ _0595_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1331_ _0666_ _0837_ _0838_ _0839_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1165__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1400_ _0659_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1262_ _0791_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1193_ _0743_ _0745_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput6 io_in_1[3] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1529_ _0996_ _0997_ _0998_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1156__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ _0465_ _0485_ _0486_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1386__A1 _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1314_ _0826_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_54_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1245_ net10 _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1176_ _0733_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1368__A1 _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1030_ _0610_ _0611_ _0612_ tt_um_rejunity_ay8913.noise_generator.lfsr\[0\] _0613_
+ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1932_ _0527_ _0530_ _0532_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1863_ _0435_ _0471_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1794_ tt_um_rejunity_ay8913.tone_B_generator.counter\[9\] _0410_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1359__A1 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1228_ _0769_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_2_2__f_wb_clk_i clknet_0_wb_clk_i clknet_2_2__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1159_ _0719_ tt_um_rejunity_ay8913.pwm_master.accumulator\[8\] tt_um_rejunity_ay8913.pwm_master.accumulator\[9\]
+ _0711_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1522__A1 _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1153__I _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1053__A3 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1038__B1 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2131_ _0081_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2062_ _0012_ clknet_leaf_12_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2200_ _0150_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.envelope_alternate vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1063__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_14_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1915_ tt_um_rejunity_ay8913.tone_A_generator.counter\[9\] _0676_ _0518_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1846_ _0455_ _0430_ _0460_ _0461_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1777_ tt_um_rejunity_ay8913.tone_C_generator.counter\[8\] _0354_ _0392_ _0398_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_8_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input12_I io_in_2[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1631_ tt_um_rejunity_ay8913.noise_generator.lfsr\[14\] _0267_ _0274_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1700_ _0324_ _0328_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1562_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\] _1020_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\]
+ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1493_ _0913_ _0917_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2114_ _0064_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input4_I io_in_1[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2045_ _0605_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1829_ tt_um_rejunity_ay8913.tone_B_generator.counter\[8\] _0443_ _0444_ tt_um_rejunity_ay8913.tone_B_generator.counter\[7\]
+ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1964__A1 _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1614_ tt_um_rejunity_ay8913.noise_generator.lfsr\[8\] _0261_ _0262_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1545_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\] _1004_ _1010_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1476_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\] _0951_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_37_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2028_ _0592_ _0594_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1261_ _0636_ _0667_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1330_ tt_um_rejunity_ay8913.amplitude_A\[0\] _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 io_in_1[4] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1192_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\] _0740_ _0741_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\]
+ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_54_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1528_ _0922_ _0995_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1459_ _0926_ _0931_ _0933_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_40_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1083__A1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1066__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_1__f_wb_clk_i clknet_0_wb_clk_i clknet_2_1__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1313_ tt_um_rejunity_ay8913.pwm_B.accumulator\[6\] _0824_ _0826_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1244_ _0779_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_19_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_19_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1175_ _0732_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1074__A1 _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1301__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1931_ _0531_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput10 io_in_1[7] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1862_ _0473_ _0474_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1793_ _0408_ _0321_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1227_ _0630_ _0765_ _0768_ tt_um_rejunity_ay8913.tone_C_generator.period\[0\] _0769_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1158_ _0718_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1089_ _0663_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1053__A4 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2130_ _0080_ clknet_leaf_11_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2061_ _0011_ clknet_leaf_12_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1914_ tt_um_rejunity_ay8913.tone_A_generator.counter\[8\] _0494_ _0513_ _0515_ _0516_
+ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_44_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1845_ _0420_ _0436_ _0424_ _0445_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_4_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1776_ _0354_ _0392_ tt_um_rejunity_ay8913.tone_C_generator.counter\[8\] _0397_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2259_ _0209_ clknet_leaf_15_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1268__A1 _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_34_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_34_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_31_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1630_ _0271_ _0273_ _0270_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1561_ _1007_ _1021_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1492_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\] _0965_ _0966_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\]
+ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_49_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2113_ _0063_ clknet_leaf_30_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2044_ _0699_ tt_um_rejunity_ay8913.pwm_A.accumulator\[7\] tt_um_rejunity_ay8913.pwm_A.accumulator\[8\]
+ _0600_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_44_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1828_ tt_um_rejunity_ay8913.tone_B_generator.period\[7\] _0444_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1759_ _0370_ _0383_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_23_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1069__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1544_ _0944_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1613_ _0236_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1475_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\] _0887_ _0885_
+ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\] _0950_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_5_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2027_ tt_um_rejunity_ay8913.pwm_A.accumulator\[3\] _0590_ _0593_ _0594_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1260_ _0629_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput8 io_in_1[5] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1191_ _0743_ _0744_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_2_0__f_wb_clk_i clknet_0_wb_clk_i clknet_2_0__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_36_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1527_ _0922_ _0995_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1458_ _0919_ _0932_ _0923_ _0922_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1389_ _0677_ _0876_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_2_1__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1791__B _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1174_ _0658_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1312_ _0824_ _0825_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1082__I _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1243_ _0778_ _0773_ _0774_ tt_um_rejunity_ay8913.tone_C_generator.period\[6\] _0779_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2014__A1 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ tt_um_rejunity_ay8913.tone_A_generator.counter\[2\] _0499_ _0491_ _0979_ _0531_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
Xinput11 io_in_2[0] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1861_ _0422_ _0471_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1792_ tt_um_rejunity_ay8913.tone_B_generator.counter\[0\] _0408_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1157_ _0679_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1226_ _0767_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1088_ _0646_ _0657_ _0660_ tt_um_rejunity_ay8913.tone_C_generator.period\[10\] _0663_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1625__I _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_4_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_4_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_53_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2060_ _0010_ clknet_leaf_12_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1913_ _0514_ tt_um_rejunity_ay8913.tone_A_generator.period\[7\] _0516_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1844_ _0413_ _0458_ _0459_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1775_ _0396_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2258_ _0208_ clknet_leaf_15_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1270__I net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2189_ _0139_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1209_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1560_ _0938_ _1020_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1491_ tt_um_rejunity_ay8913.envelope_generator.period\[0\] _0966_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2112_ _0062_ clknet_leaf_31_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_49_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2043_ _0831_ _0604_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ tt_um_rejunity_ay8913.tone_B_generator.period\[8\] _0443_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1689_ _0318_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1758_ _0345_ _0381_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_23_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1175__I _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1101__A1 _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1543_ _1007_ _1008_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1474_ _0947_ tt_um_rejunity_ay8913.envelope_generator.period\[15\] tt_um_rejunity_ay8913.envelope_generator.period\[14\]
+ _0948_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_41_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1612_ tt_um_rejunity_ay8913.noise_generator.lfsr\[9\] _0256_ _0260_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2026_ _0680_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1331__A1 _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1398__A1 _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1119__B _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 io_in_1[6] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1190_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\] _0740_ _0741_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\]
+ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1389__A1 _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1526_ _0988_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1457_ tt_um_rejunity_ay8913.envelope_generator.period\[4\] _0932_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1388_ _0871_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2009_ _0582_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_ay8913_40 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1311_ tt_um_rejunity_ay8913.pwm_B.accumulator\[5\] _0821_ _0822_ _0825_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1242_ net9 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1173_ _0726_ _0727_ _0729_ _0731_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_28_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_28_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1509_ _0893_ _0902_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1273__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1525__A1 _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1860_ _0464_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput12 io_in_2[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1791_ _0406_ _0407_ _0857_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1358__I _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1516__A1 _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1156_ _0715_ _0717_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1087_ _0662_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1225_ _0766_ _0764_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1989_ tt_um_rejunity_ay8913.active _0569_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1994__A1 _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1912_ _0514_ tt_um_rejunity_ay8913.tone_A_generator.period\[7\] tt_um_rejunity_ay8913.tone_A_generator.period\[6\]
+ _0496_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1843_ _0416_ _0441_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1774_ _0370_ _0395_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2257_ _0207_ clknet_leaf_15_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1208_ tt_um_rejunity_ay8913.pwm_C.accumulator\[5\] _0752_ _0755_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2188_ _0138_ clknet_leaf_6_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1139_ _0681_ _0704_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1490_ tt_um_rejunity_ay8913.envelope_generator.period\[1\] _0965_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2111_ _0061_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2042_ tt_um_rejunity_ay8913.pwm_A.accumulator\[8\] _0603_ _0604_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_49_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ _0421_ _0438_ _0441_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1688_ _0800_ _0891_ _0314_ tt_um_rejunity_ay8913.envelope_continue _0318_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1990__B _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1757_ _0382_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input10_I io_in_1[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1611_ _0257_ _0258_ _0259_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1542_ _0912_ _1004_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1473_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\] _0948_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I custom_settings[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1315__B _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2025_ tt_um_rejunity_ay8913.pwm_A.accumulator\[3\] _0590_ _0592_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_49_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1809_ tt_um_rejunity_ay8913.tone_B_generator.counter\[1\] _0425_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1525_ _0989_ _0994_ _0995_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1456_ _0925_ _0924_ _0928_ _0930_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1387_ tt_um_rejunity_ay8913.envelope_generator.period\[9\] _0875_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2008_ _0683_ _0577_ _0579_ tt_um_rejunity_ay8913.envelope_generator.period\[2\]
+ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_ay8913_41 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_30 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_51_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1240__A1 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1310_ tt_um_rejunity_ay8913.pwm_B.accumulator\[5\] _0821_ _0824_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1241_ _0777_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1172_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\] _0730_ _0722_ _0718_ _0731_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1059__A1 _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1231__A1 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1439_ _0913_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1508_ _0900_ _0982_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 rst_n net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1790_ tt_um_rejunity_ay8913.tone_C _0991_ _0385_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1516__A2 _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2273_ _0223_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.envelope_C vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1224_ _0639_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1155_ tt_um_rejunity_ay8913.pwm_master.accumulator\[9\] _0716_ _0717_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1086_ _0644_ _0657_ _0660_ tt_um_rejunity_ay8913.tone_C_generator.period\[9\] _0662_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1988_ net12 net11 _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1682__A1 _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1911_ tt_um_rejunity_ay8913.tone_A_generator.counter\[7\] _0514_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1842_ _0408_ _0428_ _0431_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1773_ _0354_ _0392_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1318__B _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2256_ _0206_ clknet_leaf_14_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2187_ _0137_ clknet_leaf_6_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1207_ _0752_ _0754_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1138_ _0703_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1069_ net6 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_12_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_12_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_26_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1664__A1 _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1189__I _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2110_ _0060_ clknet_leaf_30_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2041_ tt_um_rejunity_ay8913.pwm_A.accumulator\[7\] _0599_ _0603_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1825_ tt_um_rejunity_ay8913.tone_B_generator.counter\[6\] _0439_ _0440_ tt_um_rejunity_ay8913.tone_B_generator.counter\[5\]
+ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1756_ _0371_ _0380_ _0381_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1687_ _0317_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2239_ _0189_ clknet_leaf_9_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1610_ _0733_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1541_ _1006_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1472_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\] _0947_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2024_ _0590_ _0591_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_20_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1808_ _0422_ tt_um_rejunity_ay8913.tone_B_generator.period\[3\] tt_um_rejunity_ay8913.tone_B_generator.period\[2\]
+ _0423_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1739_ _0329_ _0343_ _0357_ _0366_ _0367_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_31_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1524_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\] _0993_ _0995_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1455_ _0927_ tt_um_rejunity_ay8913.envelope_generator.period\[1\] tt_um_rejunity_ay8913.envelope_generator.period\[0\]
+ _0929_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1386_ _0666_ _0872_ _0874_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2007_ _0581_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1996__B _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_ay8913_31 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_38_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1171_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\] _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1240_ _0776_ _0773_ _0774_ tt_um_rejunity_ay8913.tone_C_generator.period\[5\] _0777_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_22_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1507_ _0963_ _0973_ _0981_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_2_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1438_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\] _0913_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1369_ _0863_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_37_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_37_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1745__I _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1154_ tt_um_rejunity_ay8913.pwm_master.accumulator\[8\] _0710_ _0716_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1223_ _0764_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2272_ _0222_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.amplitude_C\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1085_ _0661_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1987_ _0567_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1691__A2 _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1910_ _0496_ tt_um_rejunity_ay8913.tone_A_generator.period\[6\] _0508_ _0511_ _0512_
+ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1772_ _0394_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1841_ _0450_ _0451_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1370__A1 _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2255_ _0205_ clknet_leaf_15_wb_clk_i tt_um_rejunity_ay8913.latched_register\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2186_ _0136_ clknet_leaf_6_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_25_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1137_ _0695_ _0694_ tt_um_rejunity_ay8913.pwm_master.accumulator\[4\] tt_um_rejunity_ay8913.pwm_master.accumulator\[5\]
+ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_18_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1206_ tt_um_rejunity_ay8913.pwm_C.accumulator\[4\] _0750_ _0753_ _0754_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1068_ _0647_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2040_ tt_um_rejunity_ay8913.pwm_A.accumulator\[7\] _0600_ _0602_ _0219_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1686_ _0798_ _0101_ _0314_ tt_um_rejunity_ay8913.envelope_attack _0317_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1824_ tt_um_rejunity_ay8913.tone_B_generator.period\[5\] _0440_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1755_ _0378_ _0379_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2238_ _0188_ clknet_leaf_8_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1343__A1 _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2169_ _0119_ clknet_leaf_18_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1334__A1 _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1540_ _0988_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1471_ _0942_ _0875_ _0943_ _0944_ _0945_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_2023_ tt_um_rejunity_ay8913.pwm_A.accumulator\[2\] _0625_ _0559_ _0591_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1807_ tt_um_rejunity_ay8913.tone_B_generator.counter\[2\] _0423_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1738_ _0324_ _0327_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1669_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\] tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\]
+ _0981_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1523_ _0925_ _0993_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1454_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\] _0929_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1385_ _0671_ tt_um_rejunity_ay8913.envelope_generator.period\[8\] _0873_ _0874_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2006_ _0677_ _0577_ _0579_ tt_um_rejunity_ay8913.envelope_generator.period\[1\]
+ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_ay8913_32 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_7_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_7_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1170_ net20 _0728_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1437_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\] _0912_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1506_ _0980_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1368_ _0640_ _0861_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1299_ _0810_ _0816_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1921__A1 _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2271_ _0221_ clknet_leaf_36_wb_clk_i net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1153_ _0674_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1222_ _0632_ _0763_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1084_ _0630_ _0657_ _0660_ tt_um_rejunity_ay8913.tone_C_generator.period\[8\] _0661_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1988__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1986_ net12 net11 _0566_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1840_ _0413_ _0447_ _0455_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1771_ _0391_ _0386_ _0392_ _0393_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_8_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2254_ _0204_ clknet_leaf_14_wb_clk_i tt_um_rejunity_ay8913.latched_register\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2185_ _0135_ clknet_leaf_5_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1136_ tt_um_rejunity_ay8913.pwm_master.accumulator\[5\] _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1067_ _0646_ _0638_ _0642_ tt_um_rejunity_ay8913.noise_generator.period\[2\] _0647_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1205_ _0698_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1969_ _0553_ _0554_ _0555_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_21_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1823_ tt_um_rejunity_ay8913.tone_B_generator.period\[6\] _0439_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1685_ _0316_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1754_ _0378_ _0379_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2237_ _0187_ clknet_leaf_8_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2168_ _0118_ clknet_leaf_19_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1119_ tt_um_rejunity_ay8913.pwm_master.accumulator\[2\] net19 _0671_ _0688_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2099_ _0049_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1470_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\] _0878_ _0875_
+ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\] _0945_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_1_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2022_ tt_um_rejunity_ay8913.pwm_A.accumulator\[2\] _0625_ _0590_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1806_ tt_um_rejunity_ay8913.tone_B_generator.counter\[3\] _0422_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1737_ _0358_ _0365_ _0329_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1668_ _0305_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1599_ tt_um_rejunity_ay8913.noise_generator.lfsr\[4\] _0250_ _0251_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1243__A1 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1522_ _0989_ _0992_ _0993_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1453_ _0927_ tt_um_rejunity_ay8913.envelope_generator.period\[1\] _0928_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2005_ _0580_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1384_ _0871_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_ay8913_33 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1225__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1216__A1 _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1436_ _0903_ _0911_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1367_ _0861_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1505_ _0979_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1298_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\] _0814_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
+ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1221_ tt_um_rejunity_ay8913.latched_register\[1\] tt_um_rejunity_ay8913.latched_register\[0\]
+ _0635_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_9_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2270_ _0220_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1083_ _0659_ _0656_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1152_ tt_um_rejunity_ay8913.pwm_master.accumulator\[8\] _0711_ _0714_ _0019_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1988__A2 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1985_ net7 net10 net9 net8 _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_15_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1419_ _0658_ tt_um_rejunity_ay8913.restart_envelope _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1102__I _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1419__A1 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1770_ tt_um_rejunity_ay8913.tone_C_generator.counter\[6\] _0389_ _0393_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2184_ _0134_ clknet_leaf_5_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2253_ _0203_ clknet_leaf_14_wb_clk_i tt_um_rejunity_ay8913.latched_register\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1204_ tt_um_rejunity_ay8913.pwm_C.accumulator\[4\] _0750_ _0752_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_34_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1135_ _0697_ _0701_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1066_ net5 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1899_ tt_um_rejunity_ay8913.tone_A_generator.period\[0\] _0502_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1968_ _0553_ _0554_ _0829_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_2_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1822_ _0424_ _0432_ _0437_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1753_ tt_um_rejunity_ay8913.tone_C_generator.counter\[2\] tt_um_rejunity_ay8913.tone_C_generator.counter\[1\]
+ tt_um_rejunity_ay8913.tone_C_generator.counter\[0\] _0979_ _0379_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1684_ _0796_ _0101_ _0314_ tt_um_rejunity_ay8913.envelope_alternate _0316_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2236_ _0186_ clknet_leaf_9_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2167_ _0117_ clknet_leaf_17_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1118_ _0669_ _0685_ _0687_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1049_ tt_um_rejunity_ay8913.latched_register\[2\] _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2098_ _0048_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2047__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2021_ _0589_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1805_ _0420_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1736_ _0355_ _0364_ _0334_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1598_ _0236_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1667_ _0303_ _0304_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2219_ _0169_ clknet_leaf_22_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1452_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\] _0927_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1521_ _0927_ _0929_ _0976_ _0978_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1383_ _0871_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ _0629_ _0577_ _0579_ tt_um_rejunity_ay8913.envelope_generator.period\[0\]
+ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1719_ tt_um_rejunity_ay8913.tone_C_generator.period\[5\] _0348_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1105__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1170__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_ay8913_23 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_34 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1225__A2 _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1504_ _0976_ _0978_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_2_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1435_ tt_um_rejunity_ay8913.envelope_generator.stop _0894_ _0897_ _0910_ _0911_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1366_ _0632_ _0782_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1297_ _0810_ _0815_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1595__I _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_15_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_15_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1220_ _0762_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1151_ tt_um_rejunity_ay8913.pwm_master.accumulator\[8\] _0711_ _0707_ _0714_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1082_ _0658_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1984_ _0831_ _0565_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1349_ _0651_ _0850_ _0851_ tt_um_rejunity_ay8913.tone_A_generator.period\[4\] _0852_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1418_ _0897_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1364__A1 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1355__A1 _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2252_ _0202_ clknet_leaf_14_wb_clk_i tt_um_rejunity_ay8913.latched_register\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2183_ _0133_ clknet_leaf_5_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1134_ _0699_ _0700_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1203_ _0750_ _0751_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1065_ _0645_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1898_ _0499_ _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1967_ tt_um_rejunity_ay8913.clk_counter\[1\] _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1034__B1 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1337__A1 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_30_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_30_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_29_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ _0315_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1821_ _0436_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_29_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1752_ tt_um_rejunity_ay8913.tone_C_generator.counter\[3\] _0378_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1040__A3 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1576__A1 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2235_ _0185_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2166_ _0116_ clknet_leaf_18_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1117_ _0686_ _0672_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2097_ _0047_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1048_ _0629_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1108__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2020_ _0780_ _0584_ _0585_ tt_um_rejunity_ay8913.envelope_generator.period\[7\]
+ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_15_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1804_ _0417_ tt_um_rejunity_ay8913.tone_B_generator.period\[5\] tt_um_rejunity_ay8913.tone_B_generator.period\[4\]
+ _0419_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1735_ _0346_ _0362_ _0363_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1666_ tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\] _0986_ _0304_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1597_ tt_um_rejunity_ay8913.noise_generator.lfsr\[5\] _0245_ _0249_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2149_ _0099_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[14\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2218_ _0168_ clknet_leaf_22_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1788__A1 _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1960__A1 _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1520_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\] _0991_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\]
+ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1451_ _0922_ _0923_ _0924_ _0925_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1382_ tt_um_rejunity_ay8913.latched_register\[3\] tt_um_rejunity_ay8913.latched_register\[2\]
+ _0763_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2003_ _0578_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_33_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1649_ _0287_ _0288_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1718_ tt_um_rejunity_ay8913.tone_C_generator.period\[6\] _0347_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_16_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_ay8913_35 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_24 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1121__I _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1740__B _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1503_ _0974_ net1 _0977_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1434_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\] tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\]
+ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\] _0892_ _0910_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1296_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\] _0814_ _0815_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1365_ _0860_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1930__A4 _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1116__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1150_ _0711_ _0713_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1081_ _0639_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1070__A1 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1983_ tt_um_rejunity_ay8913.clk_counter\[6\] _0563_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1417_ _0894_ _0896_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1348_ _0844_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_43_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1279_ _0804_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2251_ _0201_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.active vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2182_ _0132_ clknet_leaf_5_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1133_ tt_um_rejunity_ay8913.pwm_master.accumulator\[4\] _0696_ _0700_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1064_ _0644_ _0638_ _0642_ tt_um_rejunity_ay8913.noise_generator.period\[1\] _0645_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1202_ tt_um_rejunity_ay8913.pwm_C.accumulator\[3\] _0748_ _0681_ _0751_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1966_ _0553_ _0239_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_0_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_0_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1897_ tt_um_rejunity_ay8913.tone_A_generator.period\[1\] _0500_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_3_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1282__A1 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1820_ tt_um_rejunity_ay8913.tone_B_generator.counter\[4\] _0433_ _0434_ _0435_ _0436_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_17_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1682_ _0790_ _0101_ _0314_ tt_um_rejunity_ay8913.envelope_generator.hold _0315_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1751_ _0377_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2234_ _0184_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2165_ _0115_ clknet_leaf_18_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1116_ net6 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2096_ _0046_ clknet_leaf_25_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1047_ net3 _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1949_ _0525_ _0542_ _0543_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_0_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1803_ _0418_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1246__A1 _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1734_ _0349_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1665_ _0718_ _0301_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1596_ _0246_ _0247_ _0248_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2217_ _0167_ clknet_leaf_22_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2148_ _0098_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[13\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2079_ _0029_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1788__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1237__A1 _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1450_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\] _0925_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1381_ _0870_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1920__C _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2002_ _0766_ _0576_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_33_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1648__B _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1648_ tt_um_rejunity_ay8913.noise_generator.lfsr\[16\] _0233_ _0822_ _0288_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1717_ _0344_ tt_um_rejunity_ay8913.tone_C_generator.period\[5\] tt_um_rejunity_ay8913.tone_C_generator.period\[4\]
+ _0345_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1579_ tt_um_rejunity_ay8913.noise_generator.signal_edge.signal _0231_ _0235_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xwrapped_ay8913_36 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_25 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_8_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1433_ _0903_ _0909_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1502_ tt_um_rejunity_ay8913.clk_counter\[3\] tt_um_rejunity_ay8913.clk_counter\[5\]
+ tt_um_rejunity_ay8913.clk_counter\[4\] tt_um_rejunity_ay8913.clk_counter\[6\] _0977_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__1688__A1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1295_ _0809_ _0813_ _0814_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1364_ tt_um_rejunity_ay8913.noise_generator.signal_edge.signal _0719_ _0860_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_18_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_24_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_24_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1080_ _0656_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1982_ _0563_ _0564_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1347_ _0842_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1416_ _0895_ tt_um_rejunity_ay8913.envelope_generator.hold tt_um_rejunity_ay8913.envelope_generator.stop
+ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1278_ _0651_ _0802_ _0803_ tt_um_rejunity_ay8913.tone_B_generator.period\[4\] _0804_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1555__C _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2010__A1 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2250_ _0200_ clknet_leaf_1_wb_clk_i tt_um_rejunity_ay8913.clk_counter\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1201_ tt_um_rejunity_ay8913.pwm_C.accumulator\[3\] _0748_ _0750_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_34_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2181_ _0131_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1063_ net4 _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1132_ _0698_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1965_ tt_um_rejunity_ay8913.clk_counter\[0\] _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1043__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1896_ tt_um_rejunity_ay8913.tone_A_generator.counter\[1\] _0499_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1025__A2 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1320__I _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1750_ _0370_ _0376_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _0732_ _0891_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2233_ _0183_ clknet_leaf_11_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2164_ _0114_ clknet_leaf_17_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input9_I io_in_1[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1115_ _0681_ tt_um_rejunity_ay8913.tone_A_generator.period\[11\] _0685_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1046_ _0628_ net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2095_ _0045_ clknet_leaf_26_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1948_ tt_um_rejunity_ay8913.tone_A_generator.counter\[8\] _0540_ _0543_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1879_ tt_um_rejunity_ay8913.tone_B_generator.counter\[9\] _0483_ _0486_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_22_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1802_ tt_um_rejunity_ay8913.tone_B_generator.counter\[4\] _0418_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1733_ _0359_ _0361_ _0338_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1664_ _0857_ _0302_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1595_ _0733_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2147_ _0097_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[12\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2216_ _0166_ clknet_leaf_24_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.counter\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1029_ tt_um_rejunity_ay8913.tone_C tt_um_rejunity_ay8913.tone_disable_C _0613_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2078_ _0028_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1380_ _0776_ _0861_ _0863_ tt_um_rejunity_ay8913.noise_disable_C _0870_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2001_ _0576_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1716_ tt_um_rejunity_ay8913.tone_C_generator.counter\[4\] _0345_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1578_ tt_um_rejunity_ay8913.noise_generator.lfsr\[1\] _0233_ _0234_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1647_ _0236_ _0286_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_ay8913_37 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_26 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_8_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1385__A1 _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1432_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\] _0907_ _0909_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1501_ _0974_ net1 _0975_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1688__A2 _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1363_ _0723_ _0810_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_53_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1294_ _0730_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\] tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
+ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1376__A1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1981_ tt_um_rejunity_ay8913.clk_counter\[5\] _0561_ _0559_ _0564_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1415_ tt_um_rejunity_ay8913.envelope_continue _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1346_ _0849_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1277_ _0793_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_3__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1349__A1 _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1200_ _0689_ _0748_ _0749_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2180_ _0130_ clknet_leaf_0_wb_clk_i tt_um_rejunity_ay8913.noise_generator.lfsr\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1131_ _0679_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1062_ _0643_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1895_ tt_um_rejunity_ay8913.tone_A_generator.counter\[2\] _0498_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1964_ _0840_ _0549_ _0550_ _0552_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1579__A1 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1503__A1 _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1329_ _0811_ _0837_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1680_ _0298_ _0311_ _0303_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2163_ _0113_ clknet_leaf_17_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2232_ _0182_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1114_ _0669_ _0682_ _0684_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1045_ _0626_ _0627_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2094_ _0044_ clknet_leaf_24_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1947_ tt_um_rejunity_ay8913.tone_A_generator.counter\[8\] _0540_ _0542_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1972__A1 _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1878_ tt_um_rejunity_ay8913.tone_B_generator.counter\[9\] _0483_ _0485_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1801_ tt_um_rejunity_ay8913.tone_B_generator.counter\[5\] _0417_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1732_ _0331_ _0360_ _0350_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1663_ tt_um_rejunity_ay8913.noise_generator.signal_edge.signal _0301_ _0302_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1594_ tt_um_rejunity_ay8913.noise_generator.lfsr\[3\] _0237_ _0247_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2146_ _0096_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2077_ _0027_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2215_ _0165_ clknet_leaf_33_wb_clk_i tt_um_rejunity_ay8913.tone_C vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1028_ tt_um_rejunity_ay8913.noise_disable_C _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_18_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_18_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_50_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2000_ _0782_ _0836_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1646_ tt_um_rejunity_ay8913.noise_generator.lfsr\[3\] _0619_ _0285_ _0286_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1715_ tt_um_rejunity_ay8913.tone_C_generator.counter\[5\] _0344_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1577_ _0232_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2129_ _0079_ clknet_leaf_11_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_ay8913_38 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_27 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_8_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1500_ tt_um_rejunity_ay8913.clk_counter\[0\] tt_um_rejunity_ay8913.clk_counter\[1\]
+ tt_um_rejunity_ay8913.clk_counter\[2\] _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_2_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1431_ _0906_ _0908_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1293_ _0808_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\] tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
+ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1362_ _0858_ _0736_ _0859_ _0831_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_53_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1629_ tt_um_rejunity_ay8913.noise_generator.lfsr\[12\] _0272_ _0273_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1300__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1119__A2 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_33_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_33_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_15_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1980_ tt_um_rejunity_ay8913.clk_counter\[5\] _0561_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1414_ _0893_ tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
+ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1345_ _0800_ _0843_ _0845_ tt_um_rejunity_ay8913.tone_A_generator.period\[3\] _0849_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1276_ _0791_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1130_ tt_um_rejunity_ay8913.pwm_master.accumulator\[4\] _0696_ _0697_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1061_ _0630_ _0638_ _0642_ tt_um_rejunity_ay8913.noise_generator.period\[0\] _0643_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1894_ tt_um_rejunity_ay8913.tone_A_generator.period\[4\] _0497_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_43_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ tt_um_rejunity_ay8913.envelope_B _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1200__A1 _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1503__A2 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1328_ _0763_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1259_ _0789_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1742__A2 _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1258__A1 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2231_ _0181_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2162_ _0112_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1113_ _0683_ _0672_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2093_ _0043_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1044_ _0609_ _0614_ _0625_ _0622_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_0_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1946_ _0525_ _0540_ _0541_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_43_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1877_ _0465_ _0483_ _0484_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_39_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1800_ _0414_ tt_um_rejunity_ay8913.tone_B_generator.period\[7\] tt_um_rejunity_ay8913.tone_B_generator.period\[6\]
+ _0415_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1403__A1 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1731_ _0330_ tt_um_rejunity_ay8913.tone_C_generator.period\[1\] _0360_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1662_ _0297_ _0299_ _0300_ _0990_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1593_ tt_um_rejunity_ay8913.noise_generator.lfsr\[4\] _0245_ _0246_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2214_ _0164_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2145_ _0095_ clknet_leaf_17_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1027_ tt_um_rejunity_ay8913.envelope_C _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2076_ _0026_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1929_ tt_um_rejunity_ay8913.tone_A_generator.counter\[2\] _0528_ _0530_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_42_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1927__A2 _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1645_ _0280_ _0284_ tt_um_rejunity_ay8913.noise_generator.lfsr\[3\] _0619_ _0285_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1714_ _0331_ _0335_ _0342_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_13_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1576_ tt_um_rejunity_ay8913.noise_generator.signal_edge.signal _0231_ _0232_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2059_ _0009_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2128_ _0078_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xwrapped_ay8913_39 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_ay8913_28 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1430_ _0900_ _0907_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1361_ net16 _0735_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1292_ _0808_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\] _0812_ _0061_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_3_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_3_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1559_ _1006_ _1018_ _1020_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1628_ _0235_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_37_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_21_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1413_ tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal _0893_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1344_ _0848_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1275_ _0801_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1060_ _0641_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ _0666_ _0549_ _0550_ _0551_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_51_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ tt_um_rejunity_ay8913.tone_A_generator.counter\[6\] _0496_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_43_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1503__A3 _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1327_ _0835_ tt_um_rejunity_ay8913.latched_register\[2\] _0836_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1189_ _0733_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1258_ _0648_ _0784_ _0785_ tt_um_rejunity_ay8913.tone_B_generator.period\[11\] _0789_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2230_ _0180_ clknet_leaf_10_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.counter\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2161_ _0111_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1112_ net5 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2092_ _0042_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1043_ _0625_ _0623_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1945_ tt_um_rejunity_ay8913.tone_A_generator.counter\[6\] _0537_ tt_um_rejunity_ay8913.tone_A_generator.counter\[7\]
+ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_31_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1876_ tt_um_rejunity_ay8913.tone_B_generator.counter\[8\] _0481_ _0484_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1100__A1 _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1592_ _0244_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1730_ _0341_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1661_ _0298_ tt_um_rejunity_ay8913.noise_generator.period\[4\] _0300_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2144_ _0094_ clknet_leaf_17_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input7_I io_in_1[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2213_ _0163_ clknet_leaf_28_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2075_ _0025_ clknet_leaf_36_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1026_ tt_um_rejunity_ay8913.amplitude_C\[0\] _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1928_ _0527_ _0528_ _0529_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1859_ _0467_ _0471_ _0472_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_8_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_27_wb_clk_i clknet_2_2__leaf_wb_clk_i clknet_leaf_27_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_50_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1713_ _0338_ _0341_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1644_ tt_um_rejunity_ay8913.noise_generator.lfsr\[4\] tt_um_rejunity_ay8913.noise_generator.lfsr\[2\]
+ tt_um_rejunity_ay8913.noise_generator.lfsr\[1\] _0283_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_13_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1575_ tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0
+ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_21_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2127_ _0077_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xwrapped_ay8913_29 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2058_ _0008_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[11\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1854__A2 _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1360_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\] _0858_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1291_ _0808_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\] _0728_ _0811_ _0812_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_53_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1558_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\] _1003_ _1019_
+ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1489_ _0921_ _0933_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1627_ tt_um_rejunity_ay8913.noise_generator.lfsr\[13\] _0267_ _0271_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1412_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\] _0892_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1343_ _0798_ _0843_ _0845_ tt_um_rejunity_ay8913.tone_A_generator.period\[2\] _0848_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1274_ _0800_ _0792_ _0794_ tt_um_rejunity_ay8913.tone_B_generator.period\[3\] _0801_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ tt_um_rejunity_ay8913.tone_A_generator.counter\[9\] _0676_ _0494_ tt_um_rejunity_ay8913.tone_A_generator.counter\[8\]
+ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_43_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1961_ tt_um_rejunity_ay8913.amplitude_B\[0\] _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1984__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1326_ tt_um_rejunity_ay8913.latched_register\[3\] _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1188_ _0734_ _0742_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1257_ _0788_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_49_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2160_ _0110_ clknet_leaf_16_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1111_ _0681_ tt_um_rejunity_ay8913.tone_A_generator.period\[10\] _0682_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2091_ _0041_ clknet_leaf_31_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1042_ _0618_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1944_ tt_um_rejunity_ay8913.tone_A_generator.counter\[7\] tt_um_rejunity_ay8913.tone_A_generator.counter\[6\]
+ _0537_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_31_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1875_ tt_um_rejunity_ay8913.tone_B_generator.counter\[8\] _0481_ _0483_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_39_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1309_ _0821_ _0823_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1591_ _0232_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ _0289_ tt_um_rejunity_ay8913.noise_generator.period\[3\] tt_um_rejunity_ay8913.noise_generator.period\[4\]
+ _0298_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_21_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2143_ _0093_ clknet_leaf_22_wb_clk_i tt_um_rejunity_ay8913.envelope_generator.period\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2212_ _0162_ clknet_leaf_28_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1025_ tt_um_rejunity_ay8913.envelope_C _0608_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2074_ _0024_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1927_ _0491_ _0991_ _0499_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1858_ tt_um_rejunity_ay8913.tone_B_generator.counter\[2\] _0468_ _0472_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1789_ _0307_ _0385_ tt_um_rejunity_ay8913.tone_C _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1176__I _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1643_ _0281_ _0282_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1712_ _0339_ tt_um_rejunity_ay8913.tone_C_generator.period\[2\] tt_um_rejunity_ay8913.tone_C_generator.period\[3\]
+ _0340_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1574_ tt_um_rejunity_ay8913.envelope_attack _0903_ _0230_ _0124_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2126_ _0076_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[1\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2057_ _0007_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[10\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1067__A1 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1790__A2 _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1290_ _0679_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1626_ _0268_ _0269_ _0270_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1557_ _1015_ _1013_ _1009_ _0912_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1488_ _0937_ _0957_ _0962_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2109_ _0059_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_11_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_11_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_2_0__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1342_ _0847_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1411_ _0891_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1273_ net6 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1609_ tt_um_rejunity_ay8913.noise_generator.lfsr\[7\] _0250_ _0258_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1681__A1 _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1891_ tt_um_rejunity_ay8913.tone_A_generator.period\[8\] _0494_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_36_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1960_ _0811_ _0549_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1308__B _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1325_ _0834_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1256_ _0646_ _0784_ _0785_ tt_um_rejunity_ay8913.tone_B_generator.period\[10\] _0788_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1187_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\] _0740_ _0741_ tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\]
+ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1663__A1 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ _0040_ clknet_leaf_31_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1110_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1041_ _0624_ net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1943_ _0533_ _0539_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1406__A1 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1874_ _0465_ _0481_ _0482_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1239_ net8 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_39_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1308_ tt_um_rejunity_ay8913.pwm_B.accumulator\[4\] _0819_ _0822_ _0823_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1590_ _0242_ _0243_ _0239_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1024_ tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\] tt_um_rejunity_ay8913.envelope_generator.invert_output
+ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_TAPCELL_ROW_36_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2142_ _0092_ clknet_leaf_3_wb_clk_i tt_um_rejunity_ay8913.noise_disable_C vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2211_ _0161_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2073_ _0023_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1926_ _0499_ _0491_ _0321_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1857_ _0470_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1788_ _0307_ _0385_ _0405_ _0322_ _0391_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_12_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2043__A1 _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_wb_clk_i clknet_2_0__leaf_wb_clk_i clknet_leaf_36_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1642_ tt_um_rejunity_ay8913.noise_generator.lfsr\[16\] tt_um_rejunity_ay8913.noise_generator.lfsr\[15\]
+ tt_um_rejunity_ay8913.noise_generator.lfsr\[14\] tt_um_rejunity_ay8913.noise_generator.lfsr\[13\]
+ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1711_ tt_um_rejunity_ay8913.tone_C_generator.counter\[3\] _0340_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1573_ tt_um_rejunity_ay8913.envelope_generator.invert_output _0228_ _0229_ _0230_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2125_ _0075_ clknet_leaf_13_wb_clk_i tt_um_rejunity_ay8913.tone_A_generator.period\[0\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2056_ _0006_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[9\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1909_ tt_um_rejunity_ay8913.tone_A_generator.counter\[5\] _0509_ _0512_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1790__A3 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1097__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1556_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\] _1017_ _1018_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1625_ _0674_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1487_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\] _0889_ _0949_
+ _0961_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_52_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2108_ _0058_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[6\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2039_ tt_um_rejunity_ay8913.pwm_A.accumulator\[7\] _0600_ _0856_ _0602_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1410_ _0835_ _0631_ tt_um_rejunity_ay8913.latched_register\[1\] _0654_ _0891_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1341_ _0796_ _0843_ _0845_ tt_um_rejunity_ay8913.tone_A_generator.period\[1\] _0847_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1272_ _0799_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1539_ _0996_ _1004_ _1005_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1608_ tt_um_rejunity_ay8913.noise_generator.lfsr\[8\] _0256_ _0257_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1681__A2 _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1890_ tt_um_rejunity_ay8913.tone_A_generator.counter\[10\] _0493_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_36_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1186_ _0735_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1324_ _0719_ tt_um_rejunity_ay8913.pwm_B.accumulator\[7\] tt_um_rejunity_ay8913.pwm_B.accumulator\[8\]
+ _0827_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1255_ _0787_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1994__B _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1351__A1 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1040_ _0615_ _0618_ _0623_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1942_ _0496_ _0537_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_2_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1873_ tt_um_rejunity_ay8913.tone_B_generator.counter\[6\] _0479_ tt_um_rejunity_ay8913.tone_B_generator.counter\[7\]
+ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1169_ tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\] tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
+ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1307_ _0698_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1238_ _0775_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2210_ _0160_ clknet_leaf_27_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.counter\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_28_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2141_ _0091_ clknet_leaf_23_wb_clk_i tt_um_rejunity_ay8913.noise_disable_B vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2072_ _0022_ clknet_leaf_35_wb_clk_i tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1925_ _0524_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_44_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_6_wb_clk_i clknet_2_1__leaf_wb_clk_i clknet_leaf_6_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_8_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1856_ tt_um_rejunity_ay8913.tone_B_generator.counter\[2\] _0425_ tt_um_rejunity_ay8913.tone_B_generator.counter\[0\]
+ _0979_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1787_ tt_um_rejunity_ay8913.tone_C_generator.counter\[10\] _0352_ _0398_ _0405_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_12_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1572_ tt_um_rejunity_ay8913.envelope_generator.invert_output _0228_ _0900_ _0229_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1641_ tt_um_rejunity_ay8913.noise_generator.lfsr\[12\] tt_um_rejunity_ay8913.noise_generator.lfsr\[11\]
+ tt_um_rejunity_ay8913.noise_generator.lfsr\[10\] tt_um_rejunity_ay8913.noise_generator.lfsr\[9\]
+ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_13_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1710_ tt_um_rejunity_ay8913.tone_C_generator.counter\[2\] _0339_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2124_ _0074_ clknet_leaf_3_wb_clk_i tt_um_rejunity_ay8913.envelope_A vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input5_I io_in_1[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2055_ _0005_ clknet_leaf_29_wb_clk_i tt_um_rejunity_ay8913.tone_C_generator.period\[8\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1908_ tt_um_rejunity_ay8913.tone_A_generator.counter\[5\] _0509_ _0497_ _0510_ _0511_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_29_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1839_ _0454_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1507__B _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1766__A1 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1555_ _1015_ _1016_ _1017_ _0989_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_41_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1624_ tt_um_rejunity_ay8913.noise_generator.lfsr\[11\] _0261_ _0269_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1486_ _0950_ _0960_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2107_ _0057_ clknet_leaf_20_wb_clk_i tt_um_rejunity_ay8913.tone_B_generator.period\[5\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2038_ _0600_ _0601_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_15_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_9_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1340_ _0846_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_20_wb_clk_i clknet_2_3__leaf_wb_clk_i clknet_leaf_20_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1271_ _0798_ _0792_ _0794_ tt_um_rejunity_ay8913.tone_B_generator.period\[2\] _0799_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_2_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1538_ _0913_ _1002_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1469_ tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\] _0944_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1607_ _0244_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1323_ _0831_ _0833_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1185_ _0724_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1254_ _0644_ _0784_ _0785_ tt_um_rejunity_ay8913.tone_B_generator.period\[9\] _0787_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1941_ _0527_ _0537_ _0538_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1872_ tt_um_rejunity_ay8913.tone_B_generator.counter\[7\] tt_um_rejunity_ay8913.tone_B_generator.counter\[6\]
+ _0479_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_24_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1306_ tt_um_rejunity_ay8913.pwm_B.accumulator\[4\] _0819_ _0821_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1099_ _0668_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1168_ _0724_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1237_ _0651_ _0773_ _0774_ tt_um_rejunity_ay8913.tone_C_generator.period\[4\] _0775_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2140_ _0090_ clknet_leaf_4_wb_clk_i tt_um_rejunity_ay8913.noise_disable_A vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1088__A1 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2071_ _0021_ clknet_leaf_37_wb_clk_i net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1924_ _0526_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1855_ _0467_ _0468_ _0469_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1786_ _0404_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2269_ _0219_ clknet_leaf_34_wb_clk_i tt_um_rejunity_ay8913.pwm_A.accumulator\[7\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1251__A1 _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1571_ _0895_ _0226_ _0227_ _0910_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1640_ tt_um_rejunity_ay8913.noise_generator.lfsr\[8\] tt_um_rejunity_ay8913.noise_generator.lfsr\[7\]
+ tt_um_rejunity_ay8913.noise_generator.lfsr\[6\] tt_um_rejunity_ay8913.noise_generator.lfsr\[5\]
+ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_21_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1793__A2 _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2123_ _0073_ clknet_leaf_14_wb_clk_i tt_um_rejunity_ay8913.amplitude_A\[0\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2054_ _0004_ clknet_leaf_32_wb_clk_i tt_um_rejunity_ay8913.noise_generator.period\[4\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1907_ tt_um_rejunity_ay8913.tone_A_generator.counter\[4\] _0510_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1838_ _0410_ tt_um_rejunity_ay8913.tone_B_generator.period\[9\] _0450_ _0453_ _0454_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1233__A1 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1769_ tt_um_rejunity_ay8913.tone_C_generator.counter\[6\] _0389_ _0392_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_2_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1766__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1554_ _1015_ _1013_ _1009_ _1010_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_1485_ _0940_ _0959_ _0952_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1623_ tt_um_rejunity_ay8913.noise_generator.lfsr\[12\] _0267_ _0268_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

