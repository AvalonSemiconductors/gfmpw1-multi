magic
tech gf180mcuD
magscale 1 5
timestamp 1712517913
<< obsm1 >>
rect 672 855 24808 24009
<< metal2 >>
rect 3136 25100 3192 25500
rect 9520 25100 9576 25500
rect 15904 25100 15960 25500
rect 22288 25100 22344 25500
rect 560 0 616 400
rect 1456 0 1512 400
rect 2352 0 2408 400
rect 3248 0 3304 400
rect 4144 0 4200 400
rect 5040 0 5096 400
rect 5936 0 5992 400
rect 6832 0 6888 400
rect 7728 0 7784 400
rect 8624 0 8680 400
rect 9520 0 9576 400
rect 10416 0 10472 400
rect 11312 0 11368 400
rect 12208 0 12264 400
rect 13104 0 13160 400
rect 14000 0 14056 400
rect 14896 0 14952 400
rect 15792 0 15848 400
rect 16688 0 16744 400
rect 17584 0 17640 400
rect 18480 0 18536 400
rect 19376 0 19432 400
rect 20272 0 20328 400
rect 21168 0 21224 400
rect 22064 0 22120 400
rect 22960 0 23016 400
rect 23856 0 23912 400
rect 24752 0 24808 400
<< obsm2 >>
rect 574 25070 3106 25100
rect 3222 25070 9490 25100
rect 9606 25070 15874 25100
rect 15990 25070 22258 25100
rect 22374 25070 24850 25100
rect 574 430 24850 25070
rect 646 350 1426 430
rect 1542 350 2322 430
rect 2438 350 3218 430
rect 3334 350 4114 430
rect 4230 350 5010 430
rect 5126 350 5906 430
rect 6022 350 6802 430
rect 6918 350 7698 430
rect 7814 350 8594 430
rect 8710 350 9490 430
rect 9606 350 10386 430
rect 10502 350 11282 430
rect 11398 350 12178 430
rect 12294 350 13074 430
rect 13190 350 13970 430
rect 14086 350 14866 430
rect 14982 350 15762 430
rect 15878 350 16658 430
rect 16774 350 17554 430
rect 17670 350 18450 430
rect 18566 350 19346 430
rect 19462 350 20242 430
rect 20358 350 21138 430
rect 21254 350 22034 430
rect 22150 350 22930 430
rect 23046 350 23826 430
rect 23942 350 24722 430
rect 24838 350 24850 430
<< metal3 >>
rect 25100 24416 25500 24472
rect 25100 22288 25500 22344
rect 25100 20160 25500 20216
rect 25100 18032 25500 18088
rect 25100 15904 25500 15960
rect 25100 13776 25500 13832
rect 25100 11648 25500 11704
rect 25100 9520 25500 9576
rect 25100 7392 25500 7448
rect 25100 5264 25500 5320
rect 25100 3136 25500 3192
rect 25100 1008 25500 1064
<< obsm3 >>
rect 849 24386 25070 24458
rect 849 22374 25100 24386
rect 849 22258 25070 22374
rect 849 20246 25100 22258
rect 849 20130 25070 20246
rect 849 18118 25100 20130
rect 849 18002 25070 18118
rect 849 15990 25100 18002
rect 849 15874 25070 15990
rect 849 13862 25100 15874
rect 849 13746 25070 13862
rect 849 11734 25100 13746
rect 849 11618 25070 11734
rect 849 9606 25100 11618
rect 849 9490 25070 9606
rect 849 7478 25100 9490
rect 849 7362 25070 7478
rect 849 5350 25100 7362
rect 849 5234 25070 5350
rect 849 3222 25100 5234
rect 849 3106 25070 3222
rect 849 1094 25100 3106
rect 849 1022 25070 1094
<< metal4 >>
rect 2224 1538 2384 23942
rect 9904 1538 10064 23942
rect 17584 1538 17744 23942
<< obsm4 >>
rect 1694 1689 2194 23511
rect 2414 1689 9874 23511
rect 10094 1689 17554 23511
rect 17774 1689 24122 23511
<< labels >>
rlabel metal3 s 25100 18032 25500 18088 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 25100 20160 25500 20216 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 25100 22288 25500 22344 6 custom_settings[2]
port 3 nsew signal input
rlabel metal3 s 25100 24416 25500 24472 6 custom_settings[3]
port 4 nsew signal input
rlabel metal3 s 25100 1008 25500 1064 6 io_in_1[0]
port 5 nsew signal input
rlabel metal3 s 25100 3136 25500 3192 6 io_in_1[1]
port 6 nsew signal input
rlabel metal3 s 25100 5264 25500 5320 6 io_in_1[2]
port 7 nsew signal input
rlabel metal3 s 25100 7392 25500 7448 6 io_in_1[3]
port 8 nsew signal input
rlabel metal3 s 25100 9520 25500 9576 6 io_in_1[4]
port 9 nsew signal input
rlabel metal3 s 25100 11648 25500 11704 6 io_in_1[5]
port 10 nsew signal input
rlabel metal3 s 25100 13776 25500 13832 6 io_in_1[6]
port 11 nsew signal input
rlabel metal3 s 25100 15904 25500 15960 6 io_in_1[7]
port 12 nsew signal input
rlabel metal2 s 15904 25100 15960 25500 6 io_in_2[0]
port 13 nsew signal input
rlabel metal2 s 22288 25100 22344 25500 6 io_in_2[1]
port 14 nsew signal input
rlabel metal2 s 560 0 616 400 6 io_out[0]
port 15 nsew signal output
rlabel metal2 s 9520 0 9576 400 6 io_out[10]
port 16 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 io_out[11]
port 17 nsew signal output
rlabel metal2 s 11312 0 11368 400 6 io_out[12]
port 18 nsew signal output
rlabel metal2 s 12208 0 12264 400 6 io_out[13]
port 19 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 io_out[14]
port 20 nsew signal output
rlabel metal2 s 14000 0 14056 400 6 io_out[15]
port 21 nsew signal output
rlabel metal2 s 14896 0 14952 400 6 io_out[16]
port 22 nsew signal output
rlabel metal2 s 15792 0 15848 400 6 io_out[17]
port 23 nsew signal output
rlabel metal2 s 16688 0 16744 400 6 io_out[18]
port 24 nsew signal output
rlabel metal2 s 17584 0 17640 400 6 io_out[19]
port 25 nsew signal output
rlabel metal2 s 1456 0 1512 400 6 io_out[1]
port 26 nsew signal output
rlabel metal2 s 18480 0 18536 400 6 io_out[20]
port 27 nsew signal output
rlabel metal2 s 19376 0 19432 400 6 io_out[21]
port 28 nsew signal output
rlabel metal2 s 20272 0 20328 400 6 io_out[22]
port 29 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 io_out[23]
port 30 nsew signal output
rlabel metal2 s 22064 0 22120 400 6 io_out[24]
port 31 nsew signal output
rlabel metal2 s 22960 0 23016 400 6 io_out[25]
port 32 nsew signal output
rlabel metal2 s 23856 0 23912 400 6 io_out[26]
port 33 nsew signal output
rlabel metal2 s 24752 0 24808 400 6 io_out[27]
port 34 nsew signal output
rlabel metal2 s 2352 0 2408 400 6 io_out[2]
port 35 nsew signal output
rlabel metal2 s 3248 0 3304 400 6 io_out[3]
port 36 nsew signal output
rlabel metal2 s 4144 0 4200 400 6 io_out[4]
port 37 nsew signal output
rlabel metal2 s 5040 0 5096 400 6 io_out[5]
port 38 nsew signal output
rlabel metal2 s 5936 0 5992 400 6 io_out[6]
port 39 nsew signal output
rlabel metal2 s 6832 0 6888 400 6 io_out[7]
port 40 nsew signal output
rlabel metal2 s 7728 0 7784 400 6 io_out[8]
port 41 nsew signal output
rlabel metal2 s 8624 0 8680 400 6 io_out[9]
port 42 nsew signal output
rlabel metal2 s 9520 25100 9576 25500 6 rst_n
port 43 nsew signal input
rlabel metal4 s 2224 1538 2384 23942 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 23942 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 23942 6 vss
port 45 nsew ground bidirectional
rlabel metal2 s 3136 25100 3192 25500 6 wb_clk_i
port 46 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 25500 25500
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2490036
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_ay8913/runs/24_04_07_21_21/results/signoff/wrapped_ay8913.magic.gds
string GDS_START 323206
<< end >>

