magic
tech gf180mcuD
magscale 1 10
timestamp 1702046264
<< metal1 >>
rect 1344 32170 34608 32204
rect 1344 32118 5372 32170
rect 5424 32118 5476 32170
rect 5528 32118 5580 32170
rect 5632 32118 13688 32170
rect 13740 32118 13792 32170
rect 13844 32118 13896 32170
rect 13948 32118 22004 32170
rect 22056 32118 22108 32170
rect 22160 32118 22212 32170
rect 22264 32118 30320 32170
rect 30372 32118 30424 32170
rect 30476 32118 30528 32170
rect 30580 32118 34608 32170
rect 1344 32084 34608 32118
rect 1344 31386 34768 31420
rect 1344 31334 9530 31386
rect 9582 31334 9634 31386
rect 9686 31334 9738 31386
rect 9790 31334 17846 31386
rect 17898 31334 17950 31386
rect 18002 31334 18054 31386
rect 18106 31334 26162 31386
rect 26214 31334 26266 31386
rect 26318 31334 26370 31386
rect 26422 31334 34478 31386
rect 34530 31334 34582 31386
rect 34634 31334 34686 31386
rect 34738 31334 34768 31386
rect 1344 31300 34768 31334
rect 1344 30602 34608 30636
rect 1344 30550 5372 30602
rect 5424 30550 5476 30602
rect 5528 30550 5580 30602
rect 5632 30550 13688 30602
rect 13740 30550 13792 30602
rect 13844 30550 13896 30602
rect 13948 30550 22004 30602
rect 22056 30550 22108 30602
rect 22160 30550 22212 30602
rect 22264 30550 30320 30602
rect 30372 30550 30424 30602
rect 30476 30550 30528 30602
rect 30580 30550 34608 30602
rect 1344 30516 34608 30550
rect 1344 29818 34768 29852
rect 1344 29766 9530 29818
rect 9582 29766 9634 29818
rect 9686 29766 9738 29818
rect 9790 29766 17846 29818
rect 17898 29766 17950 29818
rect 18002 29766 18054 29818
rect 18106 29766 26162 29818
rect 26214 29766 26266 29818
rect 26318 29766 26370 29818
rect 26422 29766 34478 29818
rect 34530 29766 34582 29818
rect 34634 29766 34686 29818
rect 34738 29766 34768 29818
rect 1344 29732 34768 29766
rect 1344 29034 34608 29068
rect 1344 28982 5372 29034
rect 5424 28982 5476 29034
rect 5528 28982 5580 29034
rect 5632 28982 13688 29034
rect 13740 28982 13792 29034
rect 13844 28982 13896 29034
rect 13948 28982 22004 29034
rect 22056 28982 22108 29034
rect 22160 28982 22212 29034
rect 22264 28982 30320 29034
rect 30372 28982 30424 29034
rect 30476 28982 30528 29034
rect 30580 28982 34608 29034
rect 1344 28948 34608 28982
rect 11218 28702 11230 28754
rect 11282 28702 11294 28754
rect 8418 28590 8430 28642
rect 8482 28590 8494 28642
rect 9090 28478 9102 28530
rect 9154 28478 9166 28530
rect 1344 28250 34768 28284
rect 1344 28198 9530 28250
rect 9582 28198 9634 28250
rect 9686 28198 9738 28250
rect 9790 28198 17846 28250
rect 17898 28198 17950 28250
rect 18002 28198 18054 28250
rect 18106 28198 26162 28250
rect 26214 28198 26266 28250
rect 26318 28198 26370 28250
rect 26422 28198 34478 28250
rect 34530 28198 34582 28250
rect 34634 28198 34686 28250
rect 34738 28198 34768 28250
rect 1344 28164 34768 28198
rect 20302 28082 20354 28094
rect 20302 28018 20354 28030
rect 5070 27970 5122 27982
rect 5070 27906 5122 27918
rect 4510 27858 4562 27870
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 4510 27794 4562 27806
rect 4846 27858 4898 27870
rect 4846 27794 4898 27806
rect 5182 27858 5234 27870
rect 19966 27858 20018 27870
rect 10210 27806 10222 27858
rect 10274 27806 10286 27858
rect 5182 27794 5234 27806
rect 19966 27794 20018 27806
rect 20190 27858 20242 27870
rect 20190 27794 20242 27806
rect 20526 27858 20578 27870
rect 20526 27794 20578 27806
rect 3614 27746 3666 27758
rect 10994 27694 11006 27746
rect 11058 27694 11070 27746
rect 13122 27694 13134 27746
rect 13186 27694 13198 27746
rect 3614 27682 3666 27694
rect 1344 27466 34608 27500
rect 1344 27414 5372 27466
rect 5424 27414 5476 27466
rect 5528 27414 5580 27466
rect 5632 27414 13688 27466
rect 13740 27414 13792 27466
rect 13844 27414 13896 27466
rect 13948 27414 22004 27466
rect 22056 27414 22108 27466
rect 22160 27414 22212 27466
rect 22264 27414 30320 27466
rect 30372 27414 30424 27466
rect 30476 27414 30528 27466
rect 30580 27414 34608 27466
rect 1344 27380 34608 27414
rect 5854 27298 5906 27310
rect 5854 27234 5906 27246
rect 4958 27186 5010 27198
rect 12238 27186 12290 27198
rect 4610 27134 4622 27186
rect 4674 27134 4686 27186
rect 10322 27134 10334 27186
rect 10386 27134 10398 27186
rect 17154 27134 17166 27186
rect 17218 27134 17230 27186
rect 20402 27134 20414 27186
rect 20466 27134 20478 27186
rect 4958 27122 5010 27134
rect 12238 27122 12290 27134
rect 5966 27074 6018 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 5966 27010 6018 27022
rect 6190 27074 6242 27086
rect 6190 27010 6242 27022
rect 6750 27074 6802 27086
rect 12462 27074 12514 27086
rect 23774 27074 23826 27086
rect 7410 27022 7422 27074
rect 7474 27022 7486 27074
rect 14354 27022 14366 27074
rect 14418 27022 14430 27074
rect 17602 27022 17614 27074
rect 17666 27022 17678 27074
rect 24210 27022 24222 27074
rect 24274 27022 24286 27074
rect 6750 27010 6802 27022
rect 12462 27010 12514 27022
rect 23774 27010 23826 27022
rect 5070 26962 5122 26974
rect 2482 26910 2494 26962
rect 2546 26910 2558 26962
rect 5070 26898 5122 26910
rect 6302 26962 6354 26974
rect 6302 26898 6354 26910
rect 6638 26962 6690 26974
rect 6638 26898 6690 26910
rect 6862 26962 6914 26974
rect 12126 26962 12178 26974
rect 8194 26910 8206 26962
rect 8258 26910 8270 26962
rect 6862 26898 6914 26910
rect 12126 26898 12178 26910
rect 12686 26962 12738 26974
rect 15026 26910 15038 26962
rect 15090 26910 15102 26962
rect 18274 26910 18286 26962
rect 18338 26910 18350 26962
rect 24098 26910 24110 26962
rect 24162 26910 24174 26962
rect 12686 26898 12738 26910
rect 23426 26798 23438 26850
rect 23490 26798 23502 26850
rect 1344 26682 34768 26716
rect 1344 26630 9530 26682
rect 9582 26630 9634 26682
rect 9686 26630 9738 26682
rect 9790 26630 17846 26682
rect 17898 26630 17950 26682
rect 18002 26630 18054 26682
rect 18106 26630 26162 26682
rect 26214 26630 26266 26682
rect 26318 26630 26370 26682
rect 26422 26630 34478 26682
rect 34530 26630 34582 26682
rect 34634 26630 34686 26682
rect 34738 26630 34768 26682
rect 1344 26596 34768 26630
rect 9886 26514 9938 26526
rect 9886 26450 9938 26462
rect 16270 26514 16322 26526
rect 16270 26450 16322 26462
rect 18062 26514 18114 26526
rect 18062 26450 18114 26462
rect 18958 26514 19010 26526
rect 18958 26450 19010 26462
rect 25678 26514 25730 26526
rect 25678 26450 25730 26462
rect 16606 26402 16658 26414
rect 7298 26350 7310 26402
rect 7362 26350 7374 26402
rect 16606 26338 16658 26350
rect 19182 26402 19234 26414
rect 25342 26402 25394 26414
rect 20402 26350 20414 26402
rect 20466 26350 20478 26402
rect 19182 26338 19234 26350
rect 25342 26338 25394 26350
rect 12350 26290 12402 26302
rect 16158 26290 16210 26302
rect 1810 26238 1822 26290
rect 1874 26238 1886 26290
rect 7970 26238 7982 26290
rect 8034 26238 8046 26290
rect 11778 26238 11790 26290
rect 11842 26238 11854 26290
rect 15810 26238 15822 26290
rect 15874 26238 15886 26290
rect 12350 26226 12402 26238
rect 16158 26226 16210 26238
rect 16382 26290 16434 26302
rect 16382 26226 16434 26238
rect 17838 26290 17890 26302
rect 17838 26226 17890 26238
rect 18174 26290 18226 26302
rect 18174 26226 18226 26238
rect 18286 26290 18338 26302
rect 18286 26226 18338 26238
rect 18734 26290 18786 26302
rect 18734 26226 18786 26238
rect 18846 26290 18898 26302
rect 25566 26290 25618 26302
rect 19618 26238 19630 26290
rect 19682 26238 19694 26290
rect 18846 26226 18898 26238
rect 25566 26226 25618 26238
rect 25790 26290 25842 26302
rect 25790 26226 25842 26238
rect 9998 26178 10050 26190
rect 2482 26126 2494 26178
rect 2546 26126 2558 26178
rect 4610 26126 4622 26178
rect 4674 26126 4686 26178
rect 5170 26126 5182 26178
rect 5234 26126 5246 26178
rect 9998 26114 10050 26126
rect 12462 26178 12514 26190
rect 12898 26126 12910 26178
rect 12962 26126 12974 26178
rect 15026 26126 15038 26178
rect 15090 26126 15102 26178
rect 22530 26126 22542 26178
rect 22594 26126 22606 26178
rect 12462 26114 12514 26126
rect 1344 25898 34608 25932
rect 1344 25846 5372 25898
rect 5424 25846 5476 25898
rect 5528 25846 5580 25898
rect 5632 25846 13688 25898
rect 13740 25846 13792 25898
rect 13844 25846 13896 25898
rect 13948 25846 22004 25898
rect 22056 25846 22108 25898
rect 22160 25846 22212 25898
rect 22264 25846 30320 25898
rect 30372 25846 30424 25898
rect 30476 25846 30528 25898
rect 30580 25846 34608 25898
rect 1344 25812 34608 25846
rect 2606 25730 2658 25742
rect 2606 25666 2658 25678
rect 2942 25730 2994 25742
rect 2942 25666 2994 25678
rect 3278 25730 3330 25742
rect 3278 25666 3330 25678
rect 18510 25730 18562 25742
rect 18510 25666 18562 25678
rect 18958 25730 19010 25742
rect 18958 25666 19010 25678
rect 19294 25730 19346 25742
rect 19294 25666 19346 25678
rect 13582 25618 13634 25630
rect 4946 25566 4958 25618
rect 5010 25566 5022 25618
rect 9874 25566 9886 25618
rect 9938 25566 9950 25618
rect 13582 25554 13634 25566
rect 14478 25618 14530 25630
rect 14478 25554 14530 25566
rect 15374 25618 15426 25630
rect 15374 25554 15426 25566
rect 19966 25618 20018 25630
rect 22978 25566 22990 25618
rect 23042 25566 23054 25618
rect 19966 25554 20018 25566
rect 12574 25506 12626 25518
rect 2594 25454 2606 25506
rect 2658 25454 2670 25506
rect 3266 25454 3278 25506
rect 3330 25454 3342 25506
rect 4610 25454 4622 25506
rect 4674 25454 4686 25506
rect 7074 25454 7086 25506
rect 7138 25454 7150 25506
rect 12002 25454 12014 25506
rect 12066 25454 12078 25506
rect 12574 25442 12626 25454
rect 13694 25506 13746 25518
rect 13694 25442 13746 25454
rect 14142 25506 14194 25518
rect 14142 25442 14194 25454
rect 14254 25506 14306 25518
rect 14254 25442 14306 25454
rect 14702 25506 14754 25518
rect 14702 25442 14754 25454
rect 15150 25506 15202 25518
rect 15150 25442 15202 25454
rect 15486 25506 15538 25518
rect 15486 25442 15538 25454
rect 15822 25506 15874 25518
rect 15822 25442 15874 25454
rect 18622 25506 18674 25518
rect 18622 25442 18674 25454
rect 20078 25506 20130 25518
rect 26350 25506 26402 25518
rect 25890 25454 25902 25506
rect 25954 25454 25966 25506
rect 20078 25442 20130 25454
rect 26350 25442 26402 25454
rect 3614 25394 3666 25406
rect 3614 25330 3666 25342
rect 4062 25394 4114 25406
rect 12350 25394 12402 25406
rect 7746 25342 7758 25394
rect 7810 25342 7822 25394
rect 4062 25330 4114 25342
rect 12350 25330 12402 25342
rect 14926 25394 14978 25406
rect 14926 25330 14978 25342
rect 16158 25394 16210 25406
rect 16158 25330 16210 25342
rect 16606 25394 16658 25406
rect 16606 25330 16658 25342
rect 19518 25394 19570 25406
rect 19518 25330 19570 25342
rect 19854 25394 19906 25406
rect 26574 25394 26626 25406
rect 25218 25342 25230 25394
rect 25282 25342 25294 25394
rect 19854 25330 19906 25342
rect 26574 25330 26626 25342
rect 26910 25394 26962 25406
rect 26910 25330 26962 25342
rect 27358 25394 27410 25406
rect 27358 25330 27410 25342
rect 27582 25394 27634 25406
rect 27582 25330 27634 25342
rect 12462 25282 12514 25294
rect 12462 25218 12514 25230
rect 13470 25282 13522 25294
rect 13470 25218 13522 25230
rect 16270 25282 16322 25294
rect 16270 25218 16322 25230
rect 16382 25282 16434 25294
rect 16382 25218 16434 25230
rect 20302 25282 20354 25294
rect 20302 25218 20354 25230
rect 26686 25282 26738 25294
rect 26686 25218 26738 25230
rect 27470 25282 27522 25294
rect 27470 25218 27522 25230
rect 28142 25282 28194 25294
rect 28142 25218 28194 25230
rect 1344 25114 34768 25148
rect 1344 25062 9530 25114
rect 9582 25062 9634 25114
rect 9686 25062 9738 25114
rect 9790 25062 17846 25114
rect 17898 25062 17950 25114
rect 18002 25062 18054 25114
rect 18106 25062 26162 25114
rect 26214 25062 26266 25114
rect 26318 25062 26370 25114
rect 26422 25062 34478 25114
rect 34530 25062 34582 25114
rect 34634 25062 34686 25114
rect 34738 25062 34768 25114
rect 1344 25028 34768 25062
rect 8878 24946 8930 24958
rect 4722 24894 4734 24946
rect 4786 24894 4798 24946
rect 6178 24894 6190 24946
rect 6242 24894 6254 24946
rect 8878 24882 8930 24894
rect 11006 24946 11058 24958
rect 11006 24882 11058 24894
rect 11118 24946 11170 24958
rect 11118 24882 11170 24894
rect 11230 24946 11282 24958
rect 11230 24882 11282 24894
rect 12462 24946 12514 24958
rect 12462 24882 12514 24894
rect 15150 24946 15202 24958
rect 15150 24882 15202 24894
rect 15262 24946 15314 24958
rect 24334 24946 24386 24958
rect 17490 24894 17502 24946
rect 17554 24894 17566 24946
rect 18162 24894 18174 24946
rect 18226 24894 18238 24946
rect 18834 24894 18846 24946
rect 18898 24894 18910 24946
rect 15262 24882 15314 24894
rect 24334 24882 24386 24894
rect 11342 24834 11394 24846
rect 4050 24782 4062 24834
rect 4114 24782 4126 24834
rect 5842 24782 5854 24834
rect 5906 24782 5918 24834
rect 6402 24782 6414 24834
rect 6466 24782 6478 24834
rect 11342 24770 11394 24782
rect 12350 24834 12402 24846
rect 12350 24770 12402 24782
rect 12686 24834 12738 24846
rect 12686 24770 12738 24782
rect 13470 24834 13522 24846
rect 13470 24770 13522 24782
rect 14254 24834 14306 24846
rect 14254 24770 14306 24782
rect 15710 24834 15762 24846
rect 24658 24782 24670 24834
rect 24722 24782 24734 24834
rect 28690 24782 28702 24834
rect 28754 24782 28766 24834
rect 15710 24770 15762 24782
rect 4398 24722 4450 24734
rect 4398 24658 4450 24670
rect 5070 24722 5122 24734
rect 5070 24658 5122 24670
rect 5294 24722 5346 24734
rect 12238 24722 12290 24734
rect 5618 24670 5630 24722
rect 5682 24670 5694 24722
rect 11666 24670 11678 24722
rect 11730 24670 11742 24722
rect 5294 24658 5346 24670
rect 12238 24658 12290 24670
rect 12574 24722 12626 24734
rect 14142 24722 14194 24734
rect 13122 24670 13134 24722
rect 13186 24670 13198 24722
rect 12574 24658 12626 24670
rect 14142 24658 14194 24670
rect 14478 24722 14530 24734
rect 14478 24658 14530 24670
rect 14590 24722 14642 24734
rect 14590 24658 14642 24670
rect 15038 24722 15090 24734
rect 15038 24658 15090 24670
rect 17838 24722 17890 24734
rect 22654 24722 22706 24734
rect 18386 24670 18398 24722
rect 18450 24670 18462 24722
rect 19058 24670 19070 24722
rect 19122 24670 19134 24722
rect 20290 24670 20302 24722
rect 20354 24670 20366 24722
rect 23426 24670 23438 24722
rect 23490 24670 23502 24722
rect 29362 24670 29374 24722
rect 29426 24670 29438 24722
rect 17838 24658 17890 24670
rect 22654 24658 22706 24670
rect 8990 24610 9042 24622
rect 8990 24546 9042 24558
rect 13358 24610 13410 24622
rect 20514 24558 20526 24610
rect 20578 24558 20590 24610
rect 22418 24558 22430 24610
rect 22482 24558 22494 24610
rect 26450 24558 26462 24610
rect 26514 24558 26526 24610
rect 13358 24546 13410 24558
rect 15598 24498 15650 24510
rect 15598 24434 15650 24446
rect 1344 24330 34608 24364
rect 1344 24278 5372 24330
rect 5424 24278 5476 24330
rect 5528 24278 5580 24330
rect 5632 24278 13688 24330
rect 13740 24278 13792 24330
rect 13844 24278 13896 24330
rect 13948 24278 22004 24330
rect 22056 24278 22108 24330
rect 22160 24278 22212 24330
rect 22264 24278 30320 24330
rect 30372 24278 30424 24330
rect 30476 24278 30528 24330
rect 30580 24278 34608 24330
rect 1344 24244 34608 24278
rect 12126 24162 12178 24174
rect 12126 24098 12178 24110
rect 13582 24162 13634 24174
rect 13582 24098 13634 24110
rect 18846 24162 18898 24174
rect 18846 24098 18898 24110
rect 11006 24050 11058 24062
rect 20302 24050 20354 24062
rect 28030 24050 28082 24062
rect 9986 23998 9998 24050
rect 10050 23998 10062 24050
rect 14914 23998 14926 24050
rect 14978 23998 14990 24050
rect 19170 23998 19182 24050
rect 19234 23998 19246 24050
rect 19842 23998 19854 24050
rect 19906 23998 19918 24050
rect 22418 23998 22430 24050
rect 22482 23998 22494 24050
rect 11006 23986 11058 23998
rect 20302 23986 20354 23998
rect 28030 23986 28082 23998
rect 10894 23938 10946 23950
rect 13022 23938 13074 23950
rect 7074 23886 7086 23938
rect 7138 23886 7150 23938
rect 11666 23886 11678 23938
rect 11730 23886 11742 23938
rect 10894 23874 10946 23886
rect 13022 23874 13074 23886
rect 13470 23938 13522 23950
rect 13470 23874 13522 23886
rect 14142 23938 14194 23950
rect 24222 23938 24274 23950
rect 27918 23938 27970 23950
rect 17826 23886 17838 23938
rect 17890 23886 17902 23938
rect 22194 23886 22206 23938
rect 22258 23886 22270 23938
rect 22754 23886 22766 23938
rect 22818 23886 22830 23938
rect 23426 23886 23438 23938
rect 23490 23886 23502 23938
rect 24546 23886 24558 23938
rect 24610 23886 24622 23938
rect 25554 23886 25566 23938
rect 25618 23886 25630 23938
rect 14142 23874 14194 23886
rect 24222 23874 24274 23886
rect 27918 23874 27970 23886
rect 28142 23938 28194 23950
rect 28142 23874 28194 23886
rect 5070 23826 5122 23838
rect 11118 23826 11170 23838
rect 7858 23774 7870 23826
rect 7922 23774 7934 23826
rect 5070 23762 5122 23774
rect 11118 23762 11170 23774
rect 11230 23826 11282 23838
rect 11230 23762 11282 23774
rect 12014 23826 12066 23838
rect 12014 23762 12066 23774
rect 13918 23826 13970 23838
rect 19518 23826 19570 23838
rect 17154 23774 17166 23826
rect 17218 23774 17230 23826
rect 13918 23762 13970 23774
rect 19518 23762 19570 23774
rect 19742 23826 19794 23838
rect 19742 23762 19794 23774
rect 27134 23826 27186 23838
rect 27134 23762 27186 23774
rect 29150 23826 29202 23838
rect 29150 23762 29202 23774
rect 29374 23826 29426 23838
rect 29374 23762 29426 23774
rect 4846 23714 4898 23726
rect 4846 23650 4898 23662
rect 4958 23714 5010 23726
rect 4958 23650 5010 23662
rect 12126 23714 12178 23726
rect 12126 23650 12178 23662
rect 13694 23714 13746 23726
rect 13694 23650 13746 23662
rect 18510 23714 18562 23726
rect 18510 23650 18562 23662
rect 19070 23714 19122 23726
rect 27022 23714 27074 23726
rect 24770 23662 24782 23714
rect 24834 23662 24846 23714
rect 26114 23662 26126 23714
rect 26178 23662 26190 23714
rect 19070 23650 19122 23662
rect 27022 23650 27074 23662
rect 27246 23714 27298 23726
rect 27246 23650 27298 23662
rect 27470 23714 27522 23726
rect 27470 23650 27522 23662
rect 28366 23714 28418 23726
rect 28366 23650 28418 23662
rect 29262 23714 29314 23726
rect 29262 23650 29314 23662
rect 29934 23714 29986 23726
rect 29934 23650 29986 23662
rect 1344 23546 34768 23580
rect 1344 23494 9530 23546
rect 9582 23494 9634 23546
rect 9686 23494 9738 23546
rect 9790 23494 17846 23546
rect 17898 23494 17950 23546
rect 18002 23494 18054 23546
rect 18106 23494 26162 23546
rect 26214 23494 26266 23546
rect 26318 23494 26370 23546
rect 26422 23494 34478 23546
rect 34530 23494 34582 23546
rect 34634 23494 34686 23546
rect 34738 23494 34768 23546
rect 1344 23460 34768 23494
rect 8318 23378 8370 23390
rect 5506 23326 5518 23378
rect 5570 23326 5582 23378
rect 8318 23314 8370 23326
rect 8766 23378 8818 23390
rect 8766 23314 8818 23326
rect 9998 23378 10050 23390
rect 9998 23314 10050 23326
rect 12910 23378 12962 23390
rect 12910 23314 12962 23326
rect 13694 23378 13746 23390
rect 15822 23378 15874 23390
rect 14130 23326 14142 23378
rect 14194 23326 14206 23378
rect 14802 23326 14814 23378
rect 14866 23326 14878 23378
rect 13694 23314 13746 23326
rect 15822 23314 15874 23326
rect 15934 23378 15986 23390
rect 15934 23314 15986 23326
rect 16046 23378 16098 23390
rect 16046 23314 16098 23326
rect 18846 23378 18898 23390
rect 23886 23378 23938 23390
rect 22978 23326 22990 23378
rect 23042 23326 23054 23378
rect 24658 23326 24670 23378
rect 24722 23326 24734 23378
rect 25778 23326 25790 23378
rect 25842 23326 25854 23378
rect 18846 23314 18898 23326
rect 23886 23314 23938 23326
rect 9886 23266 9938 23278
rect 9886 23202 9938 23214
rect 10222 23266 10274 23278
rect 10222 23202 10274 23214
rect 10894 23266 10946 23278
rect 10894 23202 10946 23214
rect 11790 23266 11842 23278
rect 11790 23202 11842 23214
rect 12686 23266 12738 23278
rect 12686 23202 12738 23214
rect 13806 23266 13858 23278
rect 13806 23202 13858 23214
rect 18286 23266 18338 23278
rect 18286 23202 18338 23214
rect 19070 23266 19122 23278
rect 20290 23214 20302 23266
rect 20354 23214 20366 23266
rect 23538 23214 23550 23266
rect 23602 23214 23614 23266
rect 29138 23214 29150 23266
rect 29202 23214 29214 23266
rect 19070 23202 19122 23214
rect 5182 23154 5234 23166
rect 6078 23154 6130 23166
rect 1810 23102 1822 23154
rect 1874 23102 1886 23154
rect 5842 23102 5854 23154
rect 5906 23102 5918 23154
rect 5182 23090 5234 23102
rect 6078 23090 6130 23102
rect 10334 23154 10386 23166
rect 11454 23154 11506 23166
rect 13470 23154 13522 23166
rect 10658 23102 10670 23154
rect 10722 23102 10734 23154
rect 12114 23102 12126 23154
rect 12178 23102 12190 23154
rect 12450 23102 12462 23154
rect 12514 23102 12526 23154
rect 10334 23090 10386 23102
rect 11454 23090 11506 23102
rect 13470 23090 13522 23102
rect 14478 23154 14530 23166
rect 15374 23154 15426 23166
rect 15026 23102 15038 23154
rect 15090 23102 15102 23154
rect 14478 23090 14530 23102
rect 15374 23090 15426 23102
rect 18622 23154 18674 23166
rect 18622 23090 18674 23102
rect 19182 23154 19234 23166
rect 25230 23154 25282 23166
rect 19506 23102 19518 23154
rect 19570 23102 19582 23154
rect 24434 23102 24446 23154
rect 24498 23102 24510 23154
rect 19182 23090 19234 23102
rect 25230 23090 25282 23102
rect 25454 23154 25506 23166
rect 30034 23102 30046 23154
rect 30098 23102 30110 23154
rect 25454 23090 25506 23102
rect 4958 23042 5010 23054
rect 2482 22990 2494 23042
rect 2546 22990 2558 23042
rect 4610 22990 4622 23042
rect 4674 22990 4686 23042
rect 4958 22978 5010 22990
rect 8430 23042 8482 23054
rect 8430 22978 8482 22990
rect 8878 23042 8930 23054
rect 11678 23042 11730 23054
rect 17950 23042 18002 23054
rect 10770 22990 10782 23042
rect 10834 22990 10846 23042
rect 12562 22990 12574 23042
rect 12626 22990 12638 23042
rect 26786 22990 26798 23042
rect 26850 22990 26862 23042
rect 8878 22978 8930 22990
rect 11678 22978 11730 22990
rect 17950 22978 18002 22990
rect 6302 22930 6354 22942
rect 6302 22866 6354 22878
rect 6414 22930 6466 22942
rect 6414 22866 6466 22878
rect 11342 22930 11394 22942
rect 11342 22866 11394 22878
rect 17390 22930 17442 22942
rect 17390 22866 17442 22878
rect 17726 22930 17778 22942
rect 17726 22866 17778 22878
rect 1344 22762 34608 22796
rect 1344 22710 5372 22762
rect 5424 22710 5476 22762
rect 5528 22710 5580 22762
rect 5632 22710 13688 22762
rect 13740 22710 13792 22762
rect 13844 22710 13896 22762
rect 13948 22710 22004 22762
rect 22056 22710 22108 22762
rect 22160 22710 22212 22762
rect 22264 22710 30320 22762
rect 30372 22710 30424 22762
rect 30476 22710 30528 22762
rect 30580 22710 34608 22762
rect 1344 22676 34608 22710
rect 5630 22594 5682 22606
rect 5630 22530 5682 22542
rect 5742 22594 5794 22606
rect 5742 22530 5794 22542
rect 20302 22594 20354 22606
rect 26462 22594 26514 22606
rect 26114 22542 26126 22594
rect 26178 22542 26190 22594
rect 20302 22530 20354 22542
rect 26462 22530 26514 22542
rect 26686 22482 26738 22494
rect 2706 22430 2718 22482
rect 2770 22430 2782 22482
rect 4834 22430 4846 22482
rect 4898 22430 4910 22482
rect 7858 22430 7870 22482
rect 7922 22430 7934 22482
rect 24434 22430 24446 22482
rect 24498 22430 24510 22482
rect 26686 22418 26738 22430
rect 27134 22482 27186 22494
rect 27134 22418 27186 22430
rect 5966 22370 6018 22382
rect 1922 22318 1934 22370
rect 1986 22318 1998 22370
rect 5966 22306 6018 22318
rect 6078 22370 6130 22382
rect 19294 22370 19346 22382
rect 20414 22370 20466 22382
rect 25566 22370 25618 22382
rect 12898 22318 12910 22370
rect 12962 22318 12974 22370
rect 17490 22318 17502 22370
rect 17554 22318 17566 22370
rect 20066 22318 20078 22370
rect 20130 22318 20142 22370
rect 21522 22318 21534 22370
rect 21586 22318 21598 22370
rect 6078 22306 6130 22318
rect 19294 22306 19346 22318
rect 20414 22306 20466 22318
rect 25566 22306 25618 22318
rect 26910 22370 26962 22382
rect 26910 22306 26962 22318
rect 27918 22370 27970 22382
rect 27918 22306 27970 22318
rect 20638 22258 20690 22270
rect 15586 22206 15598 22258
rect 15650 22206 15662 22258
rect 19618 22206 19630 22258
rect 19682 22206 19694 22258
rect 20638 22194 20690 22206
rect 20750 22258 20802 22270
rect 22194 22206 22206 22258
rect 22258 22206 22270 22258
rect 20750 22194 20802 22206
rect 25678 22146 25730 22158
rect 25678 22082 25730 22094
rect 25902 22146 25954 22158
rect 25902 22082 25954 22094
rect 27246 22146 27298 22158
rect 27246 22082 27298 22094
rect 27470 22146 27522 22158
rect 27470 22082 27522 22094
rect 27806 22146 27858 22158
rect 27806 22082 27858 22094
rect 1344 21978 34768 22012
rect 1344 21926 9530 21978
rect 9582 21926 9634 21978
rect 9686 21926 9738 21978
rect 9790 21926 17846 21978
rect 17898 21926 17950 21978
rect 18002 21926 18054 21978
rect 18106 21926 26162 21978
rect 26214 21926 26266 21978
rect 26318 21926 26370 21978
rect 26422 21926 34478 21978
rect 34530 21926 34582 21978
rect 34634 21926 34686 21978
rect 34738 21926 34768 21978
rect 1344 21892 34768 21926
rect 3614 21810 3666 21822
rect 5518 21810 5570 21822
rect 5058 21758 5070 21810
rect 5122 21758 5134 21810
rect 3614 21746 3666 21758
rect 5518 21746 5570 21758
rect 11230 21810 11282 21822
rect 11230 21746 11282 21758
rect 11342 21810 11394 21822
rect 11342 21746 11394 21758
rect 12686 21810 12738 21822
rect 12686 21746 12738 21758
rect 13582 21810 13634 21822
rect 13582 21746 13634 21758
rect 13694 21810 13746 21822
rect 13694 21746 13746 21758
rect 13806 21810 13858 21822
rect 13806 21746 13858 21758
rect 14702 21810 14754 21822
rect 14702 21746 14754 21758
rect 14926 21810 14978 21822
rect 14926 21746 14978 21758
rect 15710 21810 15762 21822
rect 15710 21746 15762 21758
rect 16382 21810 16434 21822
rect 19406 21810 19458 21822
rect 17938 21758 17950 21810
rect 18002 21758 18014 21810
rect 16382 21746 16434 21758
rect 19406 21746 19458 21758
rect 19966 21810 20018 21822
rect 19966 21746 20018 21758
rect 20862 21810 20914 21822
rect 20862 21746 20914 21758
rect 20974 21810 21026 21822
rect 25454 21810 25506 21822
rect 24434 21758 24446 21810
rect 24498 21758 24510 21810
rect 20974 21746 21026 21758
rect 25454 21746 25506 21758
rect 3950 21698 4002 21710
rect 3950 21634 4002 21646
rect 4622 21698 4674 21710
rect 4622 21634 4674 21646
rect 5406 21698 5458 21710
rect 5406 21634 5458 21646
rect 10782 21698 10834 21710
rect 13470 21698 13522 21710
rect 12338 21646 12350 21698
rect 12402 21646 12414 21698
rect 10782 21634 10834 21646
rect 13470 21634 13522 21646
rect 14814 21698 14866 21710
rect 14814 21634 14866 21646
rect 16718 21698 16770 21710
rect 16718 21634 16770 21646
rect 19294 21698 19346 21710
rect 19294 21634 19346 21646
rect 20526 21698 20578 21710
rect 20526 21634 20578 21646
rect 20750 21698 20802 21710
rect 20750 21634 20802 21646
rect 21646 21698 21698 21710
rect 21646 21634 21698 21646
rect 25566 21698 25618 21710
rect 25566 21634 25618 21646
rect 3390 21586 3442 21598
rect 3390 21522 3442 21534
rect 3614 21586 3666 21598
rect 3614 21522 3666 21534
rect 4398 21586 4450 21598
rect 4398 21522 4450 21534
rect 4510 21586 4562 21598
rect 4510 21522 4562 21534
rect 5742 21586 5794 21598
rect 5742 21522 5794 21534
rect 10558 21586 10610 21598
rect 10558 21522 10610 21534
rect 10894 21586 10946 21598
rect 11902 21586 11954 21598
rect 15150 21586 15202 21598
rect 17614 21586 17666 21598
rect 19630 21586 19682 21598
rect 11554 21534 11566 21586
rect 11618 21534 11630 21586
rect 13122 21534 13134 21586
rect 13186 21534 13198 21586
rect 14130 21534 14142 21586
rect 14194 21534 14206 21586
rect 14466 21534 14478 21586
rect 14530 21534 14542 21586
rect 15474 21534 15486 21586
rect 15538 21534 15550 21586
rect 18162 21534 18174 21586
rect 18226 21534 18238 21586
rect 10894 21522 10946 21534
rect 11902 21522 11954 21534
rect 15150 21522 15202 21534
rect 17614 21522 17666 21534
rect 19630 21522 19682 21534
rect 20190 21586 20242 21598
rect 20190 21522 20242 21534
rect 21198 21586 21250 21598
rect 21198 21522 21250 21534
rect 21758 21586 21810 21598
rect 21758 21522 21810 21534
rect 21982 21586 22034 21598
rect 23874 21534 23886 21586
rect 23938 21534 23950 21586
rect 24434 21534 24446 21586
rect 24498 21534 24510 21586
rect 29698 21534 29710 21586
rect 29762 21534 29774 21586
rect 21982 21522 22034 21534
rect 15374 21474 15426 21486
rect 22754 21422 22766 21474
rect 22818 21422 22830 21474
rect 24658 21422 24670 21474
rect 24722 21422 24734 21474
rect 26114 21422 26126 21474
rect 26178 21422 26190 21474
rect 28802 21422 28814 21474
rect 28866 21422 28878 21474
rect 15374 21410 15426 21422
rect 25454 21362 25506 21374
rect 17266 21310 17278 21362
rect 17330 21359 17342 21362
rect 17714 21359 17726 21362
rect 17330 21313 17726 21359
rect 17330 21310 17342 21313
rect 17714 21310 17726 21313
rect 17778 21310 17790 21362
rect 25454 21298 25506 21310
rect 1344 21194 34608 21228
rect 1344 21142 5372 21194
rect 5424 21142 5476 21194
rect 5528 21142 5580 21194
rect 5632 21142 13688 21194
rect 13740 21142 13792 21194
rect 13844 21142 13896 21194
rect 13948 21142 22004 21194
rect 22056 21142 22108 21194
rect 22160 21142 22212 21194
rect 22264 21142 30320 21194
rect 30372 21142 30424 21194
rect 30476 21142 30528 21194
rect 30580 21142 34608 21194
rect 1344 21108 34608 21142
rect 2606 21026 2658 21038
rect 2606 20962 2658 20974
rect 11454 21026 11506 21038
rect 11454 20962 11506 20974
rect 12798 21026 12850 21038
rect 12798 20962 12850 20974
rect 22542 21026 22594 21038
rect 22542 20962 22594 20974
rect 12350 20914 12402 20926
rect 10994 20862 11006 20914
rect 11058 20862 11070 20914
rect 12350 20850 12402 20862
rect 15822 20914 15874 20926
rect 15822 20850 15874 20862
rect 22654 20914 22706 20926
rect 27470 20914 27522 20926
rect 26002 20862 26014 20914
rect 26066 20862 26078 20914
rect 22654 20850 22706 20862
rect 27470 20850 27522 20862
rect 3278 20802 3330 20814
rect 3278 20738 3330 20750
rect 4958 20802 5010 20814
rect 13806 20802 13858 20814
rect 16046 20802 16098 20814
rect 27022 20802 27074 20814
rect 5618 20750 5630 20802
rect 5682 20750 5694 20802
rect 7634 20750 7646 20802
rect 7698 20750 7710 20802
rect 14130 20750 14142 20802
rect 14194 20750 14206 20802
rect 17602 20750 17614 20802
rect 17666 20750 17678 20802
rect 18162 20750 18174 20802
rect 18226 20750 18238 20802
rect 22866 20750 22878 20802
rect 22930 20750 22942 20802
rect 4958 20738 5010 20750
rect 13806 20738 13858 20750
rect 16046 20738 16098 20750
rect 27022 20738 27074 20750
rect 27358 20802 27410 20814
rect 27358 20738 27410 20750
rect 27582 20802 27634 20814
rect 27582 20738 27634 20750
rect 3950 20690 4002 20702
rect 8206 20690 8258 20702
rect 5730 20638 5742 20690
rect 5794 20638 5806 20690
rect 3950 20626 4002 20638
rect 8206 20626 8258 20638
rect 10558 20690 10610 20702
rect 11342 20690 11394 20702
rect 10658 20638 10670 20690
rect 10722 20638 10734 20690
rect 10558 20626 10610 20638
rect 11342 20626 11394 20638
rect 12686 20690 12738 20702
rect 12686 20626 12738 20638
rect 13470 20690 13522 20702
rect 13470 20626 13522 20638
rect 13582 20690 13634 20702
rect 13582 20626 13634 20638
rect 14366 20690 14418 20702
rect 14366 20626 14418 20638
rect 17390 20690 17442 20702
rect 23762 20638 23774 20690
rect 23826 20638 23838 20690
rect 17390 20626 17442 20638
rect 2382 20578 2434 20590
rect 2382 20514 2434 20526
rect 2494 20578 2546 20590
rect 3614 20578 3666 20590
rect 2930 20526 2942 20578
rect 2994 20526 3006 20578
rect 2494 20514 2546 20526
rect 3614 20514 3666 20526
rect 4286 20578 4338 20590
rect 4286 20514 4338 20526
rect 4398 20578 4450 20590
rect 4398 20514 4450 20526
rect 4510 20578 4562 20590
rect 4510 20514 4562 20526
rect 8094 20578 8146 20590
rect 8094 20514 8146 20526
rect 10222 20578 10274 20590
rect 10222 20514 10274 20526
rect 10446 20578 10498 20590
rect 10446 20514 10498 20526
rect 11454 20578 11506 20590
rect 11454 20514 11506 20526
rect 12798 20578 12850 20590
rect 21422 20578 21474 20590
rect 16370 20526 16382 20578
rect 16434 20526 16446 20578
rect 18386 20526 18398 20578
rect 18450 20526 18462 20578
rect 12798 20514 12850 20526
rect 21422 20514 21474 20526
rect 1344 20410 34768 20444
rect 1344 20358 9530 20410
rect 9582 20358 9634 20410
rect 9686 20358 9738 20410
rect 9790 20358 17846 20410
rect 17898 20358 17950 20410
rect 18002 20358 18054 20410
rect 18106 20358 26162 20410
rect 26214 20358 26266 20410
rect 26318 20358 26370 20410
rect 26422 20358 34478 20410
rect 34530 20358 34582 20410
rect 34634 20358 34686 20410
rect 34738 20358 34768 20410
rect 1344 20324 34768 20358
rect 12798 20242 12850 20254
rect 12798 20178 12850 20190
rect 26686 20242 26738 20254
rect 26686 20178 26738 20190
rect 8206 20130 8258 20142
rect 2482 20078 2494 20130
rect 2546 20078 2558 20130
rect 8206 20066 8258 20078
rect 8878 20130 8930 20142
rect 12014 20130 12066 20142
rect 10322 20078 10334 20130
rect 10386 20078 10398 20130
rect 8878 20066 8930 20078
rect 12014 20066 12066 20078
rect 12462 20130 12514 20142
rect 12462 20066 12514 20078
rect 12574 20130 12626 20142
rect 23998 20130 24050 20142
rect 14018 20078 14030 20130
rect 14082 20078 14094 20130
rect 15026 20078 15038 20130
rect 15090 20078 15102 20130
rect 15362 20078 15374 20130
rect 15426 20078 15438 20130
rect 16818 20078 16830 20130
rect 16882 20078 16894 20130
rect 12574 20066 12626 20078
rect 23998 20066 24050 20078
rect 24446 20130 24498 20142
rect 24446 20066 24498 20078
rect 4846 20018 4898 20030
rect 1810 19966 1822 20018
rect 1874 19966 1886 20018
rect 4846 19954 4898 19966
rect 5182 20018 5234 20030
rect 5182 19954 5234 19966
rect 5406 20018 5458 20030
rect 10558 20018 10610 20030
rect 11454 20018 11506 20030
rect 7746 19966 7758 20018
rect 7810 19966 7822 20018
rect 9762 19966 9774 20018
rect 9826 19966 9838 20018
rect 10770 19966 10782 20018
rect 10834 19966 10846 20018
rect 5406 19954 5458 19966
rect 10558 19954 10610 19966
rect 11454 19954 11506 19966
rect 11902 20018 11954 20030
rect 11902 19954 11954 19966
rect 12126 20018 12178 20030
rect 15710 20018 15762 20030
rect 18062 20018 18114 20030
rect 14242 19966 14254 20018
rect 14306 19966 14318 20018
rect 14802 19966 14814 20018
rect 14866 19966 14878 20018
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 17714 19966 17726 20018
rect 17778 19966 17790 20018
rect 12126 19954 12178 19966
rect 15710 19954 15762 19966
rect 18062 19954 18114 19966
rect 18174 20018 18226 20030
rect 18174 19954 18226 19966
rect 18286 20018 18338 20030
rect 18286 19954 18338 19966
rect 18622 20018 18674 20030
rect 18622 19954 18674 19966
rect 18958 20018 19010 20030
rect 18958 19954 19010 19966
rect 19182 20018 19234 20030
rect 19182 19954 19234 19966
rect 20638 20018 20690 20030
rect 24670 20018 24722 20030
rect 21074 19966 21086 20018
rect 21138 19966 21150 20018
rect 22194 19966 22206 20018
rect 22258 19966 22270 20018
rect 22978 19966 22990 20018
rect 23042 19966 23054 20018
rect 20638 19954 20690 19966
rect 24670 19954 24722 19966
rect 25230 20018 25282 20030
rect 25890 19966 25902 20018
rect 25954 19966 25966 20018
rect 27122 19966 27134 20018
rect 27186 19966 27198 20018
rect 30594 19966 30606 20018
rect 30658 19966 30670 20018
rect 25230 19954 25282 19966
rect 5070 19906 5122 19918
rect 16158 19906 16210 19918
rect 4610 19854 4622 19906
rect 4674 19854 4686 19906
rect 7298 19854 7310 19906
rect 7362 19854 7374 19906
rect 9650 19854 9662 19906
rect 9714 19854 9726 19906
rect 5070 19842 5122 19854
rect 16158 19842 16210 19854
rect 19070 19906 19122 19918
rect 19070 19842 19122 19854
rect 21534 19906 21586 19918
rect 21534 19842 21586 19854
rect 21870 19906 21922 19918
rect 24322 19854 24334 19906
rect 24386 19854 24398 19906
rect 25666 19854 25678 19906
rect 25730 19854 25742 19906
rect 27794 19854 27806 19906
rect 27858 19854 27870 19906
rect 29922 19854 29934 19906
rect 29986 19854 29998 19906
rect 21870 19842 21922 19854
rect 8654 19794 8706 19806
rect 8654 19730 8706 19742
rect 8990 19794 9042 19806
rect 8990 19730 9042 19742
rect 22206 19794 22258 19806
rect 22206 19730 22258 19742
rect 27134 19794 27186 19806
rect 27134 19730 27186 19742
rect 27470 19794 27522 19806
rect 27470 19730 27522 19742
rect 1344 19626 34608 19660
rect 1344 19574 5372 19626
rect 5424 19574 5476 19626
rect 5528 19574 5580 19626
rect 5632 19574 13688 19626
rect 13740 19574 13792 19626
rect 13844 19574 13896 19626
rect 13948 19574 22004 19626
rect 22056 19574 22108 19626
rect 22160 19574 22212 19626
rect 22264 19574 30320 19626
rect 30372 19574 30424 19626
rect 30476 19574 30528 19626
rect 30580 19574 34608 19626
rect 1344 19540 34608 19574
rect 12686 19458 12738 19470
rect 12686 19394 12738 19406
rect 17614 19458 17666 19470
rect 17614 19394 17666 19406
rect 7982 19346 8034 19358
rect 2482 19294 2494 19346
rect 2546 19294 2558 19346
rect 4610 19294 4622 19346
rect 4674 19294 4686 19346
rect 7982 19282 8034 19294
rect 8990 19346 9042 19358
rect 8990 19282 9042 19294
rect 9438 19346 9490 19358
rect 9438 19282 9490 19294
rect 9774 19346 9826 19358
rect 9774 19282 9826 19294
rect 11342 19346 11394 19358
rect 11342 19282 11394 19294
rect 17390 19346 17442 19358
rect 17390 19282 17442 19294
rect 18398 19346 18450 19358
rect 22306 19294 22318 19346
rect 22370 19294 22382 19346
rect 24546 19294 24558 19346
rect 24610 19294 24622 19346
rect 26450 19294 26462 19346
rect 26514 19294 26526 19346
rect 28578 19294 28590 19346
rect 28642 19294 28654 19346
rect 18398 19282 18450 19294
rect 7086 19234 7138 19246
rect 8654 19234 8706 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 7522 19182 7534 19234
rect 7586 19182 7598 19234
rect 7086 19170 7138 19182
rect 8654 19170 8706 19182
rect 8878 19234 8930 19246
rect 8878 19170 8930 19182
rect 9214 19234 9266 19246
rect 9214 19170 9266 19182
rect 10782 19234 10834 19246
rect 10782 19170 10834 19182
rect 12238 19234 12290 19246
rect 29150 19234 29202 19246
rect 21634 19182 21646 19234
rect 21698 19182 21710 19234
rect 25666 19182 25678 19234
rect 25730 19182 25742 19234
rect 12238 19170 12290 19182
rect 29150 19170 29202 19182
rect 29822 19234 29874 19246
rect 29822 19170 29874 19182
rect 9998 19122 10050 19134
rect 9998 19058 10050 19070
rect 10558 19122 10610 19134
rect 10558 19058 10610 19070
rect 11230 19122 11282 19134
rect 11230 19058 11282 19070
rect 12798 19122 12850 19134
rect 12798 19058 12850 19070
rect 15038 19122 15090 19134
rect 15038 19058 15090 19070
rect 11006 19010 11058 19022
rect 11006 18946 11058 18958
rect 11902 19010 11954 19022
rect 11902 18946 11954 18958
rect 12126 19010 12178 19022
rect 12126 18946 12178 18958
rect 12350 19010 12402 19022
rect 29262 19010 29314 19022
rect 17938 18958 17950 19010
rect 18002 18958 18014 19010
rect 12350 18946 12402 18958
rect 29262 18946 29314 18958
rect 29374 19010 29426 19022
rect 29374 18946 29426 18958
rect 1344 18842 34768 18876
rect 1344 18790 9530 18842
rect 9582 18790 9634 18842
rect 9686 18790 9738 18842
rect 9790 18790 17846 18842
rect 17898 18790 17950 18842
rect 18002 18790 18054 18842
rect 18106 18790 26162 18842
rect 26214 18790 26266 18842
rect 26318 18790 26370 18842
rect 26422 18790 34478 18842
rect 34530 18790 34582 18842
rect 34634 18790 34686 18842
rect 34738 18790 34768 18842
rect 1344 18756 34768 18790
rect 8206 18674 8258 18686
rect 7410 18622 7422 18674
rect 7474 18622 7486 18674
rect 8206 18610 8258 18622
rect 10782 18674 10834 18686
rect 10782 18610 10834 18622
rect 11454 18674 11506 18686
rect 12674 18622 12686 18674
rect 12738 18622 12750 18674
rect 11454 18610 11506 18622
rect 7982 18562 8034 18574
rect 6514 18510 6526 18562
rect 6578 18510 6590 18562
rect 7982 18498 8034 18510
rect 8766 18562 8818 18574
rect 8766 18498 8818 18510
rect 8878 18562 8930 18574
rect 8878 18498 8930 18510
rect 9550 18562 9602 18574
rect 9550 18498 9602 18510
rect 9662 18562 9714 18574
rect 19506 18510 19518 18562
rect 19570 18510 19582 18562
rect 23202 18510 23214 18562
rect 23266 18510 23278 18562
rect 30706 18510 30718 18562
rect 30770 18510 30782 18562
rect 9662 18498 9714 18510
rect 7870 18450 7922 18462
rect 6290 18398 6302 18450
rect 6354 18398 6366 18450
rect 7870 18386 7922 18398
rect 8318 18450 8370 18462
rect 8318 18386 8370 18398
rect 9886 18450 9938 18462
rect 9886 18386 9938 18398
rect 10558 18450 10610 18462
rect 10558 18386 10610 18398
rect 10670 18450 10722 18462
rect 10670 18386 10722 18398
rect 11230 18450 11282 18462
rect 11230 18386 11282 18398
rect 11454 18450 11506 18462
rect 11454 18386 11506 18398
rect 11790 18450 11842 18462
rect 17390 18450 17442 18462
rect 14018 18398 14030 18450
rect 14082 18398 14094 18450
rect 11790 18386 11842 18398
rect 17390 18386 17442 18398
rect 17614 18450 17666 18462
rect 22878 18450 22930 18462
rect 17938 18398 17950 18450
rect 18002 18398 18014 18450
rect 18722 18398 18734 18450
rect 18786 18398 18798 18450
rect 17614 18386 17666 18398
rect 22878 18386 22930 18398
rect 23550 18450 23602 18462
rect 26798 18450 26850 18462
rect 26114 18398 26126 18450
rect 26178 18398 26190 18450
rect 27122 18398 27134 18450
rect 27186 18398 27198 18450
rect 23550 18386 23602 18398
rect 26798 18386 26850 18398
rect 6862 18338 6914 18350
rect 10334 18338 10386 18350
rect 8194 18286 8206 18338
rect 8258 18286 8270 18338
rect 6862 18274 6914 18286
rect 10334 18274 10386 18286
rect 12126 18338 12178 18350
rect 12126 18274 12178 18286
rect 12350 18338 12402 18350
rect 17502 18338 17554 18350
rect 25454 18338 25506 18350
rect 14690 18286 14702 18338
rect 14754 18286 14766 18338
rect 16818 18286 16830 18338
rect 16882 18286 16894 18338
rect 21634 18286 21646 18338
rect 21698 18286 21710 18338
rect 25890 18286 25902 18338
rect 25954 18286 25966 18338
rect 12350 18274 12402 18286
rect 17502 18274 17554 18286
rect 25454 18274 25506 18286
rect 7086 18226 7138 18238
rect 7086 18162 7138 18174
rect 8878 18226 8930 18238
rect 8878 18162 8930 18174
rect 10110 18226 10162 18238
rect 10110 18162 10162 18174
rect 1344 18058 34608 18092
rect 1344 18006 5372 18058
rect 5424 18006 5476 18058
rect 5528 18006 5580 18058
rect 5632 18006 13688 18058
rect 13740 18006 13792 18058
rect 13844 18006 13896 18058
rect 13948 18006 22004 18058
rect 22056 18006 22108 18058
rect 22160 18006 22212 18058
rect 22264 18006 30320 18058
rect 30372 18006 30424 18058
rect 30476 18006 30528 18058
rect 30580 18006 34608 18058
rect 1344 17972 34608 18006
rect 9550 17890 9602 17902
rect 6850 17838 6862 17890
rect 6914 17838 6926 17890
rect 9550 17826 9602 17838
rect 9886 17890 9938 17902
rect 9886 17826 9938 17838
rect 10782 17890 10834 17902
rect 29698 17838 29710 17890
rect 29762 17838 29774 17890
rect 10782 17826 10834 17838
rect 8430 17778 8482 17790
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 8430 17714 8482 17726
rect 16046 17778 16098 17790
rect 16046 17714 16098 17726
rect 17054 17778 17106 17790
rect 23538 17726 23550 17778
rect 23602 17726 23614 17778
rect 33282 17726 33294 17778
rect 33346 17726 33358 17778
rect 17054 17714 17106 17726
rect 6302 17666 6354 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 5730 17614 5742 17666
rect 5794 17614 5806 17666
rect 6302 17602 6354 17614
rect 6526 17666 6578 17678
rect 6526 17602 6578 17614
rect 7646 17666 7698 17678
rect 10894 17666 10946 17678
rect 7858 17614 7870 17666
rect 7922 17614 7934 17666
rect 9090 17614 9102 17666
rect 9154 17614 9166 17666
rect 10210 17614 10222 17666
rect 10274 17614 10286 17666
rect 7646 17602 7698 17614
rect 10894 17602 10946 17614
rect 15822 17666 15874 17678
rect 15822 17602 15874 17614
rect 16158 17666 16210 17678
rect 16158 17602 16210 17614
rect 16494 17666 16546 17678
rect 29374 17666 29426 17678
rect 26674 17614 26686 17666
rect 26738 17614 26750 17666
rect 30482 17614 30494 17666
rect 30546 17614 30558 17666
rect 16494 17602 16546 17614
rect 29374 17602 29426 17614
rect 7198 17554 7250 17566
rect 2482 17502 2494 17554
rect 2546 17502 2558 17554
rect 5954 17502 5966 17554
rect 6018 17502 6030 17554
rect 7198 17490 7250 17502
rect 9774 17554 9826 17566
rect 9774 17490 9826 17502
rect 10670 17554 10722 17566
rect 10670 17490 10722 17502
rect 11230 17554 11282 17566
rect 18958 17554 19010 17566
rect 17490 17502 17502 17554
rect 17554 17502 17566 17554
rect 18162 17502 18174 17554
rect 18226 17502 18238 17554
rect 11230 17490 11282 17502
rect 18958 17490 19010 17502
rect 29150 17554 29202 17566
rect 31154 17502 31166 17554
rect 31218 17502 31230 17554
rect 29150 17490 29202 17502
rect 5070 17442 5122 17454
rect 5070 17378 5122 17390
rect 7310 17442 7362 17454
rect 10446 17442 10498 17454
rect 8866 17390 8878 17442
rect 8930 17390 8942 17442
rect 7310 17378 7362 17390
rect 10446 17378 10498 17390
rect 11118 17442 11170 17454
rect 11118 17378 11170 17390
rect 17838 17442 17890 17454
rect 17838 17378 17890 17390
rect 18510 17442 18562 17454
rect 18510 17378 18562 17390
rect 19070 17442 19122 17454
rect 19070 17378 19122 17390
rect 22542 17442 22594 17454
rect 22542 17378 22594 17390
rect 1344 17274 34768 17308
rect 1344 17222 9530 17274
rect 9582 17222 9634 17274
rect 9686 17222 9738 17274
rect 9790 17222 17846 17274
rect 17898 17222 17950 17274
rect 18002 17222 18054 17274
rect 18106 17222 26162 17274
rect 26214 17222 26266 17274
rect 26318 17222 26370 17274
rect 26422 17222 34478 17274
rect 34530 17222 34582 17274
rect 34634 17222 34686 17274
rect 34738 17222 34768 17274
rect 1344 17188 34768 17222
rect 7646 17106 7698 17118
rect 7074 17054 7086 17106
rect 7138 17054 7150 17106
rect 7646 17042 7698 17054
rect 8206 17106 8258 17118
rect 8206 17042 8258 17054
rect 8430 17106 8482 17118
rect 14366 17106 14418 17118
rect 8642 17054 8654 17106
rect 8706 17054 8718 17106
rect 9874 17054 9886 17106
rect 9938 17054 9950 17106
rect 8430 17042 8482 17054
rect 14366 17042 14418 17054
rect 15262 17106 15314 17118
rect 15262 17042 15314 17054
rect 15822 17106 15874 17118
rect 15822 17042 15874 17054
rect 17390 17106 17442 17118
rect 17390 17042 17442 17054
rect 29598 17106 29650 17118
rect 29598 17042 29650 17054
rect 30046 17106 30098 17118
rect 30046 17042 30098 17054
rect 31950 17106 32002 17118
rect 31950 17042 32002 17054
rect 6750 16994 6802 17006
rect 6750 16930 6802 16942
rect 8094 16994 8146 17006
rect 8094 16930 8146 16942
rect 14142 16994 14194 17006
rect 14142 16930 14194 16942
rect 15934 16994 15986 17006
rect 15934 16930 15986 16942
rect 16718 16994 16770 17006
rect 16718 16930 16770 16942
rect 17614 16994 17666 17006
rect 17614 16930 17666 16942
rect 17726 16994 17778 17006
rect 29374 16994 29426 17006
rect 17938 16942 17950 16994
rect 18002 16942 18014 16994
rect 20626 16942 20638 16994
rect 20690 16942 20702 16994
rect 30370 16942 30382 16994
rect 30434 16942 30446 16994
rect 17726 16930 17778 16942
rect 29374 16930 29426 16942
rect 7534 16882 7586 16894
rect 9550 16882 9602 16894
rect 3266 16830 3278 16882
rect 3330 16830 3342 16882
rect 3938 16830 3950 16882
rect 4002 16830 4014 16882
rect 8866 16830 8878 16882
rect 8930 16830 8942 16882
rect 7534 16818 7586 16830
rect 9550 16818 9602 16830
rect 12238 16882 12290 16894
rect 12238 16818 12290 16830
rect 12350 16882 12402 16894
rect 15374 16882 15426 16894
rect 13570 16830 13582 16882
rect 13634 16830 13646 16882
rect 13906 16830 13918 16882
rect 13970 16830 13982 16882
rect 12350 16818 12402 16830
rect 15374 16818 15426 16830
rect 15710 16882 15762 16894
rect 15710 16818 15762 16830
rect 16382 16882 16434 16894
rect 16382 16818 16434 16830
rect 16830 16882 16882 16894
rect 29262 16882 29314 16894
rect 21298 16830 21310 16882
rect 21362 16830 21374 16882
rect 24546 16830 24558 16882
rect 24610 16830 24622 16882
rect 25330 16830 25342 16882
rect 25394 16830 25406 16882
rect 16830 16818 16882 16830
rect 29262 16818 29314 16830
rect 29710 16882 29762 16894
rect 29710 16818 29762 16830
rect 31502 16882 31554 16894
rect 31502 16818 31554 16830
rect 32174 16882 32226 16894
rect 32174 16818 32226 16830
rect 12798 16770 12850 16782
rect 32062 16770 32114 16782
rect 6066 16718 6078 16770
rect 6130 16718 6142 16770
rect 14018 16718 14030 16770
rect 14082 16718 14094 16770
rect 18162 16718 18174 16770
rect 18226 16718 18238 16770
rect 18498 16718 18510 16770
rect 18562 16718 18574 16770
rect 21746 16718 21758 16770
rect 21810 16718 21822 16770
rect 23874 16718 23886 16770
rect 23938 16718 23950 16770
rect 26002 16718 26014 16770
rect 26066 16718 26078 16770
rect 28130 16718 28142 16770
rect 28194 16718 28206 16770
rect 12798 16706 12850 16718
rect 32062 16706 32114 16718
rect 7646 16658 7698 16670
rect 7646 16594 7698 16606
rect 12686 16658 12738 16670
rect 12686 16594 12738 16606
rect 15262 16658 15314 16670
rect 15262 16594 15314 16606
rect 16718 16658 16770 16670
rect 16718 16594 16770 16606
rect 1344 16490 34608 16524
rect 1344 16438 5372 16490
rect 5424 16438 5476 16490
rect 5528 16438 5580 16490
rect 5632 16438 13688 16490
rect 13740 16438 13792 16490
rect 13844 16438 13896 16490
rect 13948 16438 22004 16490
rect 22056 16438 22108 16490
rect 22160 16438 22212 16490
rect 22264 16438 30320 16490
rect 30372 16438 30424 16490
rect 30476 16438 30528 16490
rect 30580 16438 34608 16490
rect 1344 16404 34608 16438
rect 17950 16322 18002 16334
rect 17950 16258 18002 16270
rect 27470 16322 27522 16334
rect 27470 16258 27522 16270
rect 30158 16322 30210 16334
rect 30158 16258 30210 16270
rect 23438 16210 23490 16222
rect 5058 16158 5070 16210
rect 5122 16158 5134 16210
rect 10770 16158 10782 16210
rect 10834 16158 10846 16210
rect 12898 16158 12910 16210
rect 12962 16158 12974 16210
rect 13682 16158 13694 16210
rect 13746 16158 13758 16210
rect 17378 16158 17390 16210
rect 17442 16158 17454 16210
rect 23438 16146 23490 16158
rect 24446 16210 24498 16222
rect 24446 16146 24498 16158
rect 29262 16210 29314 16222
rect 34178 16158 34190 16210
rect 34242 16158 34254 16210
rect 29262 16146 29314 16158
rect 15150 16098 15202 16110
rect 2258 16046 2270 16098
rect 2322 16046 2334 16098
rect 9986 16046 9998 16098
rect 10050 16046 10062 16098
rect 13794 16046 13806 16098
rect 13858 16046 13870 16098
rect 15150 16034 15202 16046
rect 15486 16098 15538 16110
rect 15486 16034 15538 16046
rect 15710 16098 15762 16110
rect 15710 16034 15762 16046
rect 15934 16098 15986 16110
rect 15934 16034 15986 16046
rect 16158 16098 16210 16110
rect 16158 16034 16210 16046
rect 16606 16098 16658 16110
rect 17726 16098 17778 16110
rect 22430 16098 22482 16110
rect 17266 16046 17278 16098
rect 17330 16046 17342 16098
rect 19282 16046 19294 16098
rect 19346 16046 19358 16098
rect 21858 16046 21870 16098
rect 21922 16046 21934 16098
rect 16606 16034 16658 16046
rect 17726 16034 17778 16046
rect 22430 16034 22482 16046
rect 23662 16098 23714 16110
rect 23662 16034 23714 16046
rect 26238 16098 26290 16110
rect 26238 16034 26290 16046
rect 27582 16098 27634 16110
rect 27582 16034 27634 16046
rect 29374 16098 29426 16110
rect 29374 16034 29426 16046
rect 29822 16098 29874 16110
rect 31266 16046 31278 16098
rect 31330 16046 31342 16098
rect 29822 16034 29874 16046
rect 14142 15986 14194 15998
rect 2930 15934 2942 15986
rect 2994 15934 3006 15986
rect 14142 15922 14194 15934
rect 14814 15986 14866 15998
rect 14814 15922 14866 15934
rect 15038 15986 15090 15998
rect 15038 15922 15090 15934
rect 16046 15986 16098 15998
rect 16046 15922 16098 15934
rect 16942 15986 16994 15998
rect 16942 15922 16994 15934
rect 18734 15986 18786 15998
rect 18734 15922 18786 15934
rect 21534 15986 21586 15998
rect 21534 15922 21586 15934
rect 22206 15986 22258 15998
rect 22206 15922 22258 15934
rect 22654 15986 22706 15998
rect 22654 15922 22706 15934
rect 22766 15986 22818 15998
rect 22766 15922 22818 15934
rect 24334 15986 24386 15998
rect 24334 15922 24386 15934
rect 24558 15986 24610 15998
rect 24558 15922 24610 15934
rect 26126 15986 26178 15998
rect 26126 15922 26178 15934
rect 27918 15986 27970 15998
rect 27918 15922 27970 15934
rect 28366 15986 28418 15998
rect 28366 15922 28418 15934
rect 29150 15986 29202 15998
rect 29150 15922 29202 15934
rect 30046 15986 30098 15998
rect 32050 15934 32062 15986
rect 32114 15934 32126 15986
rect 30046 15922 30098 15934
rect 5742 15874 5794 15886
rect 5742 15810 5794 15822
rect 6302 15874 6354 15886
rect 6302 15810 6354 15822
rect 9662 15874 9714 15886
rect 9662 15810 9714 15822
rect 14254 15874 14306 15886
rect 14254 15810 14306 15822
rect 14478 15874 14530 15886
rect 14478 15810 14530 15822
rect 16830 15874 16882 15886
rect 16830 15810 16882 15822
rect 18286 15874 18338 15886
rect 18286 15810 18338 15822
rect 18846 15874 18898 15886
rect 18846 15810 18898 15822
rect 19070 15874 19122 15886
rect 19070 15810 19122 15822
rect 21646 15874 21698 15886
rect 26014 15874 26066 15886
rect 23986 15822 23998 15874
rect 24050 15822 24062 15874
rect 21646 15810 21698 15822
rect 26014 15810 26066 15822
rect 27470 15874 27522 15886
rect 27470 15810 27522 15822
rect 28142 15874 28194 15886
rect 28142 15810 28194 15822
rect 28478 15874 28530 15886
rect 28478 15810 28530 15822
rect 1344 15706 34768 15740
rect 1344 15654 9530 15706
rect 9582 15654 9634 15706
rect 9686 15654 9738 15706
rect 9790 15654 17846 15706
rect 17898 15654 17950 15706
rect 18002 15654 18054 15706
rect 18106 15654 26162 15706
rect 26214 15654 26266 15706
rect 26318 15654 26370 15706
rect 26422 15654 34478 15706
rect 34530 15654 34582 15706
rect 34634 15654 34686 15706
rect 34738 15654 34768 15706
rect 1344 15620 34768 15654
rect 14926 15538 14978 15550
rect 14926 15474 14978 15486
rect 15486 15538 15538 15550
rect 15486 15474 15538 15486
rect 15710 15538 15762 15550
rect 15710 15474 15762 15486
rect 30382 15538 30434 15550
rect 33058 15486 33070 15538
rect 33122 15486 33134 15538
rect 30382 15474 30434 15486
rect 16270 15426 16322 15438
rect 11890 15374 11902 15426
rect 11954 15374 11966 15426
rect 16270 15362 16322 15374
rect 16718 15426 16770 15438
rect 16718 15362 16770 15374
rect 16830 15426 16882 15438
rect 26126 15426 26178 15438
rect 20178 15374 20190 15426
rect 20242 15374 20254 15426
rect 16830 15362 16882 15374
rect 26126 15362 26178 15374
rect 26350 15426 26402 15438
rect 26350 15362 26402 15374
rect 30942 15426 30994 15438
rect 30942 15362 30994 15374
rect 32062 15426 32114 15438
rect 32062 15362 32114 15374
rect 32286 15426 32338 15438
rect 32286 15362 32338 15374
rect 8990 15314 9042 15326
rect 14814 15314 14866 15326
rect 17950 15314 18002 15326
rect 31054 15314 31106 15326
rect 5730 15262 5742 15314
rect 5794 15262 5806 15314
rect 11218 15262 11230 15314
rect 11282 15262 11294 15314
rect 15250 15262 15262 15314
rect 15314 15262 15326 15314
rect 15922 15262 15934 15314
rect 15986 15262 15998 15314
rect 18162 15262 18174 15314
rect 18226 15262 18238 15314
rect 28802 15262 28814 15314
rect 28866 15262 28878 15314
rect 8990 15250 9042 15262
rect 14814 15250 14866 15262
rect 17950 15250 18002 15262
rect 31054 15250 31106 15262
rect 31502 15314 31554 15326
rect 33630 15314 33682 15326
rect 31714 15262 31726 15314
rect 31778 15262 31790 15314
rect 31502 15250 31554 15262
rect 33630 15250 33682 15262
rect 30494 15202 30546 15214
rect 6402 15150 6414 15202
rect 6466 15150 6478 15202
rect 8530 15150 8542 15202
rect 8594 15150 8606 15202
rect 14018 15150 14030 15202
rect 14082 15150 14094 15202
rect 15362 15150 15374 15202
rect 15426 15150 15438 15202
rect 26002 15150 26014 15202
rect 26066 15150 26078 15202
rect 30494 15138 30546 15150
rect 30606 15202 30658 15214
rect 33406 15202 33458 15214
rect 32386 15150 32398 15202
rect 32450 15150 32462 15202
rect 30606 15138 30658 15150
rect 33406 15138 33458 15150
rect 16382 15090 16434 15102
rect 16382 15026 16434 15038
rect 28478 15090 28530 15102
rect 28478 15026 28530 15038
rect 28814 15090 28866 15102
rect 28814 15026 28866 15038
rect 31278 15090 31330 15102
rect 31278 15026 31330 15038
rect 1344 14922 34608 14956
rect 1344 14870 5372 14922
rect 5424 14870 5476 14922
rect 5528 14870 5580 14922
rect 5632 14870 13688 14922
rect 13740 14870 13792 14922
rect 13844 14870 13896 14922
rect 13948 14870 22004 14922
rect 22056 14870 22108 14922
rect 22160 14870 22212 14922
rect 22264 14870 30320 14922
rect 30372 14870 30424 14922
rect 30476 14870 30528 14922
rect 30580 14870 34608 14922
rect 1344 14836 34608 14870
rect 30830 14754 30882 14766
rect 32734 14754 32786 14766
rect 18610 14702 18622 14754
rect 18674 14702 18686 14754
rect 28242 14702 28254 14754
rect 28306 14702 28318 14754
rect 32162 14702 32174 14754
rect 32226 14702 32238 14754
rect 30830 14690 30882 14702
rect 32734 14690 32786 14702
rect 32846 14754 32898 14766
rect 32846 14690 32898 14702
rect 4610 14590 4622 14642
rect 4674 14590 4686 14642
rect 18722 14590 18734 14642
rect 18786 14590 18798 14642
rect 20626 14590 20638 14642
rect 20690 14590 20702 14642
rect 21298 14590 21310 14642
rect 21362 14590 21374 14642
rect 23426 14590 23438 14642
rect 23490 14590 23502 14642
rect 16158 14530 16210 14542
rect 17278 14530 17330 14542
rect 27246 14530 27298 14542
rect 1810 14478 1822 14530
rect 1874 14478 1886 14530
rect 12674 14478 12686 14530
rect 12738 14478 12750 14530
rect 16930 14478 16942 14530
rect 16994 14478 17006 14530
rect 20738 14478 20750 14530
rect 20802 14478 20814 14530
rect 24210 14478 24222 14530
rect 24274 14478 24286 14530
rect 16158 14466 16210 14478
rect 17278 14466 17330 14478
rect 27246 14466 27298 14478
rect 27582 14530 27634 14542
rect 27582 14466 27634 14478
rect 27806 14530 27858 14542
rect 27806 14466 27858 14478
rect 31166 14530 31218 14542
rect 31166 14466 31218 14478
rect 31278 14530 31330 14542
rect 31278 14466 31330 14478
rect 31614 14530 31666 14542
rect 33070 14530 33122 14542
rect 31826 14478 31838 14530
rect 31890 14478 31902 14530
rect 31614 14466 31666 14478
rect 33070 14466 33122 14478
rect 13582 14418 13634 14430
rect 2482 14366 2494 14418
rect 2546 14366 2558 14418
rect 8418 14366 8430 14418
rect 8482 14366 8494 14418
rect 13582 14354 13634 14366
rect 15822 14418 15874 14430
rect 15822 14354 15874 14366
rect 16494 14418 16546 14430
rect 16494 14354 16546 14366
rect 17726 14418 17778 14430
rect 19518 14418 19570 14430
rect 19058 14366 19070 14418
rect 19122 14366 19134 14418
rect 17726 14354 17778 14366
rect 19518 14354 19570 14366
rect 19630 14418 19682 14430
rect 19630 14354 19682 14366
rect 20078 14418 20130 14430
rect 20078 14354 20130 14366
rect 27470 14418 27522 14430
rect 27470 14354 27522 14366
rect 29150 14418 29202 14430
rect 29150 14354 29202 14366
rect 30718 14418 30770 14430
rect 30718 14354 30770 14366
rect 5070 14306 5122 14318
rect 5070 14242 5122 14254
rect 5630 14306 5682 14318
rect 15934 14306 15986 14318
rect 5954 14254 5966 14306
rect 6018 14254 6030 14306
rect 5630 14242 5682 14254
rect 15934 14242 15986 14254
rect 19854 14306 19906 14318
rect 19854 14242 19906 14254
rect 20302 14306 20354 14318
rect 20302 14242 20354 14254
rect 20526 14306 20578 14318
rect 20526 14242 20578 14254
rect 29486 14306 29538 14318
rect 29486 14242 29538 14254
rect 32734 14306 32786 14318
rect 32734 14242 32786 14254
rect 1344 14138 34768 14172
rect 1344 14086 9530 14138
rect 9582 14086 9634 14138
rect 9686 14086 9738 14138
rect 9790 14086 17846 14138
rect 17898 14086 17950 14138
rect 18002 14086 18054 14138
rect 18106 14086 26162 14138
rect 26214 14086 26266 14138
rect 26318 14086 26370 14138
rect 26422 14086 34478 14138
rect 34530 14086 34582 14138
rect 34634 14086 34686 14138
rect 34738 14086 34768 14138
rect 1344 14052 34768 14086
rect 6750 13970 6802 13982
rect 6750 13906 6802 13918
rect 9774 13970 9826 13982
rect 9774 13906 9826 13918
rect 14142 13970 14194 13982
rect 14142 13906 14194 13918
rect 16830 13970 16882 13982
rect 16830 13906 16882 13918
rect 18398 13970 18450 13982
rect 18398 13906 18450 13918
rect 18846 13970 18898 13982
rect 23662 13970 23714 13982
rect 19842 13918 19854 13970
rect 19906 13918 19918 13970
rect 22866 13918 22878 13970
rect 22930 13918 22942 13970
rect 18846 13906 18898 13918
rect 23662 13906 23714 13918
rect 24222 13970 24274 13982
rect 24222 13906 24274 13918
rect 31166 13970 31218 13982
rect 32274 13918 32286 13970
rect 32338 13918 32350 13970
rect 31166 13906 31218 13918
rect 5966 13858 6018 13870
rect 5966 13794 6018 13806
rect 7310 13858 7362 13870
rect 7310 13794 7362 13806
rect 7422 13858 7474 13870
rect 7422 13794 7474 13806
rect 9998 13858 10050 13870
rect 9998 13794 10050 13806
rect 10110 13858 10162 13870
rect 15934 13858 15986 13870
rect 10882 13806 10894 13858
rect 10946 13806 10958 13858
rect 11106 13806 11118 13858
rect 11170 13806 11182 13858
rect 10110 13794 10162 13806
rect 15934 13794 15986 13806
rect 17390 13858 17442 13870
rect 17390 13794 17442 13806
rect 17726 13858 17778 13870
rect 25678 13858 25730 13870
rect 20514 13806 20526 13858
rect 20578 13806 20590 13858
rect 17726 13794 17778 13806
rect 25678 13794 25730 13806
rect 6302 13746 6354 13758
rect 5506 13694 5518 13746
rect 5570 13694 5582 13746
rect 6302 13682 6354 13694
rect 6526 13746 6578 13758
rect 6526 13682 6578 13694
rect 6862 13746 6914 13758
rect 15822 13746 15874 13758
rect 20190 13746 20242 13758
rect 9538 13694 9550 13746
rect 9602 13694 9614 13746
rect 11330 13694 11342 13746
rect 11394 13694 11406 13746
rect 15250 13694 15262 13746
rect 15314 13694 15326 13746
rect 18162 13694 18174 13746
rect 18226 13694 18238 13746
rect 19618 13694 19630 13746
rect 19682 13694 19694 13746
rect 6862 13682 6914 13694
rect 15822 13682 15874 13694
rect 20190 13682 20242 13694
rect 22206 13746 22258 13758
rect 23550 13746 23602 13758
rect 22642 13694 22654 13746
rect 22706 13694 22718 13746
rect 22206 13682 22258 13694
rect 23550 13682 23602 13694
rect 23886 13746 23938 13758
rect 26126 13746 26178 13758
rect 25442 13694 25454 13746
rect 25506 13694 25518 13746
rect 23886 13682 23938 13694
rect 26126 13682 26178 13694
rect 26350 13746 26402 13758
rect 26350 13682 26402 13694
rect 26686 13746 26738 13758
rect 26686 13682 26738 13694
rect 27022 13746 27074 13758
rect 27022 13682 27074 13694
rect 27358 13746 27410 13758
rect 31726 13746 31778 13758
rect 30706 13694 30718 13746
rect 30770 13694 30782 13746
rect 27358 13682 27410 13694
rect 31726 13682 31778 13694
rect 33182 13746 33234 13758
rect 33182 13682 33234 13694
rect 33630 13746 33682 13758
rect 33630 13682 33682 13694
rect 7758 13634 7810 13646
rect 10222 13634 10274 13646
rect 5618 13582 5630 13634
rect 5682 13582 5694 13634
rect 7970 13582 7982 13634
rect 8034 13582 8046 13634
rect 7758 13570 7810 13582
rect 10222 13570 10274 13582
rect 11902 13634 11954 13646
rect 11902 13570 11954 13582
rect 26462 13634 26514 13646
rect 26462 13570 26514 13582
rect 27246 13634 27298 13646
rect 31278 13634 31330 13646
rect 27794 13582 27806 13634
rect 27858 13582 27870 13634
rect 29922 13582 29934 13634
rect 29986 13582 29998 13634
rect 27246 13570 27298 13582
rect 31278 13570 31330 13582
rect 7310 13522 7362 13534
rect 7310 13458 7362 13470
rect 11790 13522 11842 13534
rect 11790 13458 11842 13470
rect 21310 13522 21362 13534
rect 21310 13458 21362 13470
rect 21758 13522 21810 13534
rect 21758 13458 21810 13470
rect 21982 13522 22034 13534
rect 21982 13458 22034 13470
rect 26910 13522 26962 13534
rect 26910 13458 26962 13470
rect 31390 13522 31442 13534
rect 31390 13458 31442 13470
rect 31950 13522 32002 13534
rect 31950 13458 32002 13470
rect 33294 13522 33346 13534
rect 33294 13458 33346 13470
rect 33518 13522 33570 13534
rect 33518 13458 33570 13470
rect 1344 13354 34608 13388
rect 1344 13302 5372 13354
rect 5424 13302 5476 13354
rect 5528 13302 5580 13354
rect 5632 13302 13688 13354
rect 13740 13302 13792 13354
rect 13844 13302 13896 13354
rect 13948 13302 22004 13354
rect 22056 13302 22108 13354
rect 22160 13302 22212 13354
rect 22264 13302 30320 13354
rect 30372 13302 30424 13354
rect 30476 13302 30528 13354
rect 30580 13302 34608 13354
rect 1344 13268 34608 13302
rect 6526 13186 6578 13198
rect 6526 13122 6578 13134
rect 20302 13186 20354 13198
rect 20302 13122 20354 13134
rect 22094 13186 22146 13198
rect 22094 13122 22146 13134
rect 29598 13186 29650 13198
rect 29598 13122 29650 13134
rect 29710 13186 29762 13198
rect 29710 13122 29762 13134
rect 3726 13074 3778 13086
rect 5630 13074 5682 13086
rect 11230 13074 11282 13086
rect 4610 13022 4622 13074
rect 4674 13022 4686 13074
rect 10770 13022 10782 13074
rect 10834 13022 10846 13074
rect 3726 13010 3778 13022
rect 5630 13010 5682 13022
rect 11230 13010 11282 13022
rect 12126 13074 12178 13086
rect 12126 13010 12178 13022
rect 12574 13074 12626 13086
rect 12574 13010 12626 13022
rect 20078 13074 20130 13086
rect 20078 13010 20130 13022
rect 22990 13074 23042 13086
rect 28590 13074 28642 13086
rect 24770 13022 24782 13074
rect 24834 13022 24846 13074
rect 26898 13022 26910 13074
rect 26962 13022 26974 13074
rect 31266 13022 31278 13074
rect 31330 13022 31342 13074
rect 33394 13022 33406 13074
rect 33458 13022 33470 13074
rect 22990 13010 23042 13022
rect 28590 13010 28642 13022
rect 4286 12962 4338 12974
rect 4286 12898 4338 12910
rect 5854 12962 5906 12974
rect 5854 12898 5906 12910
rect 6078 12962 6130 12974
rect 16942 12962 16994 12974
rect 19518 12962 19570 12974
rect 20862 12962 20914 12974
rect 22318 12962 22370 12974
rect 27470 12962 27522 12974
rect 28366 12962 28418 12974
rect 29374 12962 29426 12974
rect 7858 12910 7870 12962
rect 7922 12910 7934 12962
rect 11666 12910 11678 12962
rect 11730 12910 11742 12962
rect 16034 12910 16046 12962
rect 16098 12910 16110 12962
rect 16594 12910 16606 12962
rect 16658 12910 16670 12962
rect 17602 12910 17614 12962
rect 17666 12910 17678 12962
rect 18274 12910 18286 12962
rect 18338 12910 18350 12962
rect 18946 12910 18958 12962
rect 19010 12910 19022 12962
rect 20514 12910 20526 12962
rect 20578 12910 20590 12962
rect 21858 12910 21870 12962
rect 21922 12910 21934 12962
rect 24098 12910 24110 12962
rect 24162 12910 24174 12962
rect 28018 12910 28030 12962
rect 28082 12910 28094 12962
rect 29138 12910 29150 12962
rect 29202 12910 29214 12962
rect 34066 12910 34078 12962
rect 34130 12910 34142 12962
rect 6078 12898 6130 12910
rect 16942 12898 16994 12910
rect 19518 12898 19570 12910
rect 20862 12898 20914 12910
rect 22318 12898 22370 12910
rect 27470 12898 27522 12910
rect 28366 12898 28418 12910
rect 29374 12898 29426 12910
rect 7534 12850 7586 12862
rect 18622 12850 18674 12862
rect 7186 12798 7198 12850
rect 7250 12798 7262 12850
rect 8642 12798 8654 12850
rect 8706 12798 8718 12850
rect 14130 12798 14142 12850
rect 14194 12798 14206 12850
rect 17378 12798 17390 12850
rect 17442 12798 17454 12850
rect 7534 12786 7586 12798
rect 18622 12786 18674 12798
rect 19854 12850 19906 12862
rect 19854 12786 19906 12798
rect 21646 12850 21698 12862
rect 21646 12786 21698 12798
rect 22542 12850 22594 12862
rect 22542 12786 22594 12798
rect 22878 12850 22930 12862
rect 22878 12786 22930 12798
rect 27358 12850 27410 12862
rect 27358 12786 27410 12798
rect 3390 12738 3442 12750
rect 3390 12674 3442 12686
rect 3614 12738 3666 12750
rect 3614 12674 3666 12686
rect 3838 12738 3890 12750
rect 3838 12674 3890 12686
rect 5070 12738 5122 12750
rect 5070 12674 5122 12686
rect 11118 12738 11170 12750
rect 11118 12674 11170 12686
rect 11342 12738 11394 12750
rect 11342 12674 11394 12686
rect 12014 12738 12066 12750
rect 12014 12674 12066 12686
rect 13806 12738 13858 12750
rect 18510 12738 18562 12750
rect 14578 12686 14590 12738
rect 14642 12686 14654 12738
rect 16258 12686 16270 12738
rect 16322 12686 16334 12738
rect 13806 12674 13858 12686
rect 18510 12674 18562 12686
rect 19294 12738 19346 12750
rect 19294 12674 19346 12686
rect 19406 12738 19458 12750
rect 19406 12674 19458 12686
rect 19742 12738 19794 12750
rect 19742 12674 19794 12686
rect 22094 12738 22146 12750
rect 22094 12674 22146 12686
rect 27134 12738 27186 12750
rect 27134 12674 27186 12686
rect 1344 12570 34768 12604
rect 1344 12518 9530 12570
rect 9582 12518 9634 12570
rect 9686 12518 9738 12570
rect 9790 12518 17846 12570
rect 17898 12518 17950 12570
rect 18002 12518 18054 12570
rect 18106 12518 26162 12570
rect 26214 12518 26266 12570
rect 26318 12518 26370 12570
rect 26422 12518 34478 12570
rect 34530 12518 34582 12570
rect 34634 12518 34686 12570
rect 34738 12518 34768 12570
rect 1344 12484 34768 12518
rect 4174 12402 4226 12414
rect 4174 12338 4226 12350
rect 5406 12402 5458 12414
rect 5406 12338 5458 12350
rect 5518 12402 5570 12414
rect 5518 12338 5570 12350
rect 20638 12402 20690 12414
rect 20962 12350 20974 12402
rect 21026 12350 21038 12402
rect 20638 12338 20690 12350
rect 3726 12290 3778 12302
rect 3154 12238 3166 12290
rect 3218 12238 3230 12290
rect 3726 12226 3778 12238
rect 4958 12290 5010 12302
rect 4958 12226 5010 12238
rect 8654 12290 8706 12302
rect 8654 12226 8706 12238
rect 8990 12290 9042 12302
rect 8990 12226 9042 12238
rect 10670 12290 10722 12302
rect 18162 12238 18174 12290
rect 18226 12238 18238 12290
rect 22082 12238 22094 12290
rect 22146 12238 22158 12290
rect 10670 12226 10722 12238
rect 2830 12178 2882 12190
rect 4510 12178 4562 12190
rect 4162 12126 4174 12178
rect 4226 12126 4238 12178
rect 2830 12114 2882 12126
rect 4510 12114 4562 12126
rect 4622 12178 4674 12190
rect 4622 12114 4674 12126
rect 5294 12178 5346 12190
rect 6974 12178 7026 12190
rect 10222 12178 10274 12190
rect 5842 12126 5854 12178
rect 5906 12126 5918 12178
rect 6514 12126 6526 12178
rect 6578 12126 6590 12178
rect 7858 12126 7870 12178
rect 7922 12126 7934 12178
rect 5294 12114 5346 12126
rect 6974 12114 7026 12126
rect 10222 12114 10274 12126
rect 10782 12178 10834 12190
rect 26014 12178 26066 12190
rect 31838 12178 31890 12190
rect 12674 12126 12686 12178
rect 12738 12126 12750 12178
rect 17490 12126 17502 12178
rect 17554 12126 17566 12178
rect 21410 12126 21422 12178
rect 21474 12126 21486 12178
rect 26562 12126 26574 12178
rect 26626 12126 26638 12178
rect 31378 12126 31390 12178
rect 31442 12126 31454 12178
rect 10782 12114 10834 12126
rect 26014 12114 26066 12126
rect 31838 12114 31890 12126
rect 10446 12066 10498 12078
rect 24222 12066 24274 12078
rect 3826 12014 3838 12066
rect 3890 12014 3902 12066
rect 8194 12014 8206 12066
rect 8258 12014 8270 12066
rect 13570 12014 13582 12066
rect 13634 12014 13646 12066
rect 20290 12014 20302 12066
rect 20354 12014 20366 12066
rect 26674 12014 26686 12066
rect 26738 12014 26750 12066
rect 10446 12002 10498 12014
rect 24222 12002 24274 12014
rect 3502 11954 3554 11966
rect 3502 11890 3554 11902
rect 31614 11954 31666 11966
rect 31614 11890 31666 11902
rect 31950 11954 32002 11966
rect 31950 11890 32002 11902
rect 1344 11786 34608 11820
rect 1344 11734 5372 11786
rect 5424 11734 5476 11786
rect 5528 11734 5580 11786
rect 5632 11734 13688 11786
rect 13740 11734 13792 11786
rect 13844 11734 13896 11786
rect 13948 11734 22004 11786
rect 22056 11734 22108 11786
rect 22160 11734 22212 11786
rect 22264 11734 30320 11786
rect 30372 11734 30424 11786
rect 30476 11734 30528 11786
rect 30580 11734 34608 11786
rect 1344 11700 34608 11734
rect 6862 11618 6914 11630
rect 6862 11554 6914 11566
rect 8542 11618 8594 11630
rect 17614 11618 17666 11630
rect 20414 11618 20466 11630
rect 17266 11566 17278 11618
rect 17330 11566 17342 11618
rect 18722 11566 18734 11618
rect 18786 11615 18798 11618
rect 18946 11615 18958 11618
rect 18786 11569 18958 11615
rect 18786 11566 18798 11569
rect 18946 11566 18958 11569
rect 19010 11566 19022 11618
rect 8542 11554 8594 11566
rect 17614 11554 17666 11566
rect 20414 11554 20466 11566
rect 22878 11618 22930 11630
rect 22878 11554 22930 11566
rect 2382 11506 2434 11518
rect 2382 11442 2434 11454
rect 3054 11506 3106 11518
rect 3054 11442 3106 11454
rect 4286 11506 4338 11518
rect 4286 11442 4338 11454
rect 6414 11506 6466 11518
rect 6414 11442 6466 11454
rect 10670 11506 10722 11518
rect 18734 11506 18786 11518
rect 11330 11454 11342 11506
rect 11394 11454 11406 11506
rect 14242 11454 14254 11506
rect 14306 11454 14318 11506
rect 16370 11454 16382 11506
rect 16434 11454 16446 11506
rect 10670 11442 10722 11454
rect 18734 11442 18786 11454
rect 19070 11506 19122 11518
rect 19070 11442 19122 11454
rect 20526 11506 20578 11518
rect 20526 11442 20578 11454
rect 21534 11506 21586 11518
rect 22418 11454 22430 11506
rect 22482 11454 22494 11506
rect 27346 11454 27358 11506
rect 27410 11454 27422 11506
rect 31266 11454 31278 11506
rect 31330 11454 31342 11506
rect 33394 11454 33406 11506
rect 33458 11454 33470 11506
rect 21534 11442 21586 11454
rect 2158 11394 2210 11406
rect 2158 11330 2210 11342
rect 3278 11394 3330 11406
rect 3278 11330 3330 11342
rect 3502 11394 3554 11406
rect 3502 11330 3554 11342
rect 3614 11394 3666 11406
rect 3614 11330 3666 11342
rect 4174 11394 4226 11406
rect 5518 11394 5570 11406
rect 4610 11342 4622 11394
rect 4674 11342 4686 11394
rect 4834 11342 4846 11394
rect 4898 11342 4910 11394
rect 4174 11330 4226 11342
rect 5518 11330 5570 11342
rect 5966 11394 6018 11406
rect 5966 11330 6018 11342
rect 6078 11394 6130 11406
rect 6078 11330 6130 11342
rect 6302 11394 6354 11406
rect 6302 11330 6354 11342
rect 6526 11394 6578 11406
rect 6526 11330 6578 11342
rect 7086 11394 7138 11406
rect 7086 11330 7138 11342
rect 7534 11394 7586 11406
rect 7534 11330 7586 11342
rect 8766 11394 8818 11406
rect 8766 11330 8818 11342
rect 8878 11394 8930 11406
rect 8878 11330 8930 11342
rect 9886 11394 9938 11406
rect 9886 11330 9938 11342
rect 10446 11394 10498 11406
rect 10446 11330 10498 11342
rect 10894 11394 10946 11406
rect 17838 11394 17890 11406
rect 19630 11394 19682 11406
rect 13458 11342 13470 11394
rect 13522 11342 13534 11394
rect 19394 11342 19406 11394
rect 19458 11342 19470 11394
rect 10894 11330 10946 11342
rect 17838 11330 17890 11342
rect 19630 11330 19682 11342
rect 19854 11394 19906 11406
rect 22990 11394 23042 11406
rect 29822 11394 29874 11406
rect 20066 11342 20078 11394
rect 20130 11342 20142 11394
rect 21970 11342 21982 11394
rect 22034 11342 22046 11394
rect 24434 11342 24446 11394
rect 24498 11342 24510 11394
rect 30258 11342 30270 11394
rect 30322 11342 30334 11394
rect 34066 11342 34078 11394
rect 34130 11342 34142 11394
rect 19854 11330 19906 11342
rect 22990 11330 23042 11342
rect 29822 11330 29874 11342
rect 7422 11282 7474 11294
rect 7422 11218 7474 11230
rect 8430 11282 8482 11294
rect 8430 11218 8482 11230
rect 9326 11282 9378 11294
rect 9326 11218 9378 11230
rect 10222 11282 10274 11294
rect 10222 11218 10274 11230
rect 11118 11282 11170 11294
rect 11118 11218 11170 11230
rect 16718 11282 16770 11294
rect 25218 11230 25230 11282
rect 25282 11230 25294 11282
rect 16718 11218 16770 11230
rect 2270 11170 2322 11182
rect 2270 11106 2322 11118
rect 2494 11170 2546 11182
rect 2494 11106 2546 11118
rect 2606 11170 2658 11182
rect 2606 11106 2658 11118
rect 3726 11170 3778 11182
rect 3726 11106 3778 11118
rect 4398 11170 4450 11182
rect 4398 11106 4450 11118
rect 7310 11170 7362 11182
rect 7310 11106 7362 11118
rect 11342 11170 11394 11182
rect 11342 11106 11394 11118
rect 12910 11170 12962 11182
rect 12910 11106 12962 11118
rect 16830 11170 16882 11182
rect 16830 11106 16882 11118
rect 19742 11170 19794 11182
rect 19742 11106 19794 11118
rect 29150 11170 29202 11182
rect 29150 11106 29202 11118
rect 29262 11170 29314 11182
rect 29262 11106 29314 11118
rect 29374 11170 29426 11182
rect 30034 11118 30046 11170
rect 30098 11118 30110 11170
rect 29374 11106 29426 11118
rect 1344 11002 34768 11036
rect 1344 10950 9530 11002
rect 9582 10950 9634 11002
rect 9686 10950 9738 11002
rect 9790 10950 17846 11002
rect 17898 10950 17950 11002
rect 18002 10950 18054 11002
rect 18106 10950 26162 11002
rect 26214 10950 26266 11002
rect 26318 10950 26370 11002
rect 26422 10950 34478 11002
rect 34530 10950 34582 11002
rect 34634 10950 34686 11002
rect 34738 10950 34768 11002
rect 1344 10916 34768 10950
rect 3726 10834 3778 10846
rect 3726 10770 3778 10782
rect 4734 10834 4786 10846
rect 4734 10770 4786 10782
rect 4958 10834 5010 10846
rect 7646 10834 7698 10846
rect 7298 10782 7310 10834
rect 7362 10782 7374 10834
rect 4958 10770 5010 10782
rect 7646 10770 7698 10782
rect 10334 10834 10386 10846
rect 10334 10770 10386 10782
rect 10894 10834 10946 10846
rect 10894 10770 10946 10782
rect 16942 10834 16994 10846
rect 16942 10770 16994 10782
rect 17390 10834 17442 10846
rect 17390 10770 17442 10782
rect 22542 10834 22594 10846
rect 22542 10770 22594 10782
rect 25790 10834 25842 10846
rect 31378 10782 31390 10834
rect 31442 10782 31454 10834
rect 25790 10770 25842 10782
rect 3278 10722 3330 10734
rect 3278 10658 3330 10670
rect 3838 10722 3890 10734
rect 3838 10658 3890 10670
rect 6862 10722 6914 10734
rect 6862 10658 6914 10670
rect 8990 10722 9042 10734
rect 8990 10658 9042 10670
rect 10446 10722 10498 10734
rect 22094 10722 22146 10734
rect 13010 10670 13022 10722
rect 13074 10670 13086 10722
rect 10446 10658 10498 10670
rect 22094 10658 22146 10670
rect 26014 10722 26066 10734
rect 26014 10658 26066 10670
rect 31838 10722 31890 10734
rect 31838 10658 31890 10670
rect 2718 10610 2770 10622
rect 5070 10610 5122 10622
rect 3042 10558 3054 10610
rect 3106 10558 3118 10610
rect 2718 10546 2770 10558
rect 5070 10546 5122 10558
rect 6750 10610 6802 10622
rect 6750 10546 6802 10558
rect 7086 10610 7138 10622
rect 8878 10610 8930 10622
rect 8418 10558 8430 10610
rect 8482 10558 8494 10610
rect 7086 10546 7138 10558
rect 8878 10546 8930 10558
rect 9438 10610 9490 10622
rect 9438 10546 9490 10558
rect 9886 10610 9938 10622
rect 9886 10546 9938 10558
rect 9998 10610 10050 10622
rect 9998 10546 10050 10558
rect 10782 10610 10834 10622
rect 10782 10546 10834 10558
rect 11006 10610 11058 10622
rect 11006 10546 11058 10558
rect 11230 10610 11282 10622
rect 30382 10610 30434 10622
rect 12338 10558 12350 10610
rect 12402 10558 12414 10610
rect 18498 10558 18510 10610
rect 18562 10558 18574 10610
rect 21746 10558 21758 10610
rect 21810 10558 21822 10610
rect 27122 10558 27134 10610
rect 27186 10558 27198 10610
rect 11230 10546 11282 10558
rect 30382 10546 30434 10558
rect 30494 10610 30546 10622
rect 30494 10546 30546 10558
rect 30830 10610 30882 10622
rect 30830 10546 30882 10558
rect 30942 10610 30994 10622
rect 32162 10558 32174 10610
rect 32226 10558 32238 10610
rect 30942 10546 30994 10558
rect 2942 10498 2994 10510
rect 2942 10434 2994 10446
rect 10222 10498 10274 10510
rect 15138 10446 15150 10498
rect 15202 10446 15214 10498
rect 17826 10446 17838 10498
rect 17890 10446 17902 10498
rect 19170 10446 19182 10498
rect 19234 10446 19246 10498
rect 21298 10446 21310 10498
rect 21362 10446 21374 10498
rect 25666 10446 25678 10498
rect 25730 10446 25742 10498
rect 27794 10446 27806 10498
rect 27858 10446 27870 10498
rect 29922 10446 29934 10498
rect 29986 10446 29998 10498
rect 10222 10434 10274 10446
rect 3614 10386 3666 10398
rect 3614 10322 3666 10334
rect 8654 10386 8706 10398
rect 8654 10322 8706 10334
rect 21758 10386 21810 10398
rect 21758 10322 21810 10334
rect 32174 10386 32226 10398
rect 32174 10322 32226 10334
rect 1344 10218 34608 10252
rect 1344 10166 5372 10218
rect 5424 10166 5476 10218
rect 5528 10166 5580 10218
rect 5632 10166 13688 10218
rect 13740 10166 13792 10218
rect 13844 10166 13896 10218
rect 13948 10166 22004 10218
rect 22056 10166 22108 10218
rect 22160 10166 22212 10218
rect 22264 10166 30320 10218
rect 30372 10166 30424 10218
rect 30476 10166 30528 10218
rect 30580 10166 34608 10218
rect 1344 10132 34608 10166
rect 2270 10050 2322 10062
rect 2270 9986 2322 9998
rect 7982 10050 8034 10062
rect 7982 9986 8034 9998
rect 9214 10050 9266 10062
rect 9214 9986 9266 9998
rect 21310 10050 21362 10062
rect 21310 9986 21362 9998
rect 3166 9938 3218 9950
rect 3166 9874 3218 9886
rect 3614 9938 3666 9950
rect 3614 9874 3666 9886
rect 6078 9938 6130 9950
rect 6078 9874 6130 9886
rect 8878 9938 8930 9950
rect 12014 9938 12066 9950
rect 21422 9938 21474 9950
rect 10546 9886 10558 9938
rect 10610 9886 10622 9938
rect 12450 9886 12462 9938
rect 12514 9886 12526 9938
rect 15810 9886 15822 9938
rect 15874 9886 15886 9938
rect 8878 9874 8930 9886
rect 12014 9874 12066 9886
rect 21422 9874 21474 9886
rect 30830 9938 30882 9950
rect 31266 9886 31278 9938
rect 31330 9886 31342 9938
rect 30830 9874 30882 9886
rect 2718 9826 2770 9838
rect 2718 9762 2770 9774
rect 2942 9826 2994 9838
rect 5630 9826 5682 9838
rect 4050 9774 4062 9826
rect 4114 9774 4126 9826
rect 2942 9762 2994 9774
rect 5630 9762 5682 9774
rect 5966 9826 6018 9838
rect 11454 9826 11506 9838
rect 9538 9774 9550 9826
rect 9602 9774 9614 9826
rect 5966 9762 6018 9774
rect 11454 9762 11506 9774
rect 11566 9826 11618 9838
rect 11566 9762 11618 9774
rect 12910 9826 12962 9838
rect 12910 9762 12962 9774
rect 13694 9826 13746 9838
rect 13694 9762 13746 9774
rect 15710 9826 15762 9838
rect 18174 9826 18226 9838
rect 20638 9826 20690 9838
rect 17826 9774 17838 9826
rect 17890 9774 17902 9826
rect 20066 9774 20078 9826
rect 20130 9774 20142 9826
rect 15710 9762 15762 9774
rect 18174 9762 18226 9774
rect 20638 9762 20690 9774
rect 22094 9826 22146 9838
rect 29262 9826 29314 9838
rect 27234 9774 27246 9826
rect 27298 9774 27310 9826
rect 22094 9762 22146 9774
rect 29262 9762 29314 9774
rect 29710 9826 29762 9838
rect 29710 9762 29762 9774
rect 30382 9826 30434 9838
rect 30382 9762 30434 9774
rect 30942 9826 30994 9838
rect 34066 9774 34078 9826
rect 34130 9774 34142 9826
rect 30942 9762 30994 9774
rect 6190 9714 6242 9726
rect 6190 9650 6242 9662
rect 7982 9714 8034 9726
rect 8766 9714 8818 9726
rect 9998 9714 10050 9726
rect 7982 9650 8034 9662
rect 8094 9658 8146 9670
rect 3502 9602 3554 9614
rect 3502 9538 3554 9550
rect 3726 9602 3778 9614
rect 8978 9662 8990 9714
rect 9042 9662 9054 9714
rect 8766 9650 8818 9662
rect 9998 9650 10050 9662
rect 10334 9714 10386 9726
rect 10334 9650 10386 9662
rect 10670 9714 10722 9726
rect 11230 9714 11282 9726
rect 19630 9714 19682 9726
rect 10882 9662 10894 9714
rect 10946 9662 10958 9714
rect 14130 9662 14142 9714
rect 14194 9662 14206 9714
rect 17714 9662 17726 9714
rect 17778 9662 17790 9714
rect 18610 9662 18622 9714
rect 18674 9662 18686 9714
rect 18946 9662 18958 9714
rect 19010 9662 19022 9714
rect 10670 9650 10722 9662
rect 11230 9650 11282 9662
rect 19630 9650 19682 9662
rect 21534 9714 21586 9726
rect 29374 9714 29426 9726
rect 24434 9662 24446 9714
rect 24498 9662 24510 9714
rect 21534 9650 21586 9662
rect 29374 9650 29426 9662
rect 30606 9714 30658 9726
rect 33394 9662 33406 9714
rect 33458 9662 33470 9714
rect 30606 9650 30658 9662
rect 8094 9594 8146 9606
rect 10110 9602 10162 9614
rect 3726 9538 3778 9550
rect 10110 9538 10162 9550
rect 13582 9602 13634 9614
rect 28142 9602 28194 9614
rect 29486 9602 29538 9614
rect 18274 9550 18286 9602
rect 18338 9550 18350 9602
rect 28466 9550 28478 9602
rect 28530 9550 28542 9602
rect 13582 9538 13634 9550
rect 28142 9538 28194 9550
rect 29486 9538 29538 9550
rect 1344 9434 34768 9468
rect 1344 9382 9530 9434
rect 9582 9382 9634 9434
rect 9686 9382 9738 9434
rect 9790 9382 17846 9434
rect 17898 9382 17950 9434
rect 18002 9382 18054 9434
rect 18106 9382 26162 9434
rect 26214 9382 26266 9434
rect 26318 9382 26370 9434
rect 26422 9382 34478 9434
rect 34530 9382 34582 9434
rect 34634 9382 34686 9434
rect 34738 9382 34768 9434
rect 1344 9348 34768 9382
rect 2830 9266 2882 9278
rect 2830 9202 2882 9214
rect 3950 9266 4002 9278
rect 3950 9202 4002 9214
rect 4622 9266 4674 9278
rect 4622 9202 4674 9214
rect 5294 9266 5346 9278
rect 5294 9202 5346 9214
rect 5406 9266 5458 9278
rect 5406 9202 5458 9214
rect 7870 9266 7922 9278
rect 24670 9266 24722 9278
rect 26574 9266 26626 9278
rect 10658 9214 10670 9266
rect 10722 9214 10734 9266
rect 23986 9214 23998 9266
rect 24050 9214 24062 9266
rect 26226 9214 26238 9266
rect 26290 9214 26302 9266
rect 7870 9202 7922 9214
rect 24670 9202 24722 9214
rect 26574 9202 26626 9214
rect 33182 9266 33234 9278
rect 33182 9202 33234 9214
rect 4398 9154 4450 9166
rect 4398 9090 4450 9102
rect 5518 9154 5570 9166
rect 5518 9090 5570 9102
rect 6526 9154 6578 9166
rect 6526 9090 6578 9102
rect 9550 9154 9602 9166
rect 9550 9090 9602 9102
rect 9774 9154 9826 9166
rect 14814 9154 14866 9166
rect 12226 9102 12238 9154
rect 12290 9102 12302 9154
rect 18162 9102 18174 9154
rect 18226 9102 18238 9154
rect 18946 9102 18958 9154
rect 19010 9102 19022 9154
rect 21746 9102 21758 9154
rect 21810 9102 21822 9154
rect 31826 9102 31838 9154
rect 31890 9102 31902 9154
rect 9774 9090 9826 9102
rect 14814 9090 14866 9102
rect 3166 9042 3218 9054
rect 3166 8978 3218 8990
rect 3502 9042 3554 9054
rect 4286 9042 4338 9054
rect 6414 9042 6466 9054
rect 3714 8990 3726 9042
rect 3778 8990 3790 9042
rect 5170 8990 5182 9042
rect 5234 8990 5246 9042
rect 3502 8978 3554 8990
rect 4286 8978 4338 8990
rect 6414 8978 6466 8990
rect 6638 9042 6690 9054
rect 6638 8978 6690 8990
rect 7086 9042 7138 9054
rect 7086 8978 7138 8990
rect 7646 9042 7698 9054
rect 7646 8978 7698 8990
rect 7758 9042 7810 9054
rect 7758 8978 7810 8990
rect 8318 9042 8370 9054
rect 11902 9042 11954 9054
rect 15710 9042 15762 9054
rect 33294 9042 33346 9054
rect 9986 8990 9998 9042
rect 10050 8990 10062 9042
rect 10210 8990 10222 9042
rect 10274 8990 10286 9042
rect 10882 8990 10894 9042
rect 10946 8990 10958 9042
rect 13234 8990 13246 9042
rect 13298 8990 13310 9042
rect 13794 8990 13806 9042
rect 13858 8990 13870 9042
rect 17602 8990 17614 9042
rect 17666 8990 17678 9042
rect 19058 8990 19070 9042
rect 19122 8990 19134 9042
rect 20962 8990 20974 9042
rect 21026 8990 21038 9042
rect 25554 8990 25566 9042
rect 25618 8990 25630 9042
rect 27234 8990 27246 9042
rect 27298 8990 27310 9042
rect 33058 8990 33070 9042
rect 33122 8990 33134 9042
rect 8318 8978 8370 8990
rect 11902 8978 11954 8990
rect 15710 8978 15762 8990
rect 33294 8978 33346 8990
rect 16046 8930 16098 8942
rect 2370 8878 2382 8930
rect 2434 8878 2446 8930
rect 10322 8878 10334 8930
rect 10386 8878 10398 8930
rect 16046 8866 16098 8878
rect 16158 8930 16210 8942
rect 25342 8930 25394 8942
rect 17714 8878 17726 8930
rect 17778 8878 17790 8930
rect 16158 8866 16210 8878
rect 25342 8866 25394 8878
rect 4846 8818 4898 8830
rect 11678 8818 11730 8830
rect 3714 8766 3726 8818
rect 3778 8766 3790 8818
rect 11330 8766 11342 8818
rect 11394 8766 11406 8818
rect 4846 8754 4898 8766
rect 11678 8754 11730 8766
rect 25230 8818 25282 8830
rect 25230 8754 25282 8766
rect 33518 8818 33570 8830
rect 33518 8754 33570 8766
rect 1344 8650 34608 8684
rect 1344 8598 5372 8650
rect 5424 8598 5476 8650
rect 5528 8598 5580 8650
rect 5632 8598 13688 8650
rect 13740 8598 13792 8650
rect 13844 8598 13896 8650
rect 13948 8598 22004 8650
rect 22056 8598 22108 8650
rect 22160 8598 22212 8650
rect 22264 8598 30320 8650
rect 30372 8598 30424 8650
rect 30476 8598 30528 8650
rect 30580 8598 34608 8650
rect 1344 8564 34608 8598
rect 29934 8482 29986 8494
rect 29934 8418 29986 8430
rect 2718 8370 2770 8382
rect 5854 8370 5906 8382
rect 21422 8370 21474 8382
rect 3826 8318 3838 8370
rect 3890 8318 3902 8370
rect 9202 8318 9214 8370
rect 9266 8318 9278 8370
rect 13346 8318 13358 8370
rect 13410 8318 13422 8370
rect 17938 8318 17950 8370
rect 18002 8318 18014 8370
rect 19058 8318 19070 8370
rect 19122 8318 19134 8370
rect 2718 8306 2770 8318
rect 5854 8306 5906 8318
rect 21422 8306 21474 8318
rect 22318 8370 22370 8382
rect 30606 8370 30658 8382
rect 23762 8318 23774 8370
rect 23826 8318 23838 8370
rect 25890 8318 25902 8370
rect 25954 8318 25966 8370
rect 28130 8318 28142 8370
rect 28194 8318 28206 8370
rect 34178 8318 34190 8370
rect 34242 8318 34254 8370
rect 22318 8306 22370 8318
rect 30606 8306 30658 8318
rect 3166 8258 3218 8270
rect 3166 8194 3218 8206
rect 3390 8258 3442 8270
rect 3390 8194 3442 8206
rect 3614 8258 3666 8270
rect 3614 8194 3666 8206
rect 5630 8258 5682 8270
rect 5630 8194 5682 8206
rect 6078 8258 6130 8270
rect 6974 8258 7026 8270
rect 6514 8206 6526 8258
rect 6578 8206 6590 8258
rect 6078 8194 6130 8206
rect 6974 8194 7026 8206
rect 9886 8258 9938 8270
rect 9886 8194 9938 8206
rect 12126 8258 12178 8270
rect 22094 8258 22146 8270
rect 26910 8258 26962 8270
rect 13458 8206 13470 8258
rect 13522 8206 13534 8258
rect 15362 8206 15374 8258
rect 15426 8206 15438 8258
rect 18274 8206 18286 8258
rect 18338 8206 18350 8258
rect 18946 8206 18958 8258
rect 19010 8206 19022 8258
rect 23090 8206 23102 8258
rect 23154 8206 23166 8258
rect 12126 8194 12178 8206
rect 22094 8194 22146 8206
rect 26910 8194 26962 8206
rect 27694 8258 27746 8270
rect 27694 8194 27746 8206
rect 29486 8258 29538 8270
rect 29486 8194 29538 8206
rect 29710 8258 29762 8270
rect 30494 8258 30546 8270
rect 30146 8206 30158 8258
rect 30210 8206 30222 8258
rect 31378 8206 31390 8258
rect 31442 8206 31454 8258
rect 29710 8194 29762 8206
rect 30494 8194 30546 8206
rect 2606 8146 2658 8158
rect 2606 8082 2658 8094
rect 2830 8146 2882 8158
rect 2830 8082 2882 8094
rect 3838 8146 3890 8158
rect 3838 8082 3890 8094
rect 4846 8146 4898 8158
rect 7198 8146 7250 8158
rect 6290 8094 6302 8146
rect 6354 8094 6366 8146
rect 4846 8082 4898 8094
rect 7198 8082 7250 8094
rect 7534 8146 7586 8158
rect 7534 8082 7586 8094
rect 8654 8146 8706 8158
rect 8654 8082 8706 8094
rect 8766 8146 8818 8158
rect 9550 8146 9602 8158
rect 8866 8094 8878 8146
rect 8930 8094 8942 8146
rect 8766 8082 8818 8094
rect 9550 8082 9602 8094
rect 10110 8146 10162 8158
rect 10110 8082 10162 8094
rect 10446 8146 10498 8158
rect 10446 8082 10498 8094
rect 10782 8146 10834 8158
rect 10782 8082 10834 8094
rect 11454 8146 11506 8158
rect 11454 8082 11506 8094
rect 12462 8146 12514 8158
rect 12462 8082 12514 8094
rect 12910 8146 12962 8158
rect 28030 8146 28082 8158
rect 14914 8094 14926 8146
rect 14978 8094 14990 8146
rect 16146 8094 16158 8146
rect 16210 8094 16222 8146
rect 12910 8082 12962 8094
rect 28030 8082 28082 8094
rect 29374 8146 29426 8158
rect 32050 8094 32062 8146
rect 32114 8094 32126 8146
rect 29374 8082 29426 8094
rect 4062 8034 4114 8046
rect 4062 7970 4114 7982
rect 4510 8034 4562 8046
rect 4510 7970 4562 7982
rect 5518 8034 5570 8046
rect 5518 7970 5570 7982
rect 7086 8034 7138 8046
rect 7086 7970 7138 7982
rect 7310 8034 7362 8046
rect 7310 7970 7362 7982
rect 8430 8034 8482 8046
rect 8430 7970 8482 7982
rect 9886 8034 9938 8046
rect 9886 7970 9938 7982
rect 11118 8034 11170 8046
rect 12350 8034 12402 8046
rect 11778 7982 11790 8034
rect 11842 7982 11854 8034
rect 11118 7970 11170 7982
rect 12350 7970 12402 7982
rect 12686 8034 12738 8046
rect 12686 7970 12738 7982
rect 17166 8034 17218 8046
rect 26238 8034 26290 8046
rect 28254 8034 28306 8046
rect 21746 7982 21758 8034
rect 21810 7982 21822 8034
rect 26562 7982 26574 8034
rect 26626 7982 26638 8034
rect 27234 7982 27246 8034
rect 27298 7982 27310 8034
rect 17166 7970 17218 7982
rect 26238 7970 26290 7982
rect 28254 7970 28306 7982
rect 1344 7866 34768 7900
rect 1344 7814 9530 7866
rect 9582 7814 9634 7866
rect 9686 7814 9738 7866
rect 9790 7814 17846 7866
rect 17898 7814 17950 7866
rect 18002 7814 18054 7866
rect 18106 7814 26162 7866
rect 26214 7814 26266 7866
rect 26318 7814 26370 7866
rect 26422 7814 34478 7866
rect 34530 7814 34582 7866
rect 34634 7814 34686 7866
rect 34738 7814 34768 7866
rect 1344 7780 34768 7814
rect 2494 7698 2546 7710
rect 2494 7634 2546 7646
rect 2942 7698 2994 7710
rect 6750 7698 6802 7710
rect 27582 7698 27634 7710
rect 5170 7646 5182 7698
rect 5234 7646 5246 7698
rect 7634 7646 7646 7698
rect 7698 7646 7710 7698
rect 2942 7634 2994 7646
rect 6750 7634 6802 7646
rect 9774 7642 9826 7654
rect 4510 7586 4562 7598
rect 9438 7586 9490 7598
rect 8866 7534 8878 7586
rect 8930 7534 8942 7586
rect 4510 7522 4562 7534
rect 9438 7522 9490 7534
rect 9662 7586 9714 7598
rect 27582 7634 27634 7646
rect 28142 7698 28194 7710
rect 32062 7698 32114 7710
rect 30706 7646 30718 7698
rect 30770 7646 30782 7698
rect 28142 7634 28194 7646
rect 32062 7634 32114 7646
rect 9774 7578 9826 7590
rect 16270 7586 16322 7598
rect 23326 7586 23378 7598
rect 9662 7522 9714 7534
rect 22418 7534 22430 7586
rect 22482 7534 22494 7586
rect 16270 7522 16322 7534
rect 23326 7522 23378 7534
rect 23550 7586 23602 7598
rect 23550 7522 23602 7534
rect 25902 7586 25954 7598
rect 25902 7522 25954 7534
rect 28366 7586 28418 7598
rect 28366 7522 28418 7534
rect 29486 7586 29538 7598
rect 29486 7522 29538 7534
rect 29710 7586 29762 7598
rect 33182 7586 33234 7598
rect 32162 7534 32174 7586
rect 32226 7583 32238 7586
rect 32610 7583 32622 7586
rect 32226 7537 32622 7583
rect 32226 7534 32238 7537
rect 32610 7534 32622 7537
rect 32674 7534 32686 7586
rect 29710 7522 29762 7534
rect 33182 7522 33234 7534
rect 2830 7474 2882 7486
rect 2258 7422 2270 7474
rect 2322 7422 2334 7474
rect 2830 7410 2882 7422
rect 3054 7474 3106 7486
rect 3054 7410 3106 7422
rect 3502 7474 3554 7486
rect 3502 7410 3554 7422
rect 3838 7474 3890 7486
rect 3838 7410 3890 7422
rect 3950 7474 4002 7486
rect 3950 7410 4002 7422
rect 4398 7474 4450 7486
rect 4398 7410 4450 7422
rect 4734 7474 4786 7486
rect 5294 7474 5346 7486
rect 5058 7422 5070 7474
rect 5122 7422 5134 7474
rect 4734 7410 4786 7422
rect 5294 7410 5346 7422
rect 5518 7474 5570 7486
rect 5518 7410 5570 7422
rect 5742 7474 5794 7486
rect 5742 7410 5794 7422
rect 6638 7474 6690 7486
rect 6638 7410 6690 7422
rect 6862 7474 6914 7486
rect 6862 7410 6914 7422
rect 7310 7474 7362 7486
rect 11118 7474 11170 7486
rect 7858 7422 7870 7474
rect 7922 7422 7934 7474
rect 8754 7422 8766 7474
rect 8818 7422 8830 7474
rect 10658 7422 10670 7474
rect 10722 7422 10734 7474
rect 7310 7410 7362 7422
rect 11118 7410 11170 7422
rect 13022 7474 13074 7486
rect 15038 7474 15090 7486
rect 18286 7474 18338 7486
rect 21982 7474 22034 7486
rect 13794 7422 13806 7474
rect 13858 7422 13870 7474
rect 16818 7422 16830 7474
rect 16882 7422 16894 7474
rect 18050 7422 18062 7474
rect 18114 7422 18126 7474
rect 18834 7422 18846 7474
rect 18898 7422 18910 7474
rect 13022 7410 13074 7422
rect 15038 7410 15090 7422
rect 18286 7410 18338 7422
rect 21982 7410 22034 7422
rect 22206 7474 22258 7486
rect 22206 7410 22258 7422
rect 22766 7474 22818 7486
rect 22766 7410 22818 7422
rect 22990 7474 23042 7486
rect 22990 7410 23042 7422
rect 25566 7474 25618 7486
rect 25566 7410 25618 7422
rect 26014 7474 26066 7486
rect 26014 7410 26066 7422
rect 26238 7474 26290 7486
rect 26238 7410 26290 7422
rect 27470 7474 27522 7486
rect 29150 7474 29202 7486
rect 27682 7422 27694 7474
rect 27746 7422 27758 7474
rect 27470 7410 27522 7422
rect 29150 7410 29202 7422
rect 29822 7474 29874 7486
rect 31054 7474 31106 7486
rect 30258 7422 30270 7474
rect 30322 7422 30334 7474
rect 29822 7410 29874 7422
rect 31054 7410 31106 7422
rect 31278 7474 31330 7486
rect 31278 7410 31330 7422
rect 31950 7474 32002 7486
rect 32162 7422 32174 7474
rect 32226 7422 32238 7474
rect 33394 7422 33406 7474
rect 33458 7422 33470 7474
rect 31950 7410 32002 7422
rect 14478 7362 14530 7374
rect 8306 7310 8318 7362
rect 8370 7310 8382 7362
rect 12786 7310 12798 7362
rect 12850 7310 12862 7362
rect 14478 7298 14530 7310
rect 17390 7362 17442 7374
rect 23438 7362 23490 7374
rect 19506 7310 19518 7362
rect 19570 7310 19582 7362
rect 21634 7310 21646 7362
rect 21698 7310 21710 7362
rect 17390 7298 17442 7310
rect 23438 7298 23490 7310
rect 4174 7250 4226 7262
rect 27246 7250 27298 7262
rect 26674 7198 26686 7250
rect 26738 7198 26750 7250
rect 4174 7186 4226 7198
rect 27246 7186 27298 7198
rect 28030 7250 28082 7262
rect 28030 7186 28082 7198
rect 31726 7250 31778 7262
rect 31726 7186 31778 7198
rect 33070 7250 33122 7262
rect 33070 7186 33122 7198
rect 1344 7082 34608 7116
rect 1344 7030 5372 7082
rect 5424 7030 5476 7082
rect 5528 7030 5580 7082
rect 5632 7030 13688 7082
rect 13740 7030 13792 7082
rect 13844 7030 13896 7082
rect 13948 7030 22004 7082
rect 22056 7030 22108 7082
rect 22160 7030 22212 7082
rect 22264 7030 30320 7082
rect 30372 7030 30424 7082
rect 30476 7030 30528 7082
rect 30580 7030 34608 7082
rect 1344 6996 34608 7030
rect 3502 6802 3554 6814
rect 3502 6738 3554 6750
rect 4958 6802 5010 6814
rect 4958 6738 5010 6750
rect 5630 6802 5682 6814
rect 5630 6738 5682 6750
rect 9662 6802 9714 6814
rect 9662 6738 9714 6750
rect 10446 6802 10498 6814
rect 18174 6802 18226 6814
rect 29374 6802 29426 6814
rect 30382 6802 30434 6814
rect 14018 6750 14030 6802
rect 14082 6750 14094 6802
rect 19170 6750 19182 6802
rect 19234 6750 19246 6802
rect 22194 6750 22206 6802
rect 22258 6750 22270 6802
rect 23762 6750 23774 6802
rect 23826 6750 23838 6802
rect 29698 6750 29710 6802
rect 29762 6750 29774 6802
rect 33954 6750 33966 6802
rect 34018 6750 34030 6802
rect 10446 6738 10498 6750
rect 18174 6738 18226 6750
rect 29374 6738 29426 6750
rect 30382 6738 30434 6750
rect 5070 6690 5122 6702
rect 9774 6690 9826 6702
rect 6178 6638 6190 6690
rect 6242 6638 6254 6690
rect 8194 6638 8206 6690
rect 8258 6638 8270 6690
rect 8530 6638 8542 6690
rect 8594 6638 8606 6690
rect 5070 6626 5122 6638
rect 9774 6626 9826 6638
rect 10222 6690 10274 6702
rect 11902 6690 11954 6702
rect 11554 6638 11566 6690
rect 11618 6638 11630 6690
rect 10222 6626 10274 6638
rect 11902 6626 11954 6638
rect 12126 6690 12178 6702
rect 12126 6626 12178 6638
rect 12238 6690 12290 6702
rect 19742 6690 19794 6702
rect 14130 6638 14142 6690
rect 14194 6638 14206 6690
rect 14690 6638 14702 6690
rect 14754 6638 14766 6690
rect 15250 6638 15262 6690
rect 15314 6638 15326 6690
rect 12238 6626 12290 6638
rect 19742 6626 19794 6638
rect 22094 6690 22146 6702
rect 27022 6690 27074 6702
rect 22306 6638 22318 6690
rect 22370 6638 22382 6690
rect 23202 6638 23214 6690
rect 23266 6638 23278 6690
rect 26450 6638 26462 6690
rect 26514 6638 26526 6690
rect 22094 6626 22146 6638
rect 27022 6626 27074 6638
rect 27246 6690 27298 6702
rect 29150 6690 29202 6702
rect 27906 6638 27918 6690
rect 27970 6638 27982 6690
rect 27246 6626 27298 6638
rect 29150 6626 29202 6638
rect 30158 6690 30210 6702
rect 30706 6638 30718 6690
rect 30770 6638 30782 6690
rect 31154 6638 31166 6690
rect 31218 6638 31230 6690
rect 30158 6626 30210 6638
rect 5742 6578 5794 6590
rect 12574 6578 12626 6590
rect 22990 6578 23042 6590
rect 26798 6578 26850 6590
rect 6514 6526 6526 6578
rect 6578 6526 6590 6578
rect 9090 6526 9102 6578
rect 9154 6526 9166 6578
rect 11106 6526 11118 6578
rect 11170 6526 11182 6578
rect 11442 6526 11454 6578
rect 11506 6526 11518 6578
rect 13794 6526 13806 6578
rect 13858 6526 13870 6578
rect 16034 6526 16046 6578
rect 16098 6526 16110 6578
rect 24098 6526 24110 6578
rect 24162 6526 24174 6578
rect 24770 6526 24782 6578
rect 24834 6526 24846 6578
rect 31826 6526 31838 6578
rect 31890 6526 31902 6578
rect 5742 6514 5794 6526
rect 12574 6514 12626 6526
rect 22990 6514 23042 6526
rect 26798 6514 26850 6526
rect 3390 6466 3442 6478
rect 3390 6402 3442 6414
rect 4622 6466 4674 6478
rect 4622 6402 4674 6414
rect 4846 6466 4898 6478
rect 7870 6466 7922 6478
rect 9550 6466 9602 6478
rect 6178 6414 6190 6466
rect 6242 6414 6254 6466
rect 7970 6414 7982 6466
rect 8034 6414 8046 6466
rect 4846 6402 4898 6414
rect 7870 6402 7922 6414
rect 9550 6402 9602 6414
rect 18734 6466 18786 6478
rect 18734 6402 18786 6414
rect 27022 6466 27074 6478
rect 27682 6414 27694 6466
rect 27746 6414 27758 6466
rect 27022 6402 27074 6414
rect 1344 6298 34768 6332
rect 1344 6246 9530 6298
rect 9582 6246 9634 6298
rect 9686 6246 9738 6298
rect 9790 6246 17846 6298
rect 17898 6246 17950 6298
rect 18002 6246 18054 6298
rect 18106 6246 26162 6298
rect 26214 6246 26266 6298
rect 26318 6246 26370 6298
rect 26422 6246 34478 6298
rect 34530 6246 34582 6298
rect 34634 6246 34686 6298
rect 34738 6246 34768 6298
rect 1344 6212 34768 6246
rect 7870 6130 7922 6142
rect 3266 6078 3278 6130
rect 3330 6078 3342 6130
rect 7870 6066 7922 6078
rect 7982 6130 8034 6142
rect 11566 6130 11618 6142
rect 17950 6130 18002 6142
rect 9650 6078 9662 6130
rect 9714 6078 9726 6130
rect 13570 6078 13582 6130
rect 13634 6078 13646 6130
rect 7982 6066 8034 6078
rect 11566 6066 11618 6078
rect 17950 6066 18002 6078
rect 27694 6130 27746 6142
rect 27694 6066 27746 6078
rect 5854 6018 5906 6030
rect 8430 6018 8482 6030
rect 11118 6018 11170 6030
rect 17390 6018 17442 6030
rect 4050 5966 4062 6018
rect 4114 5966 4126 6018
rect 6514 5966 6526 6018
rect 6578 5966 6590 6018
rect 8754 5966 8766 6018
rect 8818 5966 8830 6018
rect 12450 5966 12462 6018
rect 12514 5966 12526 6018
rect 12786 5966 12798 6018
rect 12850 5966 12862 6018
rect 13682 5966 13694 6018
rect 13746 5966 13758 6018
rect 14242 5966 14254 6018
rect 14306 5966 14318 6018
rect 5854 5954 5906 5966
rect 8430 5954 8482 5966
rect 11118 5954 11170 5966
rect 17390 5954 17442 5966
rect 20526 6018 20578 6030
rect 20526 5954 20578 5966
rect 20974 6018 21026 6030
rect 20974 5954 21026 5966
rect 21310 6018 21362 6030
rect 21310 5954 21362 5966
rect 22990 6018 23042 6030
rect 22990 5954 23042 5966
rect 24670 6018 24722 6030
rect 24670 5954 24722 5966
rect 25454 6018 25506 6030
rect 25454 5954 25506 5966
rect 28702 6018 28754 6030
rect 28702 5954 28754 5966
rect 28926 6018 28978 6030
rect 28926 5954 28978 5966
rect 29822 6018 29874 6030
rect 29822 5954 29874 5966
rect 30942 6018 30994 6030
rect 30942 5954 30994 5966
rect 33406 6018 33458 6030
rect 33406 5954 33458 5966
rect 2606 5906 2658 5918
rect 3726 5906 3778 5918
rect 3042 5854 3054 5906
rect 3106 5854 3118 5906
rect 2606 5842 2658 5854
rect 3726 5842 3778 5854
rect 4398 5906 4450 5918
rect 5294 5906 5346 5918
rect 8206 5906 8258 5918
rect 9998 5906 10050 5918
rect 4834 5854 4846 5906
rect 4898 5854 4910 5906
rect 6290 5854 6302 5906
rect 6354 5854 6366 5906
rect 7410 5854 7422 5906
rect 7474 5854 7486 5906
rect 7634 5854 7646 5906
rect 7698 5854 7710 5906
rect 8642 5854 8654 5906
rect 8706 5854 8718 5906
rect 4398 5842 4450 5854
rect 5294 5842 5346 5854
rect 8206 5842 8258 5854
rect 9998 5842 10050 5854
rect 10558 5906 10610 5918
rect 10558 5842 10610 5854
rect 11454 5906 11506 5918
rect 19294 5906 19346 5918
rect 21422 5906 21474 5918
rect 13122 5854 13134 5906
rect 13186 5854 13198 5906
rect 14578 5854 14590 5906
rect 14642 5854 14654 5906
rect 15698 5854 15710 5906
rect 15762 5854 15774 5906
rect 16146 5854 16158 5906
rect 16210 5854 16222 5906
rect 18722 5854 18734 5906
rect 18786 5854 18798 5906
rect 20066 5854 20078 5906
rect 20130 5854 20142 5906
rect 11454 5842 11506 5854
rect 19294 5842 19346 5854
rect 21422 5842 21474 5854
rect 21646 5906 21698 5918
rect 21646 5842 21698 5854
rect 21758 5906 21810 5918
rect 21758 5842 21810 5854
rect 22654 5906 22706 5918
rect 25566 5906 25618 5918
rect 24210 5854 24222 5906
rect 24274 5854 24286 5906
rect 25218 5854 25230 5906
rect 25282 5854 25294 5906
rect 22654 5842 22706 5854
rect 25566 5842 25618 5854
rect 26686 5906 26738 5918
rect 26686 5842 26738 5854
rect 27470 5906 27522 5918
rect 30494 5906 30546 5918
rect 30034 5854 30046 5906
rect 30098 5854 30110 5906
rect 27470 5842 27522 5854
rect 30494 5842 30546 5854
rect 31166 5906 31218 5918
rect 31166 5842 31218 5854
rect 31614 5906 31666 5918
rect 31614 5842 31666 5854
rect 31950 5906 32002 5918
rect 31950 5842 32002 5854
rect 32958 5906 33010 5918
rect 32958 5842 33010 5854
rect 33630 5906 33682 5918
rect 33630 5842 33682 5854
rect 10222 5794 10274 5806
rect 2146 5742 2158 5794
rect 2210 5742 2222 5794
rect 6402 5742 6414 5794
rect 6466 5742 6478 5794
rect 8978 5742 8990 5794
rect 9042 5742 9054 5794
rect 10222 5730 10274 5742
rect 11902 5794 11954 5806
rect 19406 5794 19458 5806
rect 16706 5742 16718 5794
rect 16770 5742 16782 5794
rect 11902 5730 11954 5742
rect 19406 5730 19458 5742
rect 19742 5794 19794 5806
rect 19742 5730 19794 5742
rect 19854 5794 19906 5806
rect 27582 5794 27634 5806
rect 22530 5742 22542 5794
rect 22594 5742 22606 5794
rect 24322 5742 24334 5794
rect 24386 5742 24398 5794
rect 26002 5742 26014 5794
rect 26066 5742 26078 5794
rect 19854 5730 19906 5742
rect 27582 5730 27634 5742
rect 31054 5794 31106 5806
rect 31054 5730 31106 5742
rect 31726 5794 31778 5806
rect 31726 5730 31778 5742
rect 33182 5794 33234 5806
rect 33182 5730 33234 5742
rect 11566 5682 11618 5694
rect 11566 5618 11618 5630
rect 26798 5682 26850 5694
rect 26798 5618 26850 5630
rect 27022 5682 27074 5694
rect 27022 5618 27074 5630
rect 27134 5682 27186 5694
rect 27134 5618 27186 5630
rect 29038 5682 29090 5694
rect 29038 5618 29090 5630
rect 32062 5682 32114 5694
rect 32062 5618 32114 5630
rect 1344 5514 34608 5548
rect 1344 5462 5372 5514
rect 5424 5462 5476 5514
rect 5528 5462 5580 5514
rect 5632 5462 13688 5514
rect 13740 5462 13792 5514
rect 13844 5462 13896 5514
rect 13948 5462 22004 5514
rect 22056 5462 22108 5514
rect 22160 5462 22212 5514
rect 22264 5462 30320 5514
rect 30372 5462 30424 5514
rect 30476 5462 30528 5514
rect 30580 5462 34608 5514
rect 1344 5428 34608 5462
rect 4622 5346 4674 5358
rect 3938 5294 3950 5346
rect 4002 5294 4014 5346
rect 4622 5282 4674 5294
rect 21982 5346 22034 5358
rect 21982 5282 22034 5294
rect 27582 5346 27634 5358
rect 27582 5282 27634 5294
rect 29262 5346 29314 5358
rect 29262 5282 29314 5294
rect 3390 5234 3442 5246
rect 2930 5182 2942 5234
rect 2994 5182 3006 5234
rect 3390 5170 3442 5182
rect 11790 5234 11842 5246
rect 19182 5234 19234 5246
rect 12114 5182 12126 5234
rect 12178 5182 12190 5234
rect 11790 5170 11842 5182
rect 19182 5170 19234 5182
rect 21646 5234 21698 5246
rect 27806 5234 27858 5246
rect 24098 5182 24110 5234
rect 24162 5182 24174 5234
rect 32050 5182 32062 5234
rect 32114 5182 32126 5234
rect 34178 5182 34190 5234
rect 34242 5182 34254 5234
rect 21646 5170 21698 5182
rect 27806 5170 27858 5182
rect 2494 5122 2546 5134
rect 2494 5058 2546 5070
rect 3614 5122 3666 5134
rect 9326 5122 9378 5134
rect 4274 5070 4286 5122
rect 4338 5070 4350 5122
rect 4834 5070 4846 5122
rect 4898 5070 4910 5122
rect 5954 5070 5966 5122
rect 6018 5070 6030 5122
rect 7410 5070 7422 5122
rect 7474 5070 7486 5122
rect 8082 5070 8094 5122
rect 8146 5070 8158 5122
rect 8866 5070 8878 5122
rect 8930 5070 8942 5122
rect 3614 5058 3666 5070
rect 9326 5058 9378 5070
rect 10110 5122 10162 5134
rect 10110 5058 10162 5070
rect 10894 5122 10946 5134
rect 10894 5058 10946 5070
rect 11230 5122 11282 5134
rect 13470 5122 13522 5134
rect 21870 5122 21922 5134
rect 12674 5070 12686 5122
rect 12738 5070 12750 5122
rect 13906 5070 13918 5122
rect 13970 5070 13982 5122
rect 15922 5070 15934 5122
rect 15986 5070 15998 5122
rect 18162 5070 18174 5122
rect 18226 5070 18238 5122
rect 11230 5058 11282 5070
rect 13470 5058 13522 5070
rect 21870 5058 21922 5070
rect 22766 5122 22818 5134
rect 22766 5058 22818 5070
rect 23326 5122 23378 5134
rect 29486 5122 29538 5134
rect 30382 5122 30434 5134
rect 27010 5070 27022 5122
rect 27074 5070 27086 5122
rect 27346 5070 27358 5122
rect 27410 5070 27422 5122
rect 29698 5070 29710 5122
rect 29762 5070 29774 5122
rect 23326 5058 23378 5070
rect 29486 5058 29538 5070
rect 30382 5058 30434 5070
rect 30494 5122 30546 5134
rect 30494 5058 30546 5070
rect 30718 5122 30770 5134
rect 30718 5058 30770 5070
rect 30942 5122 30994 5134
rect 31266 5070 31278 5122
rect 31330 5070 31342 5122
rect 30942 5058 30994 5070
rect 5070 5010 5122 5022
rect 5070 4946 5122 4958
rect 6190 5010 6242 5022
rect 21534 5010 21586 5022
rect 7298 4958 7310 5010
rect 7362 4958 7374 5010
rect 7858 4958 7870 5010
rect 7922 4958 7934 5010
rect 9874 4958 9886 5010
rect 9938 4958 9950 5010
rect 10546 4958 10558 5010
rect 10610 4958 10622 5010
rect 12450 4958 12462 5010
rect 12514 4958 12526 5010
rect 14018 4958 14030 5010
rect 14082 4958 14094 5010
rect 17714 4958 17726 5010
rect 17778 4958 17790 5010
rect 26226 4958 26238 5010
rect 26290 4958 26302 5010
rect 6190 4946 6242 4958
rect 21534 4946 21586 4958
rect 4286 4898 4338 4910
rect 7646 4898 7698 4910
rect 6290 4846 6302 4898
rect 6354 4846 6366 4898
rect 4286 4834 4338 4846
rect 7646 4834 7698 4846
rect 13582 4898 13634 4910
rect 27470 4898 27522 4910
rect 15362 4846 15374 4898
rect 15426 4846 15438 4898
rect 13582 4834 13634 4846
rect 27470 4834 27522 4846
rect 29598 4898 29650 4910
rect 29598 4834 29650 4846
rect 1344 4730 34768 4764
rect 1344 4678 9530 4730
rect 9582 4678 9634 4730
rect 9686 4678 9738 4730
rect 9790 4678 17846 4730
rect 17898 4678 17950 4730
rect 18002 4678 18054 4730
rect 18106 4678 26162 4730
rect 26214 4678 26266 4730
rect 26318 4678 26370 4730
rect 26422 4678 34478 4730
rect 34530 4678 34582 4730
rect 34634 4678 34686 4730
rect 34738 4678 34768 4730
rect 1344 4644 34768 4678
rect 6862 4562 6914 4574
rect 11118 4562 11170 4574
rect 4722 4510 4734 4562
rect 4786 4510 4798 4562
rect 7634 4510 7646 4562
rect 7698 4510 7710 4562
rect 7970 4510 7982 4562
rect 8034 4510 8046 4562
rect 8978 4510 8990 4562
rect 9042 4510 9054 4562
rect 6862 4498 6914 4510
rect 11118 4498 11170 4510
rect 17278 4562 17330 4574
rect 17278 4498 17330 4510
rect 19070 4562 19122 4574
rect 22754 4510 22766 4562
rect 22818 4510 22830 4562
rect 33058 4510 33070 4562
rect 33122 4510 33134 4562
rect 19070 4498 19122 4510
rect 6974 4450 7026 4462
rect 2482 4398 2494 4450
rect 2546 4398 2558 4450
rect 6402 4398 6414 4450
rect 6466 4398 6478 4450
rect 10770 4398 10782 4450
rect 10834 4398 10846 4450
rect 13346 4398 13358 4450
rect 13410 4398 13422 4450
rect 27906 4398 27918 4450
rect 27970 4398 27982 4450
rect 31154 4398 31166 4450
rect 31218 4398 31230 4450
rect 6974 4386 7026 4398
rect 11230 4338 11282 4350
rect 17614 4338 17666 4350
rect 23102 4338 23154 4350
rect 1810 4286 1822 4338
rect 1874 4286 1886 4338
rect 7410 4286 7422 4338
rect 7474 4286 7486 4338
rect 8194 4286 8206 4338
rect 8258 4286 8270 4338
rect 8754 4286 8766 4338
rect 8818 4286 8830 4338
rect 12114 4286 12126 4338
rect 12178 4286 12190 4338
rect 12562 4286 12574 4338
rect 12626 4286 12638 4338
rect 18050 4286 18062 4338
rect 18114 4286 18126 4338
rect 19506 4286 19518 4338
rect 19570 4286 19582 4338
rect 11230 4274 11282 4286
rect 17614 4274 17666 4286
rect 23102 4274 23154 4286
rect 23774 4338 23826 4350
rect 33406 4338 33458 4350
rect 24210 4286 24222 4338
rect 24274 4286 24286 4338
rect 28690 4286 28702 4338
rect 28754 4286 28766 4338
rect 31938 4286 31950 4338
rect 32002 4286 32014 4338
rect 23774 4274 23826 4286
rect 33406 4274 33458 4286
rect 33630 4338 33682 4350
rect 33630 4274 33682 4286
rect 23326 4226 23378 4238
rect 11778 4174 11790 4226
rect 11842 4174 11854 4226
rect 15474 4174 15486 4226
rect 15538 4174 15550 4226
rect 17714 4174 17726 4226
rect 17778 4174 17790 4226
rect 20290 4174 20302 4226
rect 20354 4174 20366 4226
rect 22418 4174 22430 4226
rect 22482 4174 22494 4226
rect 23326 4162 23378 4174
rect 23662 4226 23714 4238
rect 25778 4174 25790 4226
rect 25842 4174 25854 4226
rect 29026 4174 29038 4226
rect 29090 4174 29102 4226
rect 23662 4162 23714 4174
rect 5854 4114 5906 4126
rect 5854 4050 5906 4062
rect 6862 4114 6914 4126
rect 6862 4050 6914 4062
rect 10222 4114 10274 4126
rect 10222 4050 10274 4062
rect 23998 4114 24050 4126
rect 23998 4050 24050 4062
rect 1344 3946 34608 3980
rect 1344 3894 5372 3946
rect 5424 3894 5476 3946
rect 5528 3894 5580 3946
rect 5632 3894 13688 3946
rect 13740 3894 13792 3946
rect 13844 3894 13896 3946
rect 13948 3894 22004 3946
rect 22056 3894 22108 3946
rect 22160 3894 22212 3946
rect 22264 3894 30320 3946
rect 30372 3894 30424 3946
rect 30476 3894 30528 3946
rect 30580 3894 34608 3946
rect 1344 3860 34608 3894
rect 7086 3778 7138 3790
rect 7086 3714 7138 3726
rect 14142 3778 14194 3790
rect 14142 3714 14194 3726
rect 14478 3778 14530 3790
rect 14478 3714 14530 3726
rect 14926 3778 14978 3790
rect 14926 3714 14978 3726
rect 15262 3778 15314 3790
rect 15262 3714 15314 3726
rect 5742 3666 5794 3678
rect 8430 3666 8482 3678
rect 12350 3666 12402 3678
rect 15486 3666 15538 3678
rect 24558 3666 24610 3678
rect 8082 3614 8094 3666
rect 8146 3614 8158 3666
rect 10210 3614 10222 3666
rect 10274 3614 10286 3666
rect 13570 3614 13582 3666
rect 13634 3614 13646 3666
rect 16930 3614 16942 3666
rect 16994 3614 17006 3666
rect 21522 3614 21534 3666
rect 21586 3614 21598 3666
rect 23650 3614 23662 3666
rect 23714 3614 23726 3666
rect 5742 3602 5794 3614
rect 8430 3602 8482 3614
rect 12350 3602 12402 3614
rect 15486 3602 15538 3614
rect 24558 3602 24610 3614
rect 24670 3666 24722 3678
rect 24670 3602 24722 3614
rect 32958 3666 33010 3678
rect 32958 3602 33010 3614
rect 6078 3554 6130 3566
rect 6078 3490 6130 3502
rect 6750 3554 6802 3566
rect 14366 3554 14418 3566
rect 6962 3502 6974 3554
rect 7026 3502 7038 3554
rect 9538 3502 9550 3554
rect 9602 3502 9614 3554
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 24882 3502 24894 3554
rect 24946 3502 24958 3554
rect 25218 3502 25230 3554
rect 25282 3502 25294 3554
rect 31490 3502 31502 3554
rect 31554 3502 31566 3554
rect 32386 3502 32398 3554
rect 32450 3502 32462 3554
rect 6750 3490 6802 3502
rect 14366 3490 14418 3502
rect 6302 3442 6354 3454
rect 6302 3378 6354 3390
rect 6526 3442 6578 3454
rect 6526 3378 6578 3390
rect 13246 3442 13298 3454
rect 32174 3442 32226 3454
rect 19058 3390 19070 3442
rect 19122 3390 19134 3442
rect 26898 3390 26910 3442
rect 26962 3390 26974 3442
rect 30034 3390 30046 3442
rect 30098 3390 30110 3442
rect 13246 3378 13298 3390
rect 32174 3378 32226 3390
rect 1344 3162 34768 3196
rect 1344 3110 9530 3162
rect 9582 3110 9634 3162
rect 9686 3110 9738 3162
rect 9790 3110 17846 3162
rect 17898 3110 17950 3162
rect 18002 3110 18054 3162
rect 18106 3110 26162 3162
rect 26214 3110 26266 3162
rect 26318 3110 26370 3162
rect 26422 3110 34478 3162
rect 34530 3110 34582 3162
rect 34634 3110 34686 3162
rect 34738 3110 34768 3162
rect 1344 3076 34768 3110
<< via1 >>
rect 5372 32118 5424 32170
rect 5476 32118 5528 32170
rect 5580 32118 5632 32170
rect 13688 32118 13740 32170
rect 13792 32118 13844 32170
rect 13896 32118 13948 32170
rect 22004 32118 22056 32170
rect 22108 32118 22160 32170
rect 22212 32118 22264 32170
rect 30320 32118 30372 32170
rect 30424 32118 30476 32170
rect 30528 32118 30580 32170
rect 9530 31334 9582 31386
rect 9634 31334 9686 31386
rect 9738 31334 9790 31386
rect 17846 31334 17898 31386
rect 17950 31334 18002 31386
rect 18054 31334 18106 31386
rect 26162 31334 26214 31386
rect 26266 31334 26318 31386
rect 26370 31334 26422 31386
rect 34478 31334 34530 31386
rect 34582 31334 34634 31386
rect 34686 31334 34738 31386
rect 5372 30550 5424 30602
rect 5476 30550 5528 30602
rect 5580 30550 5632 30602
rect 13688 30550 13740 30602
rect 13792 30550 13844 30602
rect 13896 30550 13948 30602
rect 22004 30550 22056 30602
rect 22108 30550 22160 30602
rect 22212 30550 22264 30602
rect 30320 30550 30372 30602
rect 30424 30550 30476 30602
rect 30528 30550 30580 30602
rect 9530 29766 9582 29818
rect 9634 29766 9686 29818
rect 9738 29766 9790 29818
rect 17846 29766 17898 29818
rect 17950 29766 18002 29818
rect 18054 29766 18106 29818
rect 26162 29766 26214 29818
rect 26266 29766 26318 29818
rect 26370 29766 26422 29818
rect 34478 29766 34530 29818
rect 34582 29766 34634 29818
rect 34686 29766 34738 29818
rect 5372 28982 5424 29034
rect 5476 28982 5528 29034
rect 5580 28982 5632 29034
rect 13688 28982 13740 29034
rect 13792 28982 13844 29034
rect 13896 28982 13948 29034
rect 22004 28982 22056 29034
rect 22108 28982 22160 29034
rect 22212 28982 22264 29034
rect 30320 28982 30372 29034
rect 30424 28982 30476 29034
rect 30528 28982 30580 29034
rect 11230 28702 11282 28754
rect 8430 28590 8482 28642
rect 9102 28478 9154 28530
rect 9530 28198 9582 28250
rect 9634 28198 9686 28250
rect 9738 28198 9790 28250
rect 17846 28198 17898 28250
rect 17950 28198 18002 28250
rect 18054 28198 18106 28250
rect 26162 28198 26214 28250
rect 26266 28198 26318 28250
rect 26370 28198 26422 28250
rect 34478 28198 34530 28250
rect 34582 28198 34634 28250
rect 34686 28198 34738 28250
rect 20302 28030 20354 28082
rect 5070 27918 5122 27970
rect 4286 27806 4338 27858
rect 4510 27806 4562 27858
rect 4846 27806 4898 27858
rect 5182 27806 5234 27858
rect 10222 27806 10274 27858
rect 19966 27806 20018 27858
rect 20190 27806 20242 27858
rect 20526 27806 20578 27858
rect 3614 27694 3666 27746
rect 11006 27694 11058 27746
rect 13134 27694 13186 27746
rect 5372 27414 5424 27466
rect 5476 27414 5528 27466
rect 5580 27414 5632 27466
rect 13688 27414 13740 27466
rect 13792 27414 13844 27466
rect 13896 27414 13948 27466
rect 22004 27414 22056 27466
rect 22108 27414 22160 27466
rect 22212 27414 22264 27466
rect 30320 27414 30372 27466
rect 30424 27414 30476 27466
rect 30528 27414 30580 27466
rect 5854 27246 5906 27298
rect 4622 27134 4674 27186
rect 4958 27134 5010 27186
rect 10334 27134 10386 27186
rect 12238 27134 12290 27186
rect 17166 27134 17218 27186
rect 20414 27134 20466 27186
rect 1822 27022 1874 27074
rect 5966 27022 6018 27074
rect 6190 27022 6242 27074
rect 6750 27022 6802 27074
rect 7422 27022 7474 27074
rect 12462 27022 12514 27074
rect 14366 27022 14418 27074
rect 17614 27022 17666 27074
rect 23774 27022 23826 27074
rect 24222 27022 24274 27074
rect 2494 26910 2546 26962
rect 5070 26910 5122 26962
rect 6302 26910 6354 26962
rect 6638 26910 6690 26962
rect 6862 26910 6914 26962
rect 8206 26910 8258 26962
rect 12126 26910 12178 26962
rect 12686 26910 12738 26962
rect 15038 26910 15090 26962
rect 18286 26910 18338 26962
rect 24110 26910 24162 26962
rect 23438 26798 23490 26850
rect 9530 26630 9582 26682
rect 9634 26630 9686 26682
rect 9738 26630 9790 26682
rect 17846 26630 17898 26682
rect 17950 26630 18002 26682
rect 18054 26630 18106 26682
rect 26162 26630 26214 26682
rect 26266 26630 26318 26682
rect 26370 26630 26422 26682
rect 34478 26630 34530 26682
rect 34582 26630 34634 26682
rect 34686 26630 34738 26682
rect 9886 26462 9938 26514
rect 16270 26462 16322 26514
rect 18062 26462 18114 26514
rect 18958 26462 19010 26514
rect 25678 26462 25730 26514
rect 7310 26350 7362 26402
rect 16606 26350 16658 26402
rect 19182 26350 19234 26402
rect 20414 26350 20466 26402
rect 25342 26350 25394 26402
rect 1822 26238 1874 26290
rect 7982 26238 8034 26290
rect 11790 26238 11842 26290
rect 12350 26238 12402 26290
rect 15822 26238 15874 26290
rect 16158 26238 16210 26290
rect 16382 26238 16434 26290
rect 17838 26238 17890 26290
rect 18174 26238 18226 26290
rect 18286 26238 18338 26290
rect 18734 26238 18786 26290
rect 18846 26238 18898 26290
rect 19630 26238 19682 26290
rect 25566 26238 25618 26290
rect 25790 26238 25842 26290
rect 2494 26126 2546 26178
rect 4622 26126 4674 26178
rect 5182 26126 5234 26178
rect 9998 26126 10050 26178
rect 12462 26126 12514 26178
rect 12910 26126 12962 26178
rect 15038 26126 15090 26178
rect 22542 26126 22594 26178
rect 5372 25846 5424 25898
rect 5476 25846 5528 25898
rect 5580 25846 5632 25898
rect 13688 25846 13740 25898
rect 13792 25846 13844 25898
rect 13896 25846 13948 25898
rect 22004 25846 22056 25898
rect 22108 25846 22160 25898
rect 22212 25846 22264 25898
rect 30320 25846 30372 25898
rect 30424 25846 30476 25898
rect 30528 25846 30580 25898
rect 2606 25678 2658 25730
rect 2942 25678 2994 25730
rect 3278 25678 3330 25730
rect 18510 25678 18562 25730
rect 18958 25678 19010 25730
rect 19294 25678 19346 25730
rect 4958 25566 5010 25618
rect 9886 25566 9938 25618
rect 13582 25566 13634 25618
rect 14478 25566 14530 25618
rect 15374 25566 15426 25618
rect 19966 25566 20018 25618
rect 22990 25566 23042 25618
rect 2606 25454 2658 25506
rect 3278 25454 3330 25506
rect 4622 25454 4674 25506
rect 7086 25454 7138 25506
rect 12014 25454 12066 25506
rect 12574 25454 12626 25506
rect 13694 25454 13746 25506
rect 14142 25454 14194 25506
rect 14254 25454 14306 25506
rect 14702 25454 14754 25506
rect 15150 25454 15202 25506
rect 15486 25454 15538 25506
rect 15822 25454 15874 25506
rect 18622 25454 18674 25506
rect 20078 25454 20130 25506
rect 25902 25454 25954 25506
rect 26350 25454 26402 25506
rect 3614 25342 3666 25394
rect 4062 25342 4114 25394
rect 7758 25342 7810 25394
rect 12350 25342 12402 25394
rect 14926 25342 14978 25394
rect 16158 25342 16210 25394
rect 16606 25342 16658 25394
rect 19518 25342 19570 25394
rect 19854 25342 19906 25394
rect 25230 25342 25282 25394
rect 26574 25342 26626 25394
rect 26910 25342 26962 25394
rect 27358 25342 27410 25394
rect 27582 25342 27634 25394
rect 12462 25230 12514 25282
rect 13470 25230 13522 25282
rect 16270 25230 16322 25282
rect 16382 25230 16434 25282
rect 20302 25230 20354 25282
rect 26686 25230 26738 25282
rect 27470 25230 27522 25282
rect 28142 25230 28194 25282
rect 9530 25062 9582 25114
rect 9634 25062 9686 25114
rect 9738 25062 9790 25114
rect 17846 25062 17898 25114
rect 17950 25062 18002 25114
rect 18054 25062 18106 25114
rect 26162 25062 26214 25114
rect 26266 25062 26318 25114
rect 26370 25062 26422 25114
rect 34478 25062 34530 25114
rect 34582 25062 34634 25114
rect 34686 25062 34738 25114
rect 4734 24894 4786 24946
rect 6190 24894 6242 24946
rect 8878 24894 8930 24946
rect 11006 24894 11058 24946
rect 11118 24894 11170 24946
rect 11230 24894 11282 24946
rect 12462 24894 12514 24946
rect 15150 24894 15202 24946
rect 15262 24894 15314 24946
rect 17502 24894 17554 24946
rect 18174 24894 18226 24946
rect 18846 24894 18898 24946
rect 24334 24894 24386 24946
rect 4062 24782 4114 24834
rect 5854 24782 5906 24834
rect 6414 24782 6466 24834
rect 11342 24782 11394 24834
rect 12350 24782 12402 24834
rect 12686 24782 12738 24834
rect 13470 24782 13522 24834
rect 14254 24782 14306 24834
rect 15710 24782 15762 24834
rect 24670 24782 24722 24834
rect 28702 24782 28754 24834
rect 4398 24670 4450 24722
rect 5070 24670 5122 24722
rect 5294 24670 5346 24722
rect 5630 24670 5682 24722
rect 11678 24670 11730 24722
rect 12238 24670 12290 24722
rect 12574 24670 12626 24722
rect 13134 24670 13186 24722
rect 14142 24670 14194 24722
rect 14478 24670 14530 24722
rect 14590 24670 14642 24722
rect 15038 24670 15090 24722
rect 17838 24670 17890 24722
rect 18398 24670 18450 24722
rect 19070 24670 19122 24722
rect 20302 24670 20354 24722
rect 22654 24670 22706 24722
rect 23438 24670 23490 24722
rect 29374 24670 29426 24722
rect 8990 24558 9042 24610
rect 13358 24558 13410 24610
rect 20526 24558 20578 24610
rect 22430 24558 22482 24610
rect 26462 24558 26514 24610
rect 15598 24446 15650 24498
rect 5372 24278 5424 24330
rect 5476 24278 5528 24330
rect 5580 24278 5632 24330
rect 13688 24278 13740 24330
rect 13792 24278 13844 24330
rect 13896 24278 13948 24330
rect 22004 24278 22056 24330
rect 22108 24278 22160 24330
rect 22212 24278 22264 24330
rect 30320 24278 30372 24330
rect 30424 24278 30476 24330
rect 30528 24278 30580 24330
rect 12126 24110 12178 24162
rect 13582 24110 13634 24162
rect 18846 24110 18898 24162
rect 9998 23998 10050 24050
rect 11006 23998 11058 24050
rect 14926 23998 14978 24050
rect 19182 23998 19234 24050
rect 19854 23998 19906 24050
rect 20302 23998 20354 24050
rect 22430 23998 22482 24050
rect 28030 23998 28082 24050
rect 7086 23886 7138 23938
rect 10894 23886 10946 23938
rect 11678 23886 11730 23938
rect 13022 23886 13074 23938
rect 13470 23886 13522 23938
rect 14142 23886 14194 23938
rect 17838 23886 17890 23938
rect 22206 23886 22258 23938
rect 22766 23886 22818 23938
rect 23438 23886 23490 23938
rect 24222 23886 24274 23938
rect 24558 23886 24610 23938
rect 25566 23886 25618 23938
rect 27918 23886 27970 23938
rect 28142 23886 28194 23938
rect 5070 23774 5122 23826
rect 7870 23774 7922 23826
rect 11118 23774 11170 23826
rect 11230 23774 11282 23826
rect 12014 23774 12066 23826
rect 13918 23774 13970 23826
rect 17166 23774 17218 23826
rect 19518 23774 19570 23826
rect 19742 23774 19794 23826
rect 27134 23774 27186 23826
rect 29150 23774 29202 23826
rect 29374 23774 29426 23826
rect 4846 23662 4898 23714
rect 4958 23662 5010 23714
rect 12126 23662 12178 23714
rect 13694 23662 13746 23714
rect 18510 23662 18562 23714
rect 19070 23662 19122 23714
rect 24782 23662 24834 23714
rect 26126 23662 26178 23714
rect 27022 23662 27074 23714
rect 27246 23662 27298 23714
rect 27470 23662 27522 23714
rect 28366 23662 28418 23714
rect 29262 23662 29314 23714
rect 29934 23662 29986 23714
rect 9530 23494 9582 23546
rect 9634 23494 9686 23546
rect 9738 23494 9790 23546
rect 17846 23494 17898 23546
rect 17950 23494 18002 23546
rect 18054 23494 18106 23546
rect 26162 23494 26214 23546
rect 26266 23494 26318 23546
rect 26370 23494 26422 23546
rect 34478 23494 34530 23546
rect 34582 23494 34634 23546
rect 34686 23494 34738 23546
rect 5518 23326 5570 23378
rect 8318 23326 8370 23378
rect 8766 23326 8818 23378
rect 9998 23326 10050 23378
rect 12910 23326 12962 23378
rect 13694 23326 13746 23378
rect 14142 23326 14194 23378
rect 14814 23326 14866 23378
rect 15822 23326 15874 23378
rect 15934 23326 15986 23378
rect 16046 23326 16098 23378
rect 18846 23326 18898 23378
rect 22990 23326 23042 23378
rect 23886 23326 23938 23378
rect 24670 23326 24722 23378
rect 25790 23326 25842 23378
rect 9886 23214 9938 23266
rect 10222 23214 10274 23266
rect 10894 23214 10946 23266
rect 11790 23214 11842 23266
rect 12686 23214 12738 23266
rect 13806 23214 13858 23266
rect 18286 23214 18338 23266
rect 19070 23214 19122 23266
rect 20302 23214 20354 23266
rect 23550 23214 23602 23266
rect 29150 23214 29202 23266
rect 1822 23102 1874 23154
rect 5182 23102 5234 23154
rect 5854 23102 5906 23154
rect 6078 23102 6130 23154
rect 10334 23102 10386 23154
rect 10670 23102 10722 23154
rect 11454 23102 11506 23154
rect 12126 23102 12178 23154
rect 12462 23102 12514 23154
rect 13470 23102 13522 23154
rect 14478 23102 14530 23154
rect 15038 23102 15090 23154
rect 15374 23102 15426 23154
rect 18622 23102 18674 23154
rect 19182 23102 19234 23154
rect 19518 23102 19570 23154
rect 24446 23102 24498 23154
rect 25230 23102 25282 23154
rect 25454 23102 25506 23154
rect 30046 23102 30098 23154
rect 2494 22990 2546 23042
rect 4622 22990 4674 23042
rect 4958 22990 5010 23042
rect 8430 22990 8482 23042
rect 8878 22990 8930 23042
rect 10782 22990 10834 23042
rect 11678 22990 11730 23042
rect 12574 22990 12626 23042
rect 17950 22990 18002 23042
rect 26798 22990 26850 23042
rect 6302 22878 6354 22930
rect 6414 22878 6466 22930
rect 11342 22878 11394 22930
rect 17390 22878 17442 22930
rect 17726 22878 17778 22930
rect 5372 22710 5424 22762
rect 5476 22710 5528 22762
rect 5580 22710 5632 22762
rect 13688 22710 13740 22762
rect 13792 22710 13844 22762
rect 13896 22710 13948 22762
rect 22004 22710 22056 22762
rect 22108 22710 22160 22762
rect 22212 22710 22264 22762
rect 30320 22710 30372 22762
rect 30424 22710 30476 22762
rect 30528 22710 30580 22762
rect 5630 22542 5682 22594
rect 5742 22542 5794 22594
rect 20302 22542 20354 22594
rect 26126 22542 26178 22594
rect 26462 22542 26514 22594
rect 2718 22430 2770 22482
rect 4846 22430 4898 22482
rect 7870 22430 7922 22482
rect 24446 22430 24498 22482
rect 26686 22430 26738 22482
rect 27134 22430 27186 22482
rect 1934 22318 1986 22370
rect 5966 22318 6018 22370
rect 6078 22318 6130 22370
rect 12910 22318 12962 22370
rect 17502 22318 17554 22370
rect 19294 22318 19346 22370
rect 20078 22318 20130 22370
rect 20414 22318 20466 22370
rect 21534 22318 21586 22370
rect 25566 22318 25618 22370
rect 26910 22318 26962 22370
rect 27918 22318 27970 22370
rect 15598 22206 15650 22258
rect 19630 22206 19682 22258
rect 20638 22206 20690 22258
rect 20750 22206 20802 22258
rect 22206 22206 22258 22258
rect 25678 22094 25730 22146
rect 25902 22094 25954 22146
rect 27246 22094 27298 22146
rect 27470 22094 27522 22146
rect 27806 22094 27858 22146
rect 9530 21926 9582 21978
rect 9634 21926 9686 21978
rect 9738 21926 9790 21978
rect 17846 21926 17898 21978
rect 17950 21926 18002 21978
rect 18054 21926 18106 21978
rect 26162 21926 26214 21978
rect 26266 21926 26318 21978
rect 26370 21926 26422 21978
rect 34478 21926 34530 21978
rect 34582 21926 34634 21978
rect 34686 21926 34738 21978
rect 3614 21758 3666 21810
rect 5070 21758 5122 21810
rect 5518 21758 5570 21810
rect 11230 21758 11282 21810
rect 11342 21758 11394 21810
rect 12686 21758 12738 21810
rect 13582 21758 13634 21810
rect 13694 21758 13746 21810
rect 13806 21758 13858 21810
rect 14702 21758 14754 21810
rect 14926 21758 14978 21810
rect 15710 21758 15762 21810
rect 16382 21758 16434 21810
rect 17950 21758 18002 21810
rect 19406 21758 19458 21810
rect 19966 21758 20018 21810
rect 20862 21758 20914 21810
rect 20974 21758 21026 21810
rect 24446 21758 24498 21810
rect 25454 21758 25506 21810
rect 3950 21646 4002 21698
rect 4622 21646 4674 21698
rect 5406 21646 5458 21698
rect 10782 21646 10834 21698
rect 12350 21646 12402 21698
rect 13470 21646 13522 21698
rect 14814 21646 14866 21698
rect 16718 21646 16770 21698
rect 19294 21646 19346 21698
rect 20526 21646 20578 21698
rect 20750 21646 20802 21698
rect 21646 21646 21698 21698
rect 25566 21646 25618 21698
rect 3390 21534 3442 21586
rect 3614 21534 3666 21586
rect 4398 21534 4450 21586
rect 4510 21534 4562 21586
rect 5742 21534 5794 21586
rect 10558 21534 10610 21586
rect 10894 21534 10946 21586
rect 11566 21534 11618 21586
rect 11902 21534 11954 21586
rect 13134 21534 13186 21586
rect 14142 21534 14194 21586
rect 14478 21534 14530 21586
rect 15150 21534 15202 21586
rect 15486 21534 15538 21586
rect 17614 21534 17666 21586
rect 18174 21534 18226 21586
rect 19630 21534 19682 21586
rect 20190 21534 20242 21586
rect 21198 21534 21250 21586
rect 21758 21534 21810 21586
rect 21982 21534 22034 21586
rect 23886 21534 23938 21586
rect 24446 21534 24498 21586
rect 29710 21534 29762 21586
rect 15374 21422 15426 21474
rect 22766 21422 22818 21474
rect 24670 21422 24722 21474
rect 26126 21422 26178 21474
rect 28814 21422 28866 21474
rect 17278 21310 17330 21362
rect 17726 21310 17778 21362
rect 25454 21310 25506 21362
rect 5372 21142 5424 21194
rect 5476 21142 5528 21194
rect 5580 21142 5632 21194
rect 13688 21142 13740 21194
rect 13792 21142 13844 21194
rect 13896 21142 13948 21194
rect 22004 21142 22056 21194
rect 22108 21142 22160 21194
rect 22212 21142 22264 21194
rect 30320 21142 30372 21194
rect 30424 21142 30476 21194
rect 30528 21142 30580 21194
rect 2606 20974 2658 21026
rect 11454 20974 11506 21026
rect 12798 20974 12850 21026
rect 22542 20974 22594 21026
rect 11006 20862 11058 20914
rect 12350 20862 12402 20914
rect 15822 20862 15874 20914
rect 22654 20862 22706 20914
rect 26014 20862 26066 20914
rect 27470 20862 27522 20914
rect 3278 20750 3330 20802
rect 4958 20750 5010 20802
rect 5630 20750 5682 20802
rect 7646 20750 7698 20802
rect 13806 20750 13858 20802
rect 14142 20750 14194 20802
rect 16046 20750 16098 20802
rect 17614 20750 17666 20802
rect 18174 20750 18226 20802
rect 22878 20750 22930 20802
rect 27022 20750 27074 20802
rect 27358 20750 27410 20802
rect 27582 20750 27634 20802
rect 3950 20638 4002 20690
rect 5742 20638 5794 20690
rect 8206 20638 8258 20690
rect 10558 20638 10610 20690
rect 10670 20638 10722 20690
rect 11342 20638 11394 20690
rect 12686 20638 12738 20690
rect 13470 20638 13522 20690
rect 13582 20638 13634 20690
rect 14366 20638 14418 20690
rect 17390 20638 17442 20690
rect 23774 20638 23826 20690
rect 2382 20526 2434 20578
rect 2494 20526 2546 20578
rect 2942 20526 2994 20578
rect 3614 20526 3666 20578
rect 4286 20526 4338 20578
rect 4398 20526 4450 20578
rect 4510 20526 4562 20578
rect 8094 20526 8146 20578
rect 10222 20526 10274 20578
rect 10446 20526 10498 20578
rect 11454 20526 11506 20578
rect 12798 20526 12850 20578
rect 16382 20526 16434 20578
rect 18398 20526 18450 20578
rect 21422 20526 21474 20578
rect 9530 20358 9582 20410
rect 9634 20358 9686 20410
rect 9738 20358 9790 20410
rect 17846 20358 17898 20410
rect 17950 20358 18002 20410
rect 18054 20358 18106 20410
rect 26162 20358 26214 20410
rect 26266 20358 26318 20410
rect 26370 20358 26422 20410
rect 34478 20358 34530 20410
rect 34582 20358 34634 20410
rect 34686 20358 34738 20410
rect 12798 20190 12850 20242
rect 26686 20190 26738 20242
rect 2494 20078 2546 20130
rect 8206 20078 8258 20130
rect 8878 20078 8930 20130
rect 10334 20078 10386 20130
rect 12014 20078 12066 20130
rect 12462 20078 12514 20130
rect 12574 20078 12626 20130
rect 14030 20078 14082 20130
rect 15038 20078 15090 20130
rect 15374 20078 15426 20130
rect 16830 20078 16882 20130
rect 23998 20078 24050 20130
rect 24446 20078 24498 20130
rect 1822 19966 1874 20018
rect 4846 19966 4898 20018
rect 5182 19966 5234 20018
rect 5406 19966 5458 20018
rect 7758 19966 7810 20018
rect 9774 19966 9826 20018
rect 10558 19966 10610 20018
rect 10782 19966 10834 20018
rect 11454 19966 11506 20018
rect 11902 19966 11954 20018
rect 12126 19966 12178 20018
rect 14254 19966 14306 20018
rect 14814 19966 14866 20018
rect 15710 19966 15762 20018
rect 16606 19966 16658 20018
rect 17726 19966 17778 20018
rect 18062 19966 18114 20018
rect 18174 19966 18226 20018
rect 18286 19966 18338 20018
rect 18622 19966 18674 20018
rect 18958 19966 19010 20018
rect 19182 19966 19234 20018
rect 20638 19966 20690 20018
rect 21086 19966 21138 20018
rect 22206 19966 22258 20018
rect 22990 19966 23042 20018
rect 24670 19966 24722 20018
rect 25230 19966 25282 20018
rect 25902 19966 25954 20018
rect 27134 19966 27186 20018
rect 30606 19966 30658 20018
rect 4622 19854 4674 19906
rect 5070 19854 5122 19906
rect 7310 19854 7362 19906
rect 9662 19854 9714 19906
rect 16158 19854 16210 19906
rect 19070 19854 19122 19906
rect 21534 19854 21586 19906
rect 21870 19854 21922 19906
rect 24334 19854 24386 19906
rect 25678 19854 25730 19906
rect 27806 19854 27858 19906
rect 29934 19854 29986 19906
rect 8654 19742 8706 19794
rect 8990 19742 9042 19794
rect 22206 19742 22258 19794
rect 27134 19742 27186 19794
rect 27470 19742 27522 19794
rect 5372 19574 5424 19626
rect 5476 19574 5528 19626
rect 5580 19574 5632 19626
rect 13688 19574 13740 19626
rect 13792 19574 13844 19626
rect 13896 19574 13948 19626
rect 22004 19574 22056 19626
rect 22108 19574 22160 19626
rect 22212 19574 22264 19626
rect 30320 19574 30372 19626
rect 30424 19574 30476 19626
rect 30528 19574 30580 19626
rect 12686 19406 12738 19458
rect 17614 19406 17666 19458
rect 2494 19294 2546 19346
rect 4622 19294 4674 19346
rect 7982 19294 8034 19346
rect 8990 19294 9042 19346
rect 9438 19294 9490 19346
rect 9774 19294 9826 19346
rect 11342 19294 11394 19346
rect 17390 19294 17442 19346
rect 18398 19294 18450 19346
rect 22318 19294 22370 19346
rect 24558 19294 24610 19346
rect 26462 19294 26514 19346
rect 28590 19294 28642 19346
rect 1822 19182 1874 19234
rect 7086 19182 7138 19234
rect 7534 19182 7586 19234
rect 8654 19182 8706 19234
rect 8878 19182 8930 19234
rect 9214 19182 9266 19234
rect 10782 19182 10834 19234
rect 12238 19182 12290 19234
rect 21646 19182 21698 19234
rect 25678 19182 25730 19234
rect 29150 19182 29202 19234
rect 29822 19182 29874 19234
rect 9998 19070 10050 19122
rect 10558 19070 10610 19122
rect 11230 19070 11282 19122
rect 12798 19070 12850 19122
rect 15038 19070 15090 19122
rect 11006 18958 11058 19010
rect 11902 18958 11954 19010
rect 12126 18958 12178 19010
rect 12350 18958 12402 19010
rect 17950 18958 18002 19010
rect 29262 18958 29314 19010
rect 29374 18958 29426 19010
rect 9530 18790 9582 18842
rect 9634 18790 9686 18842
rect 9738 18790 9790 18842
rect 17846 18790 17898 18842
rect 17950 18790 18002 18842
rect 18054 18790 18106 18842
rect 26162 18790 26214 18842
rect 26266 18790 26318 18842
rect 26370 18790 26422 18842
rect 34478 18790 34530 18842
rect 34582 18790 34634 18842
rect 34686 18790 34738 18842
rect 7422 18622 7474 18674
rect 8206 18622 8258 18674
rect 10782 18622 10834 18674
rect 11454 18622 11506 18674
rect 12686 18622 12738 18674
rect 6526 18510 6578 18562
rect 7982 18510 8034 18562
rect 8766 18510 8818 18562
rect 8878 18510 8930 18562
rect 9550 18510 9602 18562
rect 9662 18510 9714 18562
rect 19518 18510 19570 18562
rect 23214 18510 23266 18562
rect 30718 18510 30770 18562
rect 6302 18398 6354 18450
rect 7870 18398 7922 18450
rect 8318 18398 8370 18450
rect 9886 18398 9938 18450
rect 10558 18398 10610 18450
rect 10670 18398 10722 18450
rect 11230 18398 11282 18450
rect 11454 18398 11506 18450
rect 11790 18398 11842 18450
rect 14030 18398 14082 18450
rect 17390 18398 17442 18450
rect 17614 18398 17666 18450
rect 17950 18398 18002 18450
rect 18734 18398 18786 18450
rect 22878 18398 22930 18450
rect 23550 18398 23602 18450
rect 26126 18398 26178 18450
rect 26798 18398 26850 18450
rect 27134 18398 27186 18450
rect 6862 18286 6914 18338
rect 8206 18286 8258 18338
rect 10334 18286 10386 18338
rect 12126 18286 12178 18338
rect 12350 18286 12402 18338
rect 14702 18286 14754 18338
rect 16830 18286 16882 18338
rect 17502 18286 17554 18338
rect 21646 18286 21698 18338
rect 25454 18286 25506 18338
rect 25902 18286 25954 18338
rect 7086 18174 7138 18226
rect 8878 18174 8930 18226
rect 10110 18174 10162 18226
rect 5372 18006 5424 18058
rect 5476 18006 5528 18058
rect 5580 18006 5632 18058
rect 13688 18006 13740 18058
rect 13792 18006 13844 18058
rect 13896 18006 13948 18058
rect 22004 18006 22056 18058
rect 22108 18006 22160 18058
rect 22212 18006 22264 18058
rect 30320 18006 30372 18058
rect 30424 18006 30476 18058
rect 30528 18006 30580 18058
rect 6862 17838 6914 17890
rect 9550 17838 9602 17890
rect 9886 17838 9938 17890
rect 10782 17838 10834 17890
rect 29710 17838 29762 17890
rect 4622 17726 4674 17778
rect 8430 17726 8482 17778
rect 16046 17726 16098 17778
rect 17054 17726 17106 17778
rect 23550 17726 23602 17778
rect 33294 17726 33346 17778
rect 1822 17614 1874 17666
rect 5742 17614 5794 17666
rect 6302 17614 6354 17666
rect 6526 17614 6578 17666
rect 7646 17614 7698 17666
rect 7870 17614 7922 17666
rect 9102 17614 9154 17666
rect 10222 17614 10274 17666
rect 10894 17614 10946 17666
rect 15822 17614 15874 17666
rect 16158 17614 16210 17666
rect 16494 17614 16546 17666
rect 26686 17614 26738 17666
rect 29374 17614 29426 17666
rect 30494 17614 30546 17666
rect 2494 17502 2546 17554
rect 5966 17502 6018 17554
rect 7198 17502 7250 17554
rect 9774 17502 9826 17554
rect 10670 17502 10722 17554
rect 11230 17502 11282 17554
rect 17502 17502 17554 17554
rect 18174 17502 18226 17554
rect 18958 17502 19010 17554
rect 29150 17502 29202 17554
rect 31166 17502 31218 17554
rect 5070 17390 5122 17442
rect 7310 17390 7362 17442
rect 8878 17390 8930 17442
rect 10446 17390 10498 17442
rect 11118 17390 11170 17442
rect 17838 17390 17890 17442
rect 18510 17390 18562 17442
rect 19070 17390 19122 17442
rect 22542 17390 22594 17442
rect 9530 17222 9582 17274
rect 9634 17222 9686 17274
rect 9738 17222 9790 17274
rect 17846 17222 17898 17274
rect 17950 17222 18002 17274
rect 18054 17222 18106 17274
rect 26162 17222 26214 17274
rect 26266 17222 26318 17274
rect 26370 17222 26422 17274
rect 34478 17222 34530 17274
rect 34582 17222 34634 17274
rect 34686 17222 34738 17274
rect 7086 17054 7138 17106
rect 7646 17054 7698 17106
rect 8206 17054 8258 17106
rect 8430 17054 8482 17106
rect 8654 17054 8706 17106
rect 9886 17054 9938 17106
rect 14366 17054 14418 17106
rect 15262 17054 15314 17106
rect 15822 17054 15874 17106
rect 17390 17054 17442 17106
rect 29598 17054 29650 17106
rect 30046 17054 30098 17106
rect 31950 17054 32002 17106
rect 6750 16942 6802 16994
rect 8094 16942 8146 16994
rect 14142 16942 14194 16994
rect 15934 16942 15986 16994
rect 16718 16942 16770 16994
rect 17614 16942 17666 16994
rect 17726 16942 17778 16994
rect 17950 16942 18002 16994
rect 20638 16942 20690 16994
rect 29374 16942 29426 16994
rect 30382 16942 30434 16994
rect 3278 16830 3330 16882
rect 3950 16830 4002 16882
rect 7534 16830 7586 16882
rect 8878 16830 8930 16882
rect 9550 16830 9602 16882
rect 12238 16830 12290 16882
rect 12350 16830 12402 16882
rect 13582 16830 13634 16882
rect 13918 16830 13970 16882
rect 15374 16830 15426 16882
rect 15710 16830 15762 16882
rect 16382 16830 16434 16882
rect 16830 16830 16882 16882
rect 21310 16830 21362 16882
rect 24558 16830 24610 16882
rect 25342 16830 25394 16882
rect 29262 16830 29314 16882
rect 29710 16830 29762 16882
rect 31502 16830 31554 16882
rect 32174 16830 32226 16882
rect 6078 16718 6130 16770
rect 12798 16718 12850 16770
rect 14030 16718 14082 16770
rect 18174 16718 18226 16770
rect 18510 16718 18562 16770
rect 21758 16718 21810 16770
rect 23886 16718 23938 16770
rect 26014 16718 26066 16770
rect 28142 16718 28194 16770
rect 32062 16718 32114 16770
rect 7646 16606 7698 16658
rect 12686 16606 12738 16658
rect 15262 16606 15314 16658
rect 16718 16606 16770 16658
rect 5372 16438 5424 16490
rect 5476 16438 5528 16490
rect 5580 16438 5632 16490
rect 13688 16438 13740 16490
rect 13792 16438 13844 16490
rect 13896 16438 13948 16490
rect 22004 16438 22056 16490
rect 22108 16438 22160 16490
rect 22212 16438 22264 16490
rect 30320 16438 30372 16490
rect 30424 16438 30476 16490
rect 30528 16438 30580 16490
rect 17950 16270 18002 16322
rect 27470 16270 27522 16322
rect 30158 16270 30210 16322
rect 5070 16158 5122 16210
rect 10782 16158 10834 16210
rect 12910 16158 12962 16210
rect 13694 16158 13746 16210
rect 17390 16158 17442 16210
rect 23438 16158 23490 16210
rect 24446 16158 24498 16210
rect 29262 16158 29314 16210
rect 34190 16158 34242 16210
rect 2270 16046 2322 16098
rect 9998 16046 10050 16098
rect 13806 16046 13858 16098
rect 15150 16046 15202 16098
rect 15486 16046 15538 16098
rect 15710 16046 15762 16098
rect 15934 16046 15986 16098
rect 16158 16046 16210 16098
rect 16606 16046 16658 16098
rect 17278 16046 17330 16098
rect 17726 16046 17778 16098
rect 19294 16046 19346 16098
rect 21870 16046 21922 16098
rect 22430 16046 22482 16098
rect 23662 16046 23714 16098
rect 26238 16046 26290 16098
rect 27582 16046 27634 16098
rect 29374 16046 29426 16098
rect 29822 16046 29874 16098
rect 31278 16046 31330 16098
rect 2942 15934 2994 15986
rect 14142 15934 14194 15986
rect 14814 15934 14866 15986
rect 15038 15934 15090 15986
rect 16046 15934 16098 15986
rect 16942 15934 16994 15986
rect 18734 15934 18786 15986
rect 21534 15934 21586 15986
rect 22206 15934 22258 15986
rect 22654 15934 22706 15986
rect 22766 15934 22818 15986
rect 24334 15934 24386 15986
rect 24558 15934 24610 15986
rect 26126 15934 26178 15986
rect 27918 15934 27970 15986
rect 28366 15934 28418 15986
rect 29150 15934 29202 15986
rect 30046 15934 30098 15986
rect 32062 15934 32114 15986
rect 5742 15822 5794 15874
rect 6302 15822 6354 15874
rect 9662 15822 9714 15874
rect 14254 15822 14306 15874
rect 14478 15822 14530 15874
rect 16830 15822 16882 15874
rect 18286 15822 18338 15874
rect 18846 15822 18898 15874
rect 19070 15822 19122 15874
rect 21646 15822 21698 15874
rect 23998 15822 24050 15874
rect 26014 15822 26066 15874
rect 27470 15822 27522 15874
rect 28142 15822 28194 15874
rect 28478 15822 28530 15874
rect 9530 15654 9582 15706
rect 9634 15654 9686 15706
rect 9738 15654 9790 15706
rect 17846 15654 17898 15706
rect 17950 15654 18002 15706
rect 18054 15654 18106 15706
rect 26162 15654 26214 15706
rect 26266 15654 26318 15706
rect 26370 15654 26422 15706
rect 34478 15654 34530 15706
rect 34582 15654 34634 15706
rect 34686 15654 34738 15706
rect 14926 15486 14978 15538
rect 15486 15486 15538 15538
rect 15710 15486 15762 15538
rect 30382 15486 30434 15538
rect 33070 15486 33122 15538
rect 11902 15374 11954 15426
rect 16270 15374 16322 15426
rect 16718 15374 16770 15426
rect 16830 15374 16882 15426
rect 20190 15374 20242 15426
rect 26126 15374 26178 15426
rect 26350 15374 26402 15426
rect 30942 15374 30994 15426
rect 32062 15374 32114 15426
rect 32286 15374 32338 15426
rect 5742 15262 5794 15314
rect 8990 15262 9042 15314
rect 11230 15262 11282 15314
rect 14814 15262 14866 15314
rect 15262 15262 15314 15314
rect 15934 15262 15986 15314
rect 17950 15262 18002 15314
rect 18174 15262 18226 15314
rect 28814 15262 28866 15314
rect 31054 15262 31106 15314
rect 31502 15262 31554 15314
rect 31726 15262 31778 15314
rect 33630 15262 33682 15314
rect 6414 15150 6466 15202
rect 8542 15150 8594 15202
rect 14030 15150 14082 15202
rect 15374 15150 15426 15202
rect 26014 15150 26066 15202
rect 30494 15150 30546 15202
rect 30606 15150 30658 15202
rect 32398 15150 32450 15202
rect 33406 15150 33458 15202
rect 16382 15038 16434 15090
rect 28478 15038 28530 15090
rect 28814 15038 28866 15090
rect 31278 15038 31330 15090
rect 5372 14870 5424 14922
rect 5476 14870 5528 14922
rect 5580 14870 5632 14922
rect 13688 14870 13740 14922
rect 13792 14870 13844 14922
rect 13896 14870 13948 14922
rect 22004 14870 22056 14922
rect 22108 14870 22160 14922
rect 22212 14870 22264 14922
rect 30320 14870 30372 14922
rect 30424 14870 30476 14922
rect 30528 14870 30580 14922
rect 18622 14702 18674 14754
rect 28254 14702 28306 14754
rect 30830 14702 30882 14754
rect 32174 14702 32226 14754
rect 32734 14702 32786 14754
rect 32846 14702 32898 14754
rect 4622 14590 4674 14642
rect 18734 14590 18786 14642
rect 20638 14590 20690 14642
rect 21310 14590 21362 14642
rect 23438 14590 23490 14642
rect 1822 14478 1874 14530
rect 12686 14478 12738 14530
rect 16158 14478 16210 14530
rect 16942 14478 16994 14530
rect 17278 14478 17330 14530
rect 20750 14478 20802 14530
rect 24222 14478 24274 14530
rect 27246 14478 27298 14530
rect 27582 14478 27634 14530
rect 27806 14478 27858 14530
rect 31166 14478 31218 14530
rect 31278 14478 31330 14530
rect 31614 14478 31666 14530
rect 31838 14478 31890 14530
rect 33070 14478 33122 14530
rect 2494 14366 2546 14418
rect 8430 14366 8482 14418
rect 13582 14366 13634 14418
rect 15822 14366 15874 14418
rect 16494 14366 16546 14418
rect 17726 14366 17778 14418
rect 19070 14366 19122 14418
rect 19518 14366 19570 14418
rect 19630 14366 19682 14418
rect 20078 14366 20130 14418
rect 27470 14366 27522 14418
rect 29150 14366 29202 14418
rect 30718 14366 30770 14418
rect 5070 14254 5122 14306
rect 5630 14254 5682 14306
rect 5966 14254 6018 14306
rect 15934 14254 15986 14306
rect 19854 14254 19906 14306
rect 20302 14254 20354 14306
rect 20526 14254 20578 14306
rect 29486 14254 29538 14306
rect 32734 14254 32786 14306
rect 9530 14086 9582 14138
rect 9634 14086 9686 14138
rect 9738 14086 9790 14138
rect 17846 14086 17898 14138
rect 17950 14086 18002 14138
rect 18054 14086 18106 14138
rect 26162 14086 26214 14138
rect 26266 14086 26318 14138
rect 26370 14086 26422 14138
rect 34478 14086 34530 14138
rect 34582 14086 34634 14138
rect 34686 14086 34738 14138
rect 6750 13918 6802 13970
rect 9774 13918 9826 13970
rect 14142 13918 14194 13970
rect 16830 13918 16882 13970
rect 18398 13918 18450 13970
rect 18846 13918 18898 13970
rect 19854 13918 19906 13970
rect 22878 13918 22930 13970
rect 23662 13918 23714 13970
rect 24222 13918 24274 13970
rect 31166 13918 31218 13970
rect 32286 13918 32338 13970
rect 5966 13806 6018 13858
rect 7310 13806 7362 13858
rect 7422 13806 7474 13858
rect 9998 13806 10050 13858
rect 10110 13806 10162 13858
rect 10894 13806 10946 13858
rect 11118 13806 11170 13858
rect 15934 13806 15986 13858
rect 17390 13806 17442 13858
rect 17726 13806 17778 13858
rect 20526 13806 20578 13858
rect 25678 13806 25730 13858
rect 5518 13694 5570 13746
rect 6302 13694 6354 13746
rect 6526 13694 6578 13746
rect 6862 13694 6914 13746
rect 9550 13694 9602 13746
rect 11342 13694 11394 13746
rect 15262 13694 15314 13746
rect 15822 13694 15874 13746
rect 18174 13694 18226 13746
rect 19630 13694 19682 13746
rect 20190 13694 20242 13746
rect 22206 13694 22258 13746
rect 22654 13694 22706 13746
rect 23550 13694 23602 13746
rect 23886 13694 23938 13746
rect 25454 13694 25506 13746
rect 26126 13694 26178 13746
rect 26350 13694 26402 13746
rect 26686 13694 26738 13746
rect 27022 13694 27074 13746
rect 27358 13694 27410 13746
rect 30718 13694 30770 13746
rect 31726 13694 31778 13746
rect 33182 13694 33234 13746
rect 33630 13694 33682 13746
rect 5630 13582 5682 13634
rect 7758 13582 7810 13634
rect 7982 13582 8034 13634
rect 10222 13582 10274 13634
rect 11902 13582 11954 13634
rect 26462 13582 26514 13634
rect 27246 13582 27298 13634
rect 27806 13582 27858 13634
rect 29934 13582 29986 13634
rect 31278 13582 31330 13634
rect 7310 13470 7362 13522
rect 11790 13470 11842 13522
rect 21310 13470 21362 13522
rect 21758 13470 21810 13522
rect 21982 13470 22034 13522
rect 26910 13470 26962 13522
rect 31390 13470 31442 13522
rect 31950 13470 32002 13522
rect 33294 13470 33346 13522
rect 33518 13470 33570 13522
rect 5372 13302 5424 13354
rect 5476 13302 5528 13354
rect 5580 13302 5632 13354
rect 13688 13302 13740 13354
rect 13792 13302 13844 13354
rect 13896 13302 13948 13354
rect 22004 13302 22056 13354
rect 22108 13302 22160 13354
rect 22212 13302 22264 13354
rect 30320 13302 30372 13354
rect 30424 13302 30476 13354
rect 30528 13302 30580 13354
rect 6526 13134 6578 13186
rect 20302 13134 20354 13186
rect 22094 13134 22146 13186
rect 29598 13134 29650 13186
rect 29710 13134 29762 13186
rect 3726 13022 3778 13074
rect 4622 13022 4674 13074
rect 5630 13022 5682 13074
rect 10782 13022 10834 13074
rect 11230 13022 11282 13074
rect 12126 13022 12178 13074
rect 12574 13022 12626 13074
rect 20078 13022 20130 13074
rect 22990 13022 23042 13074
rect 24782 13022 24834 13074
rect 26910 13022 26962 13074
rect 28590 13022 28642 13074
rect 31278 13022 31330 13074
rect 33406 13022 33458 13074
rect 4286 12910 4338 12962
rect 5854 12910 5906 12962
rect 6078 12910 6130 12962
rect 7870 12910 7922 12962
rect 11678 12910 11730 12962
rect 16046 12910 16098 12962
rect 16606 12910 16658 12962
rect 16942 12910 16994 12962
rect 17614 12910 17666 12962
rect 18286 12910 18338 12962
rect 18958 12910 19010 12962
rect 19518 12910 19570 12962
rect 20526 12910 20578 12962
rect 20862 12910 20914 12962
rect 21870 12910 21922 12962
rect 22318 12910 22370 12962
rect 24110 12910 24162 12962
rect 27470 12910 27522 12962
rect 28030 12910 28082 12962
rect 28366 12910 28418 12962
rect 29150 12910 29202 12962
rect 29374 12910 29426 12962
rect 34078 12910 34130 12962
rect 7198 12798 7250 12850
rect 7534 12798 7586 12850
rect 8654 12798 8706 12850
rect 14142 12798 14194 12850
rect 17390 12798 17442 12850
rect 18622 12798 18674 12850
rect 19854 12798 19906 12850
rect 21646 12798 21698 12850
rect 22542 12798 22594 12850
rect 22878 12798 22930 12850
rect 27358 12798 27410 12850
rect 3390 12686 3442 12738
rect 3614 12686 3666 12738
rect 3838 12686 3890 12738
rect 5070 12686 5122 12738
rect 11118 12686 11170 12738
rect 11342 12686 11394 12738
rect 12014 12686 12066 12738
rect 13806 12686 13858 12738
rect 14590 12686 14642 12738
rect 16270 12686 16322 12738
rect 18510 12686 18562 12738
rect 19294 12686 19346 12738
rect 19406 12686 19458 12738
rect 19742 12686 19794 12738
rect 22094 12686 22146 12738
rect 27134 12686 27186 12738
rect 9530 12518 9582 12570
rect 9634 12518 9686 12570
rect 9738 12518 9790 12570
rect 17846 12518 17898 12570
rect 17950 12518 18002 12570
rect 18054 12518 18106 12570
rect 26162 12518 26214 12570
rect 26266 12518 26318 12570
rect 26370 12518 26422 12570
rect 34478 12518 34530 12570
rect 34582 12518 34634 12570
rect 34686 12518 34738 12570
rect 4174 12350 4226 12402
rect 5406 12350 5458 12402
rect 5518 12350 5570 12402
rect 20638 12350 20690 12402
rect 20974 12350 21026 12402
rect 3166 12238 3218 12290
rect 3726 12238 3778 12290
rect 4958 12238 5010 12290
rect 8654 12238 8706 12290
rect 8990 12238 9042 12290
rect 10670 12238 10722 12290
rect 18174 12238 18226 12290
rect 22094 12238 22146 12290
rect 2830 12126 2882 12178
rect 4174 12126 4226 12178
rect 4510 12126 4562 12178
rect 4622 12126 4674 12178
rect 5294 12126 5346 12178
rect 5854 12126 5906 12178
rect 6526 12126 6578 12178
rect 6974 12126 7026 12178
rect 7870 12126 7922 12178
rect 10222 12126 10274 12178
rect 10782 12126 10834 12178
rect 12686 12126 12738 12178
rect 17502 12126 17554 12178
rect 21422 12126 21474 12178
rect 26014 12126 26066 12178
rect 26574 12126 26626 12178
rect 31390 12126 31442 12178
rect 31838 12126 31890 12178
rect 3838 12014 3890 12066
rect 8206 12014 8258 12066
rect 10446 12014 10498 12066
rect 13582 12014 13634 12066
rect 20302 12014 20354 12066
rect 24222 12014 24274 12066
rect 26686 12014 26738 12066
rect 3502 11902 3554 11954
rect 31614 11902 31666 11954
rect 31950 11902 32002 11954
rect 5372 11734 5424 11786
rect 5476 11734 5528 11786
rect 5580 11734 5632 11786
rect 13688 11734 13740 11786
rect 13792 11734 13844 11786
rect 13896 11734 13948 11786
rect 22004 11734 22056 11786
rect 22108 11734 22160 11786
rect 22212 11734 22264 11786
rect 30320 11734 30372 11786
rect 30424 11734 30476 11786
rect 30528 11734 30580 11786
rect 6862 11566 6914 11618
rect 8542 11566 8594 11618
rect 17278 11566 17330 11618
rect 17614 11566 17666 11618
rect 18734 11566 18786 11618
rect 18958 11566 19010 11618
rect 20414 11566 20466 11618
rect 22878 11566 22930 11618
rect 2382 11454 2434 11506
rect 3054 11454 3106 11506
rect 4286 11454 4338 11506
rect 6414 11454 6466 11506
rect 10670 11454 10722 11506
rect 11342 11454 11394 11506
rect 14254 11454 14306 11506
rect 16382 11454 16434 11506
rect 18734 11454 18786 11506
rect 19070 11454 19122 11506
rect 20526 11454 20578 11506
rect 21534 11454 21586 11506
rect 22430 11454 22482 11506
rect 27358 11454 27410 11506
rect 31278 11454 31330 11506
rect 33406 11454 33458 11506
rect 2158 11342 2210 11394
rect 3278 11342 3330 11394
rect 3502 11342 3554 11394
rect 3614 11342 3666 11394
rect 4174 11342 4226 11394
rect 4622 11342 4674 11394
rect 4846 11342 4898 11394
rect 5518 11342 5570 11394
rect 5966 11342 6018 11394
rect 6078 11342 6130 11394
rect 6302 11342 6354 11394
rect 6526 11342 6578 11394
rect 7086 11342 7138 11394
rect 7534 11342 7586 11394
rect 8766 11342 8818 11394
rect 8878 11342 8930 11394
rect 9886 11342 9938 11394
rect 10446 11342 10498 11394
rect 10894 11342 10946 11394
rect 13470 11342 13522 11394
rect 17838 11342 17890 11394
rect 19406 11342 19458 11394
rect 19630 11342 19682 11394
rect 19854 11342 19906 11394
rect 20078 11342 20130 11394
rect 21982 11342 22034 11394
rect 22990 11342 23042 11394
rect 24446 11342 24498 11394
rect 29822 11342 29874 11394
rect 30270 11342 30322 11394
rect 34078 11342 34130 11394
rect 7422 11230 7474 11282
rect 8430 11230 8482 11282
rect 9326 11230 9378 11282
rect 10222 11230 10274 11282
rect 11118 11230 11170 11282
rect 16718 11230 16770 11282
rect 25230 11230 25282 11282
rect 2270 11118 2322 11170
rect 2494 11118 2546 11170
rect 2606 11118 2658 11170
rect 3726 11118 3778 11170
rect 4398 11118 4450 11170
rect 7310 11118 7362 11170
rect 11342 11118 11394 11170
rect 12910 11118 12962 11170
rect 16830 11118 16882 11170
rect 19742 11118 19794 11170
rect 29150 11118 29202 11170
rect 29262 11118 29314 11170
rect 29374 11118 29426 11170
rect 30046 11118 30098 11170
rect 9530 10950 9582 11002
rect 9634 10950 9686 11002
rect 9738 10950 9790 11002
rect 17846 10950 17898 11002
rect 17950 10950 18002 11002
rect 18054 10950 18106 11002
rect 26162 10950 26214 11002
rect 26266 10950 26318 11002
rect 26370 10950 26422 11002
rect 34478 10950 34530 11002
rect 34582 10950 34634 11002
rect 34686 10950 34738 11002
rect 3726 10782 3778 10834
rect 4734 10782 4786 10834
rect 4958 10782 5010 10834
rect 7310 10782 7362 10834
rect 7646 10782 7698 10834
rect 10334 10782 10386 10834
rect 10894 10782 10946 10834
rect 16942 10782 16994 10834
rect 17390 10782 17442 10834
rect 22542 10782 22594 10834
rect 25790 10782 25842 10834
rect 31390 10782 31442 10834
rect 3278 10670 3330 10722
rect 3838 10670 3890 10722
rect 6862 10670 6914 10722
rect 8990 10670 9042 10722
rect 10446 10670 10498 10722
rect 13022 10670 13074 10722
rect 22094 10670 22146 10722
rect 26014 10670 26066 10722
rect 31838 10670 31890 10722
rect 2718 10558 2770 10610
rect 3054 10558 3106 10610
rect 5070 10558 5122 10610
rect 6750 10558 6802 10610
rect 7086 10558 7138 10610
rect 8430 10558 8482 10610
rect 8878 10558 8930 10610
rect 9438 10558 9490 10610
rect 9886 10558 9938 10610
rect 9998 10558 10050 10610
rect 10782 10558 10834 10610
rect 11006 10558 11058 10610
rect 11230 10558 11282 10610
rect 12350 10558 12402 10610
rect 18510 10558 18562 10610
rect 21758 10558 21810 10610
rect 27134 10558 27186 10610
rect 30382 10558 30434 10610
rect 30494 10558 30546 10610
rect 30830 10558 30882 10610
rect 30942 10558 30994 10610
rect 32174 10558 32226 10610
rect 2942 10446 2994 10498
rect 10222 10446 10274 10498
rect 15150 10446 15202 10498
rect 17838 10446 17890 10498
rect 19182 10446 19234 10498
rect 21310 10446 21362 10498
rect 25678 10446 25730 10498
rect 27806 10446 27858 10498
rect 29934 10446 29986 10498
rect 3614 10334 3666 10386
rect 8654 10334 8706 10386
rect 21758 10334 21810 10386
rect 32174 10334 32226 10386
rect 5372 10166 5424 10218
rect 5476 10166 5528 10218
rect 5580 10166 5632 10218
rect 13688 10166 13740 10218
rect 13792 10166 13844 10218
rect 13896 10166 13948 10218
rect 22004 10166 22056 10218
rect 22108 10166 22160 10218
rect 22212 10166 22264 10218
rect 30320 10166 30372 10218
rect 30424 10166 30476 10218
rect 30528 10166 30580 10218
rect 2270 9998 2322 10050
rect 7982 9998 8034 10050
rect 9214 9998 9266 10050
rect 21310 9998 21362 10050
rect 3166 9886 3218 9938
rect 3614 9886 3666 9938
rect 6078 9886 6130 9938
rect 8878 9886 8930 9938
rect 10558 9886 10610 9938
rect 12014 9886 12066 9938
rect 12462 9886 12514 9938
rect 15822 9886 15874 9938
rect 21422 9886 21474 9938
rect 30830 9886 30882 9938
rect 31278 9886 31330 9938
rect 2718 9774 2770 9826
rect 2942 9774 2994 9826
rect 4062 9774 4114 9826
rect 5630 9774 5682 9826
rect 5966 9774 6018 9826
rect 9550 9774 9602 9826
rect 11454 9774 11506 9826
rect 11566 9774 11618 9826
rect 12910 9774 12962 9826
rect 13694 9774 13746 9826
rect 15710 9774 15762 9826
rect 17838 9774 17890 9826
rect 18174 9774 18226 9826
rect 20078 9774 20130 9826
rect 20638 9774 20690 9826
rect 22094 9774 22146 9826
rect 27246 9774 27298 9826
rect 29262 9774 29314 9826
rect 29710 9774 29762 9826
rect 30382 9774 30434 9826
rect 30942 9774 30994 9826
rect 34078 9774 34130 9826
rect 6190 9662 6242 9714
rect 7982 9662 8034 9714
rect 3502 9550 3554 9602
rect 3726 9550 3778 9602
rect 8094 9606 8146 9658
rect 8766 9662 8818 9714
rect 8990 9662 9042 9714
rect 9998 9662 10050 9714
rect 10334 9662 10386 9714
rect 10670 9662 10722 9714
rect 10894 9662 10946 9714
rect 11230 9662 11282 9714
rect 14142 9662 14194 9714
rect 17726 9662 17778 9714
rect 18622 9662 18674 9714
rect 18958 9662 19010 9714
rect 19630 9662 19682 9714
rect 21534 9662 21586 9714
rect 24446 9662 24498 9714
rect 29374 9662 29426 9714
rect 30606 9662 30658 9714
rect 33406 9662 33458 9714
rect 10110 9550 10162 9602
rect 13582 9550 13634 9602
rect 18286 9550 18338 9602
rect 28142 9550 28194 9602
rect 28478 9550 28530 9602
rect 29486 9550 29538 9602
rect 9530 9382 9582 9434
rect 9634 9382 9686 9434
rect 9738 9382 9790 9434
rect 17846 9382 17898 9434
rect 17950 9382 18002 9434
rect 18054 9382 18106 9434
rect 26162 9382 26214 9434
rect 26266 9382 26318 9434
rect 26370 9382 26422 9434
rect 34478 9382 34530 9434
rect 34582 9382 34634 9434
rect 34686 9382 34738 9434
rect 2830 9214 2882 9266
rect 3950 9214 4002 9266
rect 4622 9214 4674 9266
rect 5294 9214 5346 9266
rect 5406 9214 5458 9266
rect 7870 9214 7922 9266
rect 10670 9214 10722 9266
rect 23998 9214 24050 9266
rect 24670 9214 24722 9266
rect 26238 9214 26290 9266
rect 26574 9214 26626 9266
rect 33182 9214 33234 9266
rect 4398 9102 4450 9154
rect 5518 9102 5570 9154
rect 6526 9102 6578 9154
rect 9550 9102 9602 9154
rect 9774 9102 9826 9154
rect 12238 9102 12290 9154
rect 14814 9102 14866 9154
rect 18174 9102 18226 9154
rect 18958 9102 19010 9154
rect 21758 9102 21810 9154
rect 31838 9102 31890 9154
rect 3166 8990 3218 9042
rect 3502 8990 3554 9042
rect 3726 8990 3778 9042
rect 4286 8990 4338 9042
rect 5182 8990 5234 9042
rect 6414 8990 6466 9042
rect 6638 8990 6690 9042
rect 7086 8990 7138 9042
rect 7646 8990 7698 9042
rect 7758 8990 7810 9042
rect 8318 8990 8370 9042
rect 9998 8990 10050 9042
rect 10222 8990 10274 9042
rect 10894 8990 10946 9042
rect 11902 8990 11954 9042
rect 13246 8990 13298 9042
rect 13806 8990 13858 9042
rect 15710 8990 15762 9042
rect 17614 8990 17666 9042
rect 19070 8990 19122 9042
rect 20974 8990 21026 9042
rect 25566 8990 25618 9042
rect 27246 8990 27298 9042
rect 33070 8990 33122 9042
rect 33294 8990 33346 9042
rect 2382 8878 2434 8930
rect 10334 8878 10386 8930
rect 16046 8878 16098 8930
rect 16158 8878 16210 8930
rect 17726 8878 17778 8930
rect 25342 8878 25394 8930
rect 3726 8766 3778 8818
rect 4846 8766 4898 8818
rect 11342 8766 11394 8818
rect 11678 8766 11730 8818
rect 25230 8766 25282 8818
rect 33518 8766 33570 8818
rect 5372 8598 5424 8650
rect 5476 8598 5528 8650
rect 5580 8598 5632 8650
rect 13688 8598 13740 8650
rect 13792 8598 13844 8650
rect 13896 8598 13948 8650
rect 22004 8598 22056 8650
rect 22108 8598 22160 8650
rect 22212 8598 22264 8650
rect 30320 8598 30372 8650
rect 30424 8598 30476 8650
rect 30528 8598 30580 8650
rect 29934 8430 29986 8482
rect 2718 8318 2770 8370
rect 3838 8318 3890 8370
rect 5854 8318 5906 8370
rect 9214 8318 9266 8370
rect 13358 8318 13410 8370
rect 17950 8318 18002 8370
rect 19070 8318 19122 8370
rect 21422 8318 21474 8370
rect 22318 8318 22370 8370
rect 23774 8318 23826 8370
rect 25902 8318 25954 8370
rect 28142 8318 28194 8370
rect 30606 8318 30658 8370
rect 34190 8318 34242 8370
rect 3166 8206 3218 8258
rect 3390 8206 3442 8258
rect 3614 8206 3666 8258
rect 5630 8206 5682 8258
rect 6078 8206 6130 8258
rect 6526 8206 6578 8258
rect 6974 8206 7026 8258
rect 9886 8206 9938 8258
rect 12126 8206 12178 8258
rect 13470 8206 13522 8258
rect 15374 8206 15426 8258
rect 18286 8206 18338 8258
rect 18958 8206 19010 8258
rect 22094 8206 22146 8258
rect 23102 8206 23154 8258
rect 26910 8206 26962 8258
rect 27694 8206 27746 8258
rect 29486 8206 29538 8258
rect 29710 8206 29762 8258
rect 30158 8206 30210 8258
rect 30494 8206 30546 8258
rect 31390 8206 31442 8258
rect 2606 8094 2658 8146
rect 2830 8094 2882 8146
rect 3838 8094 3890 8146
rect 4846 8094 4898 8146
rect 6302 8094 6354 8146
rect 7198 8094 7250 8146
rect 7534 8094 7586 8146
rect 8654 8094 8706 8146
rect 8766 8094 8818 8146
rect 8878 8094 8930 8146
rect 9550 8094 9602 8146
rect 10110 8094 10162 8146
rect 10446 8094 10498 8146
rect 10782 8094 10834 8146
rect 11454 8094 11506 8146
rect 12462 8094 12514 8146
rect 12910 8094 12962 8146
rect 14926 8094 14978 8146
rect 16158 8094 16210 8146
rect 28030 8094 28082 8146
rect 29374 8094 29426 8146
rect 32062 8094 32114 8146
rect 4062 7982 4114 8034
rect 4510 7982 4562 8034
rect 5518 7982 5570 8034
rect 7086 7982 7138 8034
rect 7310 7982 7362 8034
rect 8430 7982 8482 8034
rect 9886 7982 9938 8034
rect 11118 7982 11170 8034
rect 11790 7982 11842 8034
rect 12350 7982 12402 8034
rect 12686 7982 12738 8034
rect 17166 7982 17218 8034
rect 21758 7982 21810 8034
rect 26238 7982 26290 8034
rect 26574 7982 26626 8034
rect 27246 7982 27298 8034
rect 28254 7982 28306 8034
rect 9530 7814 9582 7866
rect 9634 7814 9686 7866
rect 9738 7814 9790 7866
rect 17846 7814 17898 7866
rect 17950 7814 18002 7866
rect 18054 7814 18106 7866
rect 26162 7814 26214 7866
rect 26266 7814 26318 7866
rect 26370 7814 26422 7866
rect 34478 7814 34530 7866
rect 34582 7814 34634 7866
rect 34686 7814 34738 7866
rect 2494 7646 2546 7698
rect 2942 7646 2994 7698
rect 5182 7646 5234 7698
rect 6750 7646 6802 7698
rect 7646 7646 7698 7698
rect 4510 7534 4562 7586
rect 8878 7534 8930 7586
rect 9438 7534 9490 7586
rect 9662 7534 9714 7586
rect 9774 7590 9826 7642
rect 27582 7646 27634 7698
rect 28142 7646 28194 7698
rect 30718 7646 30770 7698
rect 32062 7646 32114 7698
rect 16270 7534 16322 7586
rect 22430 7534 22482 7586
rect 23326 7534 23378 7586
rect 23550 7534 23602 7586
rect 25902 7534 25954 7586
rect 28366 7534 28418 7586
rect 29486 7534 29538 7586
rect 29710 7534 29762 7586
rect 32174 7534 32226 7586
rect 32622 7534 32674 7586
rect 33182 7534 33234 7586
rect 2270 7422 2322 7474
rect 2830 7422 2882 7474
rect 3054 7422 3106 7474
rect 3502 7422 3554 7474
rect 3838 7422 3890 7474
rect 3950 7422 4002 7474
rect 4398 7422 4450 7474
rect 4734 7422 4786 7474
rect 5070 7422 5122 7474
rect 5294 7422 5346 7474
rect 5518 7422 5570 7474
rect 5742 7422 5794 7474
rect 6638 7422 6690 7474
rect 6862 7422 6914 7474
rect 7310 7422 7362 7474
rect 7870 7422 7922 7474
rect 8766 7422 8818 7474
rect 10670 7422 10722 7474
rect 11118 7422 11170 7474
rect 13022 7422 13074 7474
rect 13806 7422 13858 7474
rect 15038 7422 15090 7474
rect 16830 7422 16882 7474
rect 18062 7422 18114 7474
rect 18286 7422 18338 7474
rect 18846 7422 18898 7474
rect 21982 7422 22034 7474
rect 22206 7422 22258 7474
rect 22766 7422 22818 7474
rect 22990 7422 23042 7474
rect 25566 7422 25618 7474
rect 26014 7422 26066 7474
rect 26238 7422 26290 7474
rect 27470 7422 27522 7474
rect 27694 7422 27746 7474
rect 29150 7422 29202 7474
rect 29822 7422 29874 7474
rect 30270 7422 30322 7474
rect 31054 7422 31106 7474
rect 31278 7422 31330 7474
rect 31950 7422 32002 7474
rect 32174 7422 32226 7474
rect 33406 7422 33458 7474
rect 8318 7310 8370 7362
rect 12798 7310 12850 7362
rect 14478 7310 14530 7362
rect 17390 7310 17442 7362
rect 19518 7310 19570 7362
rect 21646 7310 21698 7362
rect 23438 7310 23490 7362
rect 4174 7198 4226 7250
rect 26686 7198 26738 7250
rect 27246 7198 27298 7250
rect 28030 7198 28082 7250
rect 31726 7198 31778 7250
rect 33070 7198 33122 7250
rect 5372 7030 5424 7082
rect 5476 7030 5528 7082
rect 5580 7030 5632 7082
rect 13688 7030 13740 7082
rect 13792 7030 13844 7082
rect 13896 7030 13948 7082
rect 22004 7030 22056 7082
rect 22108 7030 22160 7082
rect 22212 7030 22264 7082
rect 30320 7030 30372 7082
rect 30424 7030 30476 7082
rect 30528 7030 30580 7082
rect 3502 6750 3554 6802
rect 4958 6750 5010 6802
rect 5630 6750 5682 6802
rect 9662 6750 9714 6802
rect 10446 6750 10498 6802
rect 14030 6750 14082 6802
rect 18174 6750 18226 6802
rect 19182 6750 19234 6802
rect 22206 6750 22258 6802
rect 23774 6750 23826 6802
rect 29374 6750 29426 6802
rect 29710 6750 29762 6802
rect 30382 6750 30434 6802
rect 33966 6750 34018 6802
rect 5070 6638 5122 6690
rect 6190 6638 6242 6690
rect 8206 6638 8258 6690
rect 8542 6638 8594 6690
rect 9774 6638 9826 6690
rect 10222 6638 10274 6690
rect 11566 6638 11618 6690
rect 11902 6638 11954 6690
rect 12126 6638 12178 6690
rect 12238 6638 12290 6690
rect 14142 6638 14194 6690
rect 14702 6638 14754 6690
rect 15262 6638 15314 6690
rect 19742 6638 19794 6690
rect 22094 6638 22146 6690
rect 22318 6638 22370 6690
rect 23214 6638 23266 6690
rect 26462 6638 26514 6690
rect 27022 6638 27074 6690
rect 27246 6638 27298 6690
rect 27918 6638 27970 6690
rect 29150 6638 29202 6690
rect 30158 6638 30210 6690
rect 30718 6638 30770 6690
rect 31166 6638 31218 6690
rect 5742 6526 5794 6578
rect 6526 6526 6578 6578
rect 9102 6526 9154 6578
rect 11118 6526 11170 6578
rect 11454 6526 11506 6578
rect 12574 6526 12626 6578
rect 13806 6526 13858 6578
rect 16046 6526 16098 6578
rect 22990 6526 23042 6578
rect 24110 6526 24162 6578
rect 24782 6526 24834 6578
rect 26798 6526 26850 6578
rect 31838 6526 31890 6578
rect 3390 6414 3442 6466
rect 4622 6414 4674 6466
rect 4846 6414 4898 6466
rect 6190 6414 6242 6466
rect 7870 6414 7922 6466
rect 7982 6414 8034 6466
rect 9550 6414 9602 6466
rect 18734 6414 18786 6466
rect 27022 6414 27074 6466
rect 27694 6414 27746 6466
rect 9530 6246 9582 6298
rect 9634 6246 9686 6298
rect 9738 6246 9790 6298
rect 17846 6246 17898 6298
rect 17950 6246 18002 6298
rect 18054 6246 18106 6298
rect 26162 6246 26214 6298
rect 26266 6246 26318 6298
rect 26370 6246 26422 6298
rect 34478 6246 34530 6298
rect 34582 6246 34634 6298
rect 34686 6246 34738 6298
rect 3278 6078 3330 6130
rect 7870 6078 7922 6130
rect 7982 6078 8034 6130
rect 9662 6078 9714 6130
rect 11566 6078 11618 6130
rect 13582 6078 13634 6130
rect 17950 6078 18002 6130
rect 27694 6078 27746 6130
rect 4062 5966 4114 6018
rect 5854 5966 5906 6018
rect 6526 5966 6578 6018
rect 8430 5966 8482 6018
rect 8766 5966 8818 6018
rect 11118 5966 11170 6018
rect 12462 5966 12514 6018
rect 12798 5966 12850 6018
rect 13694 5966 13746 6018
rect 14254 5966 14306 6018
rect 17390 5966 17442 6018
rect 20526 5966 20578 6018
rect 20974 5966 21026 6018
rect 21310 5966 21362 6018
rect 22990 5966 23042 6018
rect 24670 5966 24722 6018
rect 25454 5966 25506 6018
rect 28702 5966 28754 6018
rect 28926 5966 28978 6018
rect 29822 5966 29874 6018
rect 30942 5966 30994 6018
rect 33406 5966 33458 6018
rect 2606 5854 2658 5906
rect 3054 5854 3106 5906
rect 3726 5854 3778 5906
rect 4398 5854 4450 5906
rect 4846 5854 4898 5906
rect 5294 5854 5346 5906
rect 6302 5854 6354 5906
rect 7422 5854 7474 5906
rect 7646 5854 7698 5906
rect 8206 5854 8258 5906
rect 8654 5854 8706 5906
rect 9998 5854 10050 5906
rect 10558 5854 10610 5906
rect 11454 5854 11506 5906
rect 13134 5854 13186 5906
rect 14590 5854 14642 5906
rect 15710 5854 15762 5906
rect 16158 5854 16210 5906
rect 18734 5854 18786 5906
rect 19294 5854 19346 5906
rect 20078 5854 20130 5906
rect 21422 5854 21474 5906
rect 21646 5854 21698 5906
rect 21758 5854 21810 5906
rect 22654 5854 22706 5906
rect 24222 5854 24274 5906
rect 25230 5854 25282 5906
rect 25566 5854 25618 5906
rect 26686 5854 26738 5906
rect 27470 5854 27522 5906
rect 30046 5854 30098 5906
rect 30494 5854 30546 5906
rect 31166 5854 31218 5906
rect 31614 5854 31666 5906
rect 31950 5854 32002 5906
rect 32958 5854 33010 5906
rect 33630 5854 33682 5906
rect 2158 5742 2210 5794
rect 6414 5742 6466 5794
rect 8990 5742 9042 5794
rect 10222 5742 10274 5794
rect 11902 5742 11954 5794
rect 16718 5742 16770 5794
rect 19406 5742 19458 5794
rect 19742 5742 19794 5794
rect 19854 5742 19906 5794
rect 22542 5742 22594 5794
rect 24334 5742 24386 5794
rect 26014 5742 26066 5794
rect 27582 5742 27634 5794
rect 31054 5742 31106 5794
rect 31726 5742 31778 5794
rect 33182 5742 33234 5794
rect 11566 5630 11618 5682
rect 26798 5630 26850 5682
rect 27022 5630 27074 5682
rect 27134 5630 27186 5682
rect 29038 5630 29090 5682
rect 32062 5630 32114 5682
rect 5372 5462 5424 5514
rect 5476 5462 5528 5514
rect 5580 5462 5632 5514
rect 13688 5462 13740 5514
rect 13792 5462 13844 5514
rect 13896 5462 13948 5514
rect 22004 5462 22056 5514
rect 22108 5462 22160 5514
rect 22212 5462 22264 5514
rect 30320 5462 30372 5514
rect 30424 5462 30476 5514
rect 30528 5462 30580 5514
rect 3950 5294 4002 5346
rect 4622 5294 4674 5346
rect 21982 5294 22034 5346
rect 27582 5294 27634 5346
rect 29262 5294 29314 5346
rect 2942 5182 2994 5234
rect 3390 5182 3442 5234
rect 11790 5182 11842 5234
rect 12126 5182 12178 5234
rect 19182 5182 19234 5234
rect 21646 5182 21698 5234
rect 24110 5182 24162 5234
rect 27806 5182 27858 5234
rect 32062 5182 32114 5234
rect 34190 5182 34242 5234
rect 2494 5070 2546 5122
rect 3614 5070 3666 5122
rect 4286 5070 4338 5122
rect 4846 5070 4898 5122
rect 5966 5070 6018 5122
rect 7422 5070 7474 5122
rect 8094 5070 8146 5122
rect 8878 5070 8930 5122
rect 9326 5070 9378 5122
rect 10110 5070 10162 5122
rect 10894 5070 10946 5122
rect 11230 5070 11282 5122
rect 12686 5070 12738 5122
rect 13470 5070 13522 5122
rect 13918 5070 13970 5122
rect 15934 5070 15986 5122
rect 18174 5070 18226 5122
rect 21870 5070 21922 5122
rect 22766 5070 22818 5122
rect 23326 5070 23378 5122
rect 27022 5070 27074 5122
rect 27358 5070 27410 5122
rect 29486 5070 29538 5122
rect 29710 5070 29762 5122
rect 30382 5070 30434 5122
rect 30494 5070 30546 5122
rect 30718 5070 30770 5122
rect 30942 5070 30994 5122
rect 31278 5070 31330 5122
rect 5070 4958 5122 5010
rect 6190 4958 6242 5010
rect 7310 4958 7362 5010
rect 7870 4958 7922 5010
rect 9886 4958 9938 5010
rect 10558 4958 10610 5010
rect 12462 4958 12514 5010
rect 14030 4958 14082 5010
rect 17726 4958 17778 5010
rect 21534 4958 21586 5010
rect 26238 4958 26290 5010
rect 4286 4846 4338 4898
rect 6302 4846 6354 4898
rect 7646 4846 7698 4898
rect 13582 4846 13634 4898
rect 15374 4846 15426 4898
rect 27470 4846 27522 4898
rect 29598 4846 29650 4898
rect 9530 4678 9582 4730
rect 9634 4678 9686 4730
rect 9738 4678 9790 4730
rect 17846 4678 17898 4730
rect 17950 4678 18002 4730
rect 18054 4678 18106 4730
rect 26162 4678 26214 4730
rect 26266 4678 26318 4730
rect 26370 4678 26422 4730
rect 34478 4678 34530 4730
rect 34582 4678 34634 4730
rect 34686 4678 34738 4730
rect 4734 4510 4786 4562
rect 6862 4510 6914 4562
rect 7646 4510 7698 4562
rect 7982 4510 8034 4562
rect 8990 4510 9042 4562
rect 11118 4510 11170 4562
rect 17278 4510 17330 4562
rect 19070 4510 19122 4562
rect 22766 4510 22818 4562
rect 33070 4510 33122 4562
rect 2494 4398 2546 4450
rect 6414 4398 6466 4450
rect 6974 4398 7026 4450
rect 10782 4398 10834 4450
rect 13358 4398 13410 4450
rect 27918 4398 27970 4450
rect 31166 4398 31218 4450
rect 1822 4286 1874 4338
rect 7422 4286 7474 4338
rect 8206 4286 8258 4338
rect 8766 4286 8818 4338
rect 11230 4286 11282 4338
rect 12126 4286 12178 4338
rect 12574 4286 12626 4338
rect 17614 4286 17666 4338
rect 18062 4286 18114 4338
rect 19518 4286 19570 4338
rect 23102 4286 23154 4338
rect 23774 4286 23826 4338
rect 24222 4286 24274 4338
rect 28702 4286 28754 4338
rect 31950 4286 32002 4338
rect 33406 4286 33458 4338
rect 33630 4286 33682 4338
rect 11790 4174 11842 4226
rect 15486 4174 15538 4226
rect 17726 4174 17778 4226
rect 20302 4174 20354 4226
rect 22430 4174 22482 4226
rect 23326 4174 23378 4226
rect 23662 4174 23714 4226
rect 25790 4174 25842 4226
rect 29038 4174 29090 4226
rect 5854 4062 5906 4114
rect 6862 4062 6914 4114
rect 10222 4062 10274 4114
rect 23998 4062 24050 4114
rect 5372 3894 5424 3946
rect 5476 3894 5528 3946
rect 5580 3894 5632 3946
rect 13688 3894 13740 3946
rect 13792 3894 13844 3946
rect 13896 3894 13948 3946
rect 22004 3894 22056 3946
rect 22108 3894 22160 3946
rect 22212 3894 22264 3946
rect 30320 3894 30372 3946
rect 30424 3894 30476 3946
rect 30528 3894 30580 3946
rect 7086 3726 7138 3778
rect 14142 3726 14194 3778
rect 14478 3726 14530 3778
rect 14926 3726 14978 3778
rect 15262 3726 15314 3778
rect 5742 3614 5794 3666
rect 8094 3614 8146 3666
rect 8430 3614 8482 3666
rect 10222 3614 10274 3666
rect 12350 3614 12402 3666
rect 13582 3614 13634 3666
rect 15486 3614 15538 3666
rect 16942 3614 16994 3666
rect 21534 3614 21586 3666
rect 23662 3614 23714 3666
rect 24558 3614 24610 3666
rect 24670 3614 24722 3666
rect 32958 3614 33010 3666
rect 6078 3502 6130 3554
rect 6750 3502 6802 3554
rect 6974 3502 7026 3554
rect 9550 3502 9602 3554
rect 14366 3502 14418 3554
rect 19742 3502 19794 3554
rect 20750 3502 20802 3554
rect 24894 3502 24946 3554
rect 25230 3502 25282 3554
rect 31502 3502 31554 3554
rect 32398 3502 32450 3554
rect 6302 3390 6354 3442
rect 6526 3390 6578 3442
rect 13246 3390 13298 3442
rect 19070 3390 19122 3442
rect 26910 3390 26962 3442
rect 30046 3390 30098 3442
rect 32174 3390 32226 3442
rect 9530 3110 9582 3162
rect 9634 3110 9686 3162
rect 9738 3110 9790 3162
rect 17846 3110 17898 3162
rect 17950 3110 18002 3162
rect 18054 3110 18106 3162
rect 26162 3110 26214 3162
rect 26266 3110 26318 3162
rect 26370 3110 26422 3162
rect 34478 3110 34530 3162
rect 34582 3110 34634 3162
rect 34686 3110 34738 3162
<< metal2 >>
rect 5370 32172 5634 32182
rect 5426 32116 5474 32172
rect 5530 32116 5578 32172
rect 5370 32106 5634 32116
rect 13686 32172 13950 32182
rect 13742 32116 13790 32172
rect 13846 32116 13894 32172
rect 13686 32106 13950 32116
rect 22002 32172 22266 32182
rect 22058 32116 22106 32172
rect 22162 32116 22210 32172
rect 22002 32106 22266 32116
rect 30318 32172 30582 32182
rect 30374 32116 30422 32172
rect 30478 32116 30526 32172
rect 30318 32106 30582 32116
rect 9528 31388 9792 31398
rect 9584 31332 9632 31388
rect 9688 31332 9736 31388
rect 9528 31322 9792 31332
rect 17844 31388 18108 31398
rect 17900 31332 17948 31388
rect 18004 31332 18052 31388
rect 17844 31322 18108 31332
rect 26160 31388 26424 31398
rect 26216 31332 26264 31388
rect 26320 31332 26368 31388
rect 26160 31322 26424 31332
rect 34476 31388 34740 31398
rect 34532 31332 34580 31388
rect 34636 31332 34684 31388
rect 34476 31322 34740 31332
rect 5370 30604 5634 30614
rect 5426 30548 5474 30604
rect 5530 30548 5578 30604
rect 5370 30538 5634 30548
rect 13686 30604 13950 30614
rect 13742 30548 13790 30604
rect 13846 30548 13894 30604
rect 13686 30538 13950 30548
rect 22002 30604 22266 30614
rect 22058 30548 22106 30604
rect 22162 30548 22210 30604
rect 22002 30538 22266 30548
rect 30318 30604 30582 30614
rect 30374 30548 30422 30604
rect 30478 30548 30526 30604
rect 30318 30538 30582 30548
rect 9528 29820 9792 29830
rect 9584 29764 9632 29820
rect 9688 29764 9736 29820
rect 9528 29754 9792 29764
rect 17844 29820 18108 29830
rect 17900 29764 17948 29820
rect 18004 29764 18052 29820
rect 17844 29754 18108 29764
rect 26160 29820 26424 29830
rect 26216 29764 26264 29820
rect 26320 29764 26368 29820
rect 26160 29754 26424 29764
rect 34476 29820 34740 29830
rect 34532 29764 34580 29820
rect 34636 29764 34684 29820
rect 34476 29754 34740 29764
rect 5370 29036 5634 29046
rect 5426 28980 5474 29036
rect 5530 28980 5578 29036
rect 5370 28970 5634 28980
rect 13686 29036 13950 29046
rect 13742 28980 13790 29036
rect 13846 28980 13894 29036
rect 13686 28970 13950 28980
rect 22002 29036 22266 29046
rect 22058 28980 22106 29036
rect 22162 28980 22210 29036
rect 22002 28970 22266 28980
rect 30318 29036 30582 29046
rect 30374 28980 30422 29036
rect 30478 28980 30526 29036
rect 30318 28970 30582 28980
rect 11228 28756 11284 28766
rect 11228 28754 11732 28756
rect 11228 28702 11230 28754
rect 11282 28702 11732 28754
rect 11228 28700 11732 28702
rect 11228 28690 11284 28700
rect 8428 28642 8484 28654
rect 8428 28590 8430 28642
rect 8482 28590 8484 28642
rect 5068 27970 5124 27982
rect 5068 27918 5070 27970
rect 5122 27918 5124 27970
rect 4284 27858 4340 27870
rect 4284 27806 4286 27858
rect 4338 27806 4340 27858
rect 3612 27748 3668 27758
rect 2940 27746 3668 27748
rect 2940 27694 3614 27746
rect 3666 27694 3668 27746
rect 2940 27692 3668 27694
rect 1820 27074 1876 27086
rect 1820 27022 1822 27074
rect 1874 27022 1876 27074
rect 1820 26290 1876 27022
rect 2492 26962 2548 26974
rect 2492 26910 2494 26962
rect 2546 26910 2548 26962
rect 2492 26404 2548 26910
rect 2492 26338 2548 26348
rect 1820 26238 1822 26290
rect 1874 26238 1876 26290
rect 1820 25508 1876 26238
rect 2492 26180 2548 26190
rect 2492 26178 2660 26180
rect 2492 26126 2494 26178
rect 2546 26126 2660 26178
rect 2492 26124 2660 26126
rect 2492 26114 2548 26124
rect 2604 25730 2660 26124
rect 2604 25678 2606 25730
rect 2658 25678 2660 25730
rect 2604 25666 2660 25678
rect 2940 25730 2996 27692
rect 3612 27682 3668 27692
rect 4284 26908 4340 27806
rect 4508 27860 4564 27870
rect 4844 27860 4900 27870
rect 4508 27858 4900 27860
rect 4508 27806 4510 27858
rect 4562 27806 4846 27858
rect 4898 27806 4900 27858
rect 4508 27804 4900 27806
rect 4508 27794 4564 27804
rect 4844 27794 4900 27804
rect 4620 27188 4676 27198
rect 4956 27188 5012 27198
rect 5068 27188 5124 27918
rect 5180 27858 5236 27870
rect 5180 27806 5182 27858
rect 5234 27806 5236 27858
rect 5180 27300 5236 27806
rect 8428 27860 8484 28590
rect 9100 28532 9156 28542
rect 9100 28530 9940 28532
rect 9100 28478 9102 28530
rect 9154 28478 9940 28530
rect 9100 28476 9940 28478
rect 9100 28466 9156 28476
rect 9528 28252 9792 28262
rect 9584 28196 9632 28252
rect 9688 28196 9736 28252
rect 9528 28186 9792 28196
rect 5370 27468 5634 27478
rect 5426 27412 5474 27468
rect 5530 27412 5578 27468
rect 5370 27402 5634 27412
rect 5180 27234 5236 27244
rect 5852 27300 5908 27310
rect 5852 27206 5908 27244
rect 4620 27186 5124 27188
rect 4620 27134 4622 27186
rect 4674 27134 4958 27186
rect 5010 27134 5124 27186
rect 4620 27132 5124 27134
rect 4620 27122 4676 27132
rect 4956 27122 5012 27132
rect 5964 27076 6020 27086
rect 5964 26982 6020 27020
rect 6188 27074 6244 27086
rect 6188 27022 6190 27074
rect 6242 27022 6244 27074
rect 4956 26964 5012 26974
rect 4284 26852 4564 26908
rect 2940 25678 2942 25730
rect 2994 25678 2996 25730
rect 2940 25666 2996 25678
rect 3276 26404 3332 26414
rect 3276 25730 3332 26348
rect 3276 25678 3278 25730
rect 3330 25678 3332 25730
rect 3276 25666 3332 25678
rect 4508 26180 4564 26852
rect 4620 26180 4676 26190
rect 4508 26178 4676 26180
rect 4508 26126 4622 26178
rect 4674 26126 4676 26178
rect 4508 26124 4676 26126
rect 1820 23156 1876 25452
rect 2604 25508 2660 25518
rect 3276 25508 3332 25518
rect 2604 25506 3332 25508
rect 2604 25454 2606 25506
rect 2658 25454 3278 25506
rect 3330 25454 3332 25506
rect 2604 25452 3332 25454
rect 1820 23154 1988 23156
rect 1820 23102 1822 23154
rect 1874 23102 1988 23154
rect 1820 23100 1988 23102
rect 1820 23090 1876 23100
rect 1932 22370 1988 23100
rect 2492 23042 2548 23054
rect 2492 22990 2494 23042
rect 2546 22990 2548 23042
rect 2492 22596 2548 22990
rect 2492 22530 2548 22540
rect 1932 22318 1934 22370
rect 1986 22318 1988 22370
rect 1820 20020 1876 20030
rect 1932 20020 1988 22318
rect 2604 21026 2660 25452
rect 3276 24948 3332 25452
rect 3612 25396 3668 25406
rect 4060 25396 4116 25406
rect 3612 25394 4116 25396
rect 3612 25342 3614 25394
rect 3666 25342 4062 25394
rect 4114 25342 4116 25394
rect 3612 25340 4116 25342
rect 3612 25330 3668 25340
rect 4060 25330 4116 25340
rect 3276 24882 3332 24892
rect 4060 24836 4116 24846
rect 4060 24742 4116 24780
rect 4396 24722 4452 24734
rect 4396 24670 4398 24722
rect 4450 24670 4452 24722
rect 4396 24164 4452 24670
rect 4508 24724 4564 26124
rect 4620 26114 4676 26124
rect 4956 25620 5012 26908
rect 4732 25618 5012 25620
rect 4732 25566 4958 25618
rect 5010 25566 5012 25618
rect 4732 25564 5012 25566
rect 4620 25506 4676 25518
rect 4620 25454 4622 25506
rect 4674 25454 4676 25506
rect 4620 25396 4676 25454
rect 4620 25330 4676 25340
rect 4732 24946 4788 25564
rect 4956 25554 5012 25564
rect 5068 26962 5124 26974
rect 5068 26910 5070 26962
rect 5122 26910 5124 26962
rect 5068 25396 5124 26910
rect 5068 25330 5124 25340
rect 5180 26964 5236 26974
rect 5180 26178 5236 26908
rect 5180 26126 5182 26178
rect 5234 26126 5236 26178
rect 4732 24894 4734 24946
rect 4786 24894 4788 24946
rect 4732 24882 4788 24894
rect 5068 24948 5124 24958
rect 4620 24724 4676 24734
rect 4508 24668 4620 24724
rect 4620 24658 4676 24668
rect 5068 24722 5124 24892
rect 5068 24670 5070 24722
rect 5122 24670 5124 24722
rect 5068 24164 5124 24670
rect 5180 24724 5236 26126
rect 5370 25900 5634 25910
rect 5426 25844 5474 25900
rect 5530 25844 5578 25900
rect 5370 25834 5634 25844
rect 5852 25396 5908 25406
rect 5740 24836 5796 24846
rect 5292 24724 5348 24734
rect 5180 24722 5348 24724
rect 5180 24670 5294 24722
rect 5346 24670 5348 24722
rect 5180 24668 5348 24670
rect 5292 24658 5348 24668
rect 5628 24724 5684 24734
rect 5628 24630 5684 24668
rect 5370 24332 5634 24342
rect 5426 24276 5474 24332
rect 5530 24276 5578 24332
rect 5370 24266 5634 24276
rect 5068 24108 5572 24164
rect 4396 24098 4452 24108
rect 5068 23828 5124 23838
rect 5068 23826 5236 23828
rect 5068 23774 5070 23826
rect 5122 23774 5236 23826
rect 5068 23772 5236 23774
rect 5068 23762 5124 23772
rect 4844 23714 4900 23726
rect 4844 23662 4846 23714
rect 4898 23662 4900 23714
rect 4620 23042 4676 23054
rect 4620 22990 4622 23042
rect 4674 22990 4676 23042
rect 2716 22932 2772 22942
rect 2716 22482 2772 22876
rect 2716 22430 2718 22482
rect 2770 22430 2772 22482
rect 2716 22418 2772 22430
rect 3612 22372 3668 22382
rect 3612 21810 3668 22316
rect 3612 21758 3614 21810
rect 3666 21758 3668 21810
rect 3612 21746 3668 21758
rect 3948 21700 4004 21710
rect 3948 21606 4004 21644
rect 4620 21700 4676 22990
rect 4844 23044 4900 23662
rect 4956 23714 5012 23726
rect 4956 23662 4958 23714
rect 5010 23662 5012 23714
rect 4956 23268 5012 23662
rect 4956 23202 5012 23212
rect 5180 23156 5236 23772
rect 5516 23378 5572 24108
rect 5516 23326 5518 23378
rect 5570 23326 5572 23378
rect 5516 23314 5572 23326
rect 5068 23154 5236 23156
rect 5068 23102 5182 23154
rect 5234 23102 5236 23154
rect 5068 23100 5236 23102
rect 4956 23044 5012 23054
rect 4844 23042 5012 23044
rect 4844 22990 4958 23042
rect 5010 22990 5012 23042
rect 4844 22988 5012 22990
rect 4844 22482 4900 22988
rect 4956 22978 5012 22988
rect 4844 22430 4846 22482
rect 4898 22430 4900 22482
rect 4844 21812 4900 22430
rect 4844 21746 4900 21756
rect 5068 22148 5124 23100
rect 5180 23090 5236 23100
rect 5370 22764 5634 22774
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5370 22698 5634 22708
rect 5628 22596 5684 22606
rect 5628 22502 5684 22540
rect 5740 22594 5796 24780
rect 5852 24834 5908 25340
rect 6188 25172 6244 27022
rect 6748 27076 6804 27086
rect 6748 26982 6804 27020
rect 7420 27074 7476 27086
rect 7420 27022 7422 27074
rect 7474 27022 7476 27074
rect 6300 26962 6356 26974
rect 6300 26910 6302 26962
rect 6354 26910 6356 26962
rect 6300 26404 6356 26910
rect 6300 26338 6356 26348
rect 6412 26964 6468 26974
rect 6188 25116 6356 25172
rect 5852 24782 5854 24834
rect 5906 24782 5908 24834
rect 5852 24770 5908 24782
rect 6076 24948 6132 24958
rect 5852 23268 5908 23278
rect 5852 23154 5908 23212
rect 5852 23102 5854 23154
rect 5906 23102 5908 23154
rect 5852 23090 5908 23102
rect 6076 23154 6132 24892
rect 6076 23102 6078 23154
rect 6130 23102 6132 23154
rect 6076 23090 6132 23102
rect 6188 24946 6244 24958
rect 6188 24894 6190 24946
rect 6242 24894 6244 24946
rect 5740 22542 5742 22594
rect 5794 22542 5796 22594
rect 5740 22530 5796 22542
rect 5964 22370 6020 22382
rect 5964 22318 5966 22370
rect 6018 22318 6020 22370
rect 5964 22148 6020 22318
rect 6076 22372 6132 22382
rect 6076 22278 6132 22316
rect 5068 22092 6020 22148
rect 5068 21810 5124 22092
rect 5068 21758 5070 21810
rect 5122 21758 5124 21810
rect 5068 21746 5124 21758
rect 5516 21812 5572 21822
rect 5516 21718 5572 21756
rect 4620 21606 4676 21644
rect 5404 21700 5460 21710
rect 5404 21606 5460 21644
rect 2604 20974 2606 21026
rect 2658 20974 2660 21026
rect 2604 20962 2660 20974
rect 3388 21586 3444 21598
rect 3388 21534 3390 21586
rect 3442 21534 3444 21586
rect 3276 20804 3332 20814
rect 3276 20710 3332 20748
rect 2380 20580 2436 20590
rect 2380 20486 2436 20524
rect 2492 20578 2548 20590
rect 2492 20526 2494 20578
rect 2546 20526 2548 20578
rect 2492 20130 2548 20526
rect 2940 20580 2996 20590
rect 2940 20486 2996 20524
rect 3388 20580 3444 21534
rect 3388 20514 3444 20524
rect 3612 21586 3668 21598
rect 3612 21534 3614 21586
rect 3666 21534 3668 21586
rect 3612 20578 3668 21534
rect 4396 21586 4452 21598
rect 4396 21534 4398 21586
rect 4450 21534 4452 21586
rect 4396 20916 4452 21534
rect 4508 21586 4564 21598
rect 4508 21534 4510 21586
rect 4562 21534 4564 21586
rect 4508 21028 4564 21534
rect 5740 21586 5796 21598
rect 5740 21534 5742 21586
rect 5794 21534 5796 21586
rect 5370 21196 5634 21206
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5370 21130 5634 21140
rect 4508 20972 4788 21028
rect 4396 20860 4564 20916
rect 4284 20804 4340 20814
rect 4172 20748 4284 20804
rect 3948 20692 4004 20702
rect 3948 20598 4004 20636
rect 3612 20526 3614 20578
rect 3666 20526 3668 20578
rect 2492 20078 2494 20130
rect 2546 20078 2548 20130
rect 2492 20066 2548 20078
rect 1820 20018 1988 20020
rect 1820 19966 1822 20018
rect 1874 19966 1988 20018
rect 1820 19964 1988 19966
rect 3612 20020 3668 20526
rect 1820 19234 1876 19964
rect 3612 19954 3668 19964
rect 2492 19908 2548 19918
rect 2492 19346 2548 19852
rect 4172 19796 4228 20748
rect 4284 20738 4340 20748
rect 4284 20580 4340 20590
rect 4284 20486 4340 20524
rect 4396 20578 4452 20590
rect 4396 20526 4398 20578
rect 4450 20526 4452 20578
rect 4396 20132 4452 20526
rect 4396 20066 4452 20076
rect 4508 20578 4564 20860
rect 4732 20804 4788 20972
rect 4732 20738 4788 20748
rect 4956 20802 5012 20814
rect 4956 20750 4958 20802
rect 5010 20750 5012 20802
rect 4508 20526 4510 20578
rect 4562 20526 4564 20578
rect 4508 20020 4564 20526
rect 4620 20692 4676 20702
rect 4620 20132 4676 20636
rect 4844 20580 4900 20590
rect 4620 20076 4788 20132
rect 4508 19954 4564 19964
rect 4620 19906 4676 19918
rect 4620 19854 4622 19906
rect 4674 19854 4676 19906
rect 4620 19796 4676 19854
rect 4172 19740 4676 19796
rect 2492 19294 2494 19346
rect 2546 19294 2548 19346
rect 2492 19282 2548 19294
rect 4620 19348 4676 19358
rect 4732 19348 4788 20076
rect 4844 20018 4900 20524
rect 4956 20244 5012 20750
rect 5628 20802 5684 20814
rect 5628 20750 5630 20802
rect 5682 20750 5684 20802
rect 5628 20468 5684 20750
rect 5740 20690 5796 21534
rect 5740 20638 5742 20690
rect 5794 20638 5796 20690
rect 5740 20626 5796 20638
rect 6188 20468 6244 24894
rect 6300 24164 6356 25116
rect 6412 24834 6468 26908
rect 6636 26962 6692 26974
rect 6636 26910 6638 26962
rect 6690 26910 6692 26962
rect 6636 24948 6692 26910
rect 6860 26964 6916 26974
rect 6860 26870 6916 26908
rect 7308 26404 7364 26414
rect 7308 26310 7364 26348
rect 6636 24882 6692 24892
rect 7084 25508 7140 25518
rect 6412 24782 6414 24834
rect 6466 24782 6468 24834
rect 6412 24770 6468 24782
rect 6300 22930 6356 24108
rect 7084 23938 7140 25452
rect 7420 25508 7476 27022
rect 8204 26962 8260 26974
rect 8428 26964 8484 27804
rect 8204 26910 8206 26962
rect 8258 26910 8260 26962
rect 8204 26516 8260 26910
rect 8204 26450 8260 26460
rect 8316 26908 8484 26964
rect 7420 25442 7476 25452
rect 7980 26292 8036 26302
rect 8316 26292 8372 26908
rect 9528 26684 9792 26694
rect 9584 26628 9632 26684
rect 9688 26628 9736 26684
rect 9528 26618 9792 26628
rect 7980 26290 8372 26292
rect 7980 26238 7982 26290
rect 8034 26238 8372 26290
rect 7980 26236 8372 26238
rect 8876 26516 8932 26526
rect 7980 25508 8036 26236
rect 7980 25442 8036 25452
rect 7756 25394 7812 25406
rect 7756 25342 7758 25394
rect 7810 25342 7812 25394
rect 7756 24164 7812 25342
rect 8876 24946 8932 26460
rect 9884 26514 9940 28476
rect 10220 27860 10276 27870
rect 10220 27766 10276 27804
rect 11004 27748 11060 27758
rect 11004 27654 11060 27692
rect 9884 26462 9886 26514
rect 9938 26462 9940 26514
rect 9884 26450 9940 26462
rect 10332 27186 10388 27198
rect 10332 27134 10334 27186
rect 10386 27134 10388 27186
rect 9996 26178 10052 26190
rect 9996 26126 9998 26178
rect 10050 26126 10052 26178
rect 9884 25618 9940 25630
rect 9884 25566 9886 25618
rect 9938 25566 9940 25618
rect 9528 25116 9792 25126
rect 9584 25060 9632 25116
rect 9688 25060 9736 25116
rect 9528 25050 9792 25060
rect 8876 24894 8878 24946
rect 8930 24894 8932 24946
rect 8876 24882 8932 24894
rect 8988 24610 9044 24622
rect 8988 24558 8990 24610
rect 9042 24558 9044 24610
rect 7756 24098 7812 24108
rect 8764 24164 8820 24174
rect 7084 23886 7086 23938
rect 7138 23886 7140 23938
rect 6300 22878 6302 22930
rect 6354 22878 6356 22930
rect 6300 22596 6356 22878
rect 6412 22932 6468 22942
rect 6412 22838 6468 22876
rect 6300 22530 6356 22540
rect 7084 22484 7140 23886
rect 7868 23828 7924 23838
rect 7868 23826 8372 23828
rect 7868 23774 7870 23826
rect 7922 23774 8372 23826
rect 7868 23772 8372 23774
rect 7868 23762 7924 23772
rect 8316 23378 8372 23772
rect 8316 23326 8318 23378
rect 8370 23326 8372 23378
rect 8316 23314 8372 23326
rect 8764 23378 8820 24108
rect 8988 24052 9044 24558
rect 8988 23986 9044 23996
rect 9528 23548 9792 23558
rect 9584 23492 9632 23548
rect 9688 23492 9736 23548
rect 9528 23482 9792 23492
rect 8764 23326 8766 23378
rect 8818 23326 8820 23378
rect 8764 23314 8820 23326
rect 9884 23268 9940 25566
rect 9996 24948 10052 26126
rect 9996 24882 10052 24892
rect 10332 24612 10388 27134
rect 11676 26964 11732 28700
rect 17844 28252 18108 28262
rect 17900 28196 17948 28252
rect 18004 28196 18052 28252
rect 17844 28186 18108 28196
rect 26160 28252 26424 28262
rect 26216 28196 26264 28252
rect 26320 28196 26368 28252
rect 26160 28186 26424 28196
rect 34476 28252 34740 28262
rect 34532 28196 34580 28252
rect 34636 28196 34684 28252
rect 34476 28186 34740 28196
rect 20300 28082 20356 28094
rect 20300 28030 20302 28082
rect 20354 28030 20356 28082
rect 19068 27860 19124 27870
rect 12236 27748 12292 27758
rect 12236 27186 12292 27692
rect 12236 27134 12238 27186
rect 12290 27134 12292 27186
rect 12236 27122 12292 27134
rect 13132 27746 13188 27758
rect 13132 27694 13134 27746
rect 13186 27694 13188 27746
rect 12460 27076 12516 27086
rect 12460 26982 12516 27020
rect 11676 26908 11844 26964
rect 11788 26290 11844 26908
rect 11788 26238 11790 26290
rect 11842 26238 11844 26290
rect 11004 25732 11060 25742
rect 11004 24948 11060 25676
rect 11788 25172 11844 26238
rect 12124 26962 12180 26974
rect 12124 26910 12126 26962
rect 12178 26910 12180 26962
rect 12012 25508 12068 25518
rect 12012 25414 12068 25452
rect 11228 25116 11844 25172
rect 10332 24546 10388 24556
rect 10892 24946 11060 24948
rect 10892 24894 11006 24946
rect 11058 24894 11060 24946
rect 10892 24892 11060 24894
rect 9996 24164 10052 24174
rect 9996 24050 10052 24108
rect 9996 23998 9998 24050
rect 10050 23998 10052 24050
rect 9996 23986 10052 23998
rect 10780 23940 10836 23950
rect 9996 23380 10052 23390
rect 9996 23286 10052 23324
rect 9884 23174 9940 23212
rect 10220 23266 10276 23278
rect 10220 23214 10222 23266
rect 10274 23214 10276 23266
rect 10220 23156 10276 23214
rect 10332 23156 10388 23166
rect 10220 23154 10388 23156
rect 10220 23102 10334 23154
rect 10386 23102 10388 23154
rect 10220 23100 10388 23102
rect 10332 23090 10388 23100
rect 10668 23154 10724 23166
rect 10668 23102 10670 23154
rect 10722 23102 10724 23154
rect 8428 23042 8484 23054
rect 8428 22990 8430 23042
rect 8482 22990 8484 23042
rect 7084 22418 7140 22428
rect 7868 22484 7924 22494
rect 7868 22390 7924 22428
rect 8428 22260 8484 22990
rect 8876 23044 8932 23054
rect 8876 22950 8932 22988
rect 8428 22194 8484 22204
rect 9528 21980 9792 21990
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9528 21914 9792 21924
rect 10332 21588 10388 21598
rect 7644 20804 7700 20814
rect 7644 20710 7700 20748
rect 8204 20692 8260 20702
rect 8204 20598 8260 20636
rect 5628 20412 6244 20468
rect 8092 20578 8148 20590
rect 8092 20526 8094 20578
rect 8146 20526 8148 20578
rect 4956 20178 5012 20188
rect 5404 20132 5460 20142
rect 4844 19966 4846 20018
rect 4898 19966 4900 20018
rect 4844 19954 4900 19966
rect 5180 20020 5236 20030
rect 5180 19926 5236 19964
rect 5404 20018 5460 20076
rect 5404 19966 5406 20018
rect 5458 19966 5460 20018
rect 5404 19954 5460 19966
rect 7308 20020 7364 20030
rect 5068 19908 5124 19918
rect 7308 19908 7364 19964
rect 5068 19814 5124 19852
rect 7196 19906 7364 19908
rect 7196 19854 7310 19906
rect 7362 19854 7364 19906
rect 7196 19852 7364 19854
rect 5370 19628 5634 19638
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5370 19562 5634 19572
rect 4620 19346 4788 19348
rect 4620 19294 4622 19346
rect 4674 19294 4788 19346
rect 4620 19292 4788 19294
rect 4620 19282 4676 19292
rect 1820 19182 1822 19234
rect 1874 19182 1876 19234
rect 1820 19170 1876 19182
rect 7084 19234 7140 19246
rect 7084 19182 7086 19234
rect 7138 19182 7140 19234
rect 6972 18788 7028 18798
rect 6524 18564 6580 18574
rect 6748 18564 6804 18574
rect 6524 18562 6748 18564
rect 6524 18510 6526 18562
rect 6578 18510 6748 18562
rect 6524 18508 6748 18510
rect 6524 18498 6580 18508
rect 6748 18498 6804 18508
rect 6300 18450 6356 18462
rect 6300 18398 6302 18450
rect 6354 18398 6356 18450
rect 6300 18340 6356 18398
rect 6860 18340 6916 18350
rect 6300 18338 6916 18340
rect 6300 18286 6862 18338
rect 6914 18286 6916 18338
rect 6300 18284 6916 18286
rect 5370 18060 5634 18070
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5370 17994 5634 18004
rect 4620 17778 4676 17790
rect 4620 17726 4622 17778
rect 4674 17726 4676 17778
rect 1820 17666 1876 17678
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1596 15204 1652 15214
rect 1596 4228 1652 15148
rect 1820 15092 1876 17614
rect 4620 17668 4676 17726
rect 4620 17602 4676 17612
rect 5740 17668 5796 17678
rect 5740 17574 5796 17612
rect 6300 17666 6356 17678
rect 6300 17614 6302 17666
rect 6354 17614 6356 17666
rect 2492 17556 2548 17566
rect 2380 17554 2548 17556
rect 2380 17502 2494 17554
rect 2546 17502 2548 17554
rect 2380 17500 2548 17502
rect 1820 14530 1876 15036
rect 2268 16098 2324 16110
rect 2268 16046 2270 16098
rect 2322 16046 2324 16098
rect 2268 15092 2324 16046
rect 2268 15026 2324 15036
rect 1820 14478 1822 14530
rect 1874 14478 1876 14530
rect 1820 14466 1876 14478
rect 2380 11506 2436 17500
rect 2492 17490 2548 17500
rect 5964 17556 6020 17566
rect 5964 17462 6020 17500
rect 5068 17444 5124 17454
rect 5068 17442 5236 17444
rect 5068 17390 5070 17442
rect 5122 17390 5236 17442
rect 5068 17388 5236 17390
rect 5068 17378 5124 17388
rect 5068 16996 5124 17006
rect 3276 16882 3332 16894
rect 3276 16830 3278 16882
rect 3330 16830 3332 16882
rect 2940 15986 2996 15998
rect 2940 15934 2942 15986
rect 2994 15934 2996 15986
rect 2492 14418 2548 14430
rect 2492 14366 2494 14418
rect 2546 14366 2548 14418
rect 2492 11620 2548 14366
rect 2940 14308 2996 15934
rect 3276 15092 3332 16830
rect 3948 16884 4004 16894
rect 3948 16790 4004 16828
rect 5068 16210 5124 16940
rect 5068 16158 5070 16210
rect 5122 16158 5124 16210
rect 5068 16146 5124 16158
rect 5180 15148 5236 17388
rect 5852 16884 5908 16894
rect 5370 16492 5634 16502
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5370 16426 5634 16436
rect 3276 15026 3332 15036
rect 5068 15092 5236 15148
rect 5740 15874 5796 15886
rect 5740 15822 5742 15874
rect 5794 15822 5796 15874
rect 5740 15314 5796 15822
rect 5740 15262 5742 15314
rect 5794 15262 5796 15314
rect 5740 15092 5796 15262
rect 5852 15148 5908 16828
rect 6300 16884 6356 17614
rect 6524 17668 6580 17678
rect 6524 17574 6580 17612
rect 6748 16996 6804 18284
rect 6860 18274 6916 18284
rect 6860 17892 6916 17902
rect 6860 17798 6916 17836
rect 6972 17108 7028 18732
rect 7084 18226 7140 19182
rect 7084 18174 7086 18226
rect 7138 18174 7140 18226
rect 7084 17556 7140 18174
rect 7196 17892 7252 19852
rect 7308 19842 7364 19852
rect 7756 20018 7812 20030
rect 7756 19966 7758 20018
rect 7810 19966 7812 20018
rect 7532 19236 7588 19246
rect 7756 19236 7812 19966
rect 7980 19908 8036 19918
rect 7980 19346 8036 19852
rect 7980 19294 7982 19346
rect 8034 19294 8036 19346
rect 7980 19282 8036 19294
rect 7532 19234 7812 19236
rect 7532 19182 7534 19234
rect 7586 19182 7812 19234
rect 7532 19180 7812 19182
rect 7532 19170 7588 19180
rect 7420 18676 7476 18686
rect 7420 18582 7476 18620
rect 7196 17826 7252 17836
rect 7756 18564 7812 19180
rect 7644 17668 7700 17678
rect 7644 17574 7700 17612
rect 7084 17490 7140 17500
rect 7196 17554 7252 17566
rect 7196 17502 7198 17554
rect 7250 17502 7252 17554
rect 7084 17108 7140 17118
rect 6972 17106 7140 17108
rect 6972 17054 7086 17106
rect 7138 17054 7140 17106
rect 6972 17052 7140 17054
rect 7084 17042 7140 17052
rect 6748 16902 6804 16940
rect 7196 16996 7252 17502
rect 7308 17444 7364 17454
rect 7308 17442 7700 17444
rect 7308 17390 7310 17442
rect 7362 17390 7700 17442
rect 7308 17388 7700 17390
rect 7308 17378 7364 17388
rect 7644 17106 7700 17388
rect 7644 17054 7646 17106
rect 7698 17054 7700 17106
rect 7644 17042 7700 17054
rect 7756 17108 7812 18508
rect 7980 18564 8036 18574
rect 7980 18470 8036 18508
rect 7756 17042 7812 17052
rect 7868 18450 7924 18462
rect 7868 18398 7870 18450
rect 7922 18398 7924 18450
rect 7868 17666 7924 18398
rect 7868 17614 7870 17666
rect 7922 17614 7924 17666
rect 7196 16930 7252 16940
rect 6076 16772 6132 16782
rect 6300 16772 6356 16828
rect 7532 16884 7588 16894
rect 7868 16884 7924 17614
rect 8092 17668 8148 20526
rect 9884 20580 9940 20590
rect 9528 20412 9792 20422
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9528 20346 9792 20356
rect 8204 20132 8260 20142
rect 8204 20038 8260 20076
rect 8876 20130 8932 20142
rect 8876 20078 8878 20130
rect 8930 20078 8932 20130
rect 8876 20020 8932 20078
rect 8876 19954 8932 19964
rect 9436 20020 9492 20030
rect 9772 20020 9828 20030
rect 9884 20020 9940 20524
rect 10220 20578 10276 20590
rect 10220 20526 10222 20578
rect 10274 20526 10276 20578
rect 9492 19964 9604 20020
rect 9436 19954 9492 19964
rect 8652 19794 8708 19806
rect 8652 19742 8654 19794
rect 8706 19742 8708 19794
rect 8652 19236 8708 19742
rect 8988 19796 9044 19806
rect 8988 19794 9156 19796
rect 8988 19742 8990 19794
rect 9042 19742 9156 19794
rect 8988 19740 9156 19742
rect 8988 19730 9044 19740
rect 8988 19348 9044 19358
rect 8988 19254 9044 19292
rect 8428 19234 8708 19236
rect 8428 19182 8654 19234
rect 8706 19182 8708 19234
rect 8428 19180 8708 19182
rect 8204 18788 8260 18798
rect 8204 18674 8260 18732
rect 8204 18622 8206 18674
rect 8258 18622 8260 18674
rect 8204 18610 8260 18622
rect 8316 18450 8372 18462
rect 8316 18398 8318 18450
rect 8370 18398 8372 18450
rect 8204 18338 8260 18350
rect 8204 18286 8206 18338
rect 8258 18286 8260 18338
rect 8204 18116 8260 18286
rect 8204 18050 8260 18060
rect 8316 17668 8372 18398
rect 8092 17612 8260 17668
rect 8092 17332 8148 17342
rect 8204 17332 8260 17612
rect 8316 17602 8372 17612
rect 8428 17892 8484 19180
rect 8652 19170 8708 19180
rect 8876 19234 8932 19246
rect 8876 19182 8878 19234
rect 8930 19182 8932 19234
rect 8876 19124 8932 19182
rect 9100 19124 9156 19740
rect 9548 19460 9604 19964
rect 9772 20018 9940 20020
rect 9772 19966 9774 20018
rect 9826 19966 9940 20018
rect 9772 19964 9940 19966
rect 9996 20244 10052 20254
rect 9996 20020 10052 20188
rect 10220 20132 10276 20526
rect 10332 20356 10388 21532
rect 10556 21586 10612 21598
rect 10556 21534 10558 21586
rect 10610 21534 10612 21586
rect 10556 20690 10612 21534
rect 10668 21476 10724 23102
rect 10780 23042 10836 23884
rect 10892 23938 10948 24892
rect 11004 24882 11060 24892
rect 11116 24948 11172 24958
rect 11116 24854 11172 24892
rect 11228 24946 11284 25116
rect 11228 24894 11230 24946
rect 11282 24894 11284 24946
rect 11228 24882 11284 24894
rect 11340 24834 11396 24846
rect 11340 24782 11342 24834
rect 11394 24782 11396 24834
rect 11116 24612 11172 24622
rect 11004 24052 11060 24062
rect 11004 23958 11060 23996
rect 10892 23886 10894 23938
rect 10946 23886 10948 23938
rect 10892 23874 10948 23886
rect 11116 23828 11172 24556
rect 11116 23734 11172 23772
rect 11228 23940 11284 23950
rect 11228 23826 11284 23884
rect 11228 23774 11230 23826
rect 11282 23774 11284 23826
rect 11228 23762 11284 23774
rect 10780 22990 10782 23042
rect 10834 22990 10836 23042
rect 10780 22978 10836 22990
rect 10892 23266 10948 23278
rect 10892 23214 10894 23266
rect 10946 23214 10948 23266
rect 10892 22932 10948 23214
rect 11340 23156 11396 24782
rect 11788 24836 11844 25116
rect 12124 24948 12180 26910
rect 12684 26962 12740 26974
rect 12684 26910 12686 26962
rect 12738 26910 12740 26962
rect 12348 26292 12404 26302
rect 12348 26198 12404 26236
rect 12460 26178 12516 26190
rect 12460 26126 12462 26178
rect 12514 26126 12516 26178
rect 12460 25508 12516 26126
rect 12684 25620 12740 26910
rect 13132 26292 13188 27694
rect 13686 27468 13950 27478
rect 13742 27412 13790 27468
rect 13846 27412 13894 27468
rect 13686 27402 13950 27412
rect 16380 27188 16436 27198
rect 14364 27074 14420 27086
rect 14364 27022 14366 27074
rect 14418 27022 14420 27074
rect 14364 26964 14420 27022
rect 14364 26898 14420 26908
rect 15036 26962 15092 26974
rect 15036 26910 15038 26962
rect 15090 26910 15092 26962
rect 15036 26404 15092 26910
rect 15484 26964 15540 26974
rect 15484 26852 15652 26908
rect 15596 26516 15652 26852
rect 16268 26516 16324 26526
rect 15596 26460 15876 26516
rect 15036 26348 15428 26404
rect 12684 25554 12740 25564
rect 12908 26178 12964 26190
rect 12908 26126 12910 26178
rect 12962 26126 12964 26178
rect 12572 25508 12628 25518
rect 12460 25506 12628 25508
rect 12460 25454 12574 25506
rect 12626 25454 12628 25506
rect 12460 25452 12628 25454
rect 12572 25442 12628 25452
rect 12348 25396 12404 25406
rect 12348 25302 12404 25340
rect 12908 25396 12964 26126
rect 13132 25508 13188 26236
rect 15036 26180 15092 26190
rect 14476 26178 15092 26180
rect 14476 26126 15038 26178
rect 15090 26126 15092 26178
rect 14476 26124 15092 26126
rect 13686 25900 13950 25910
rect 13742 25844 13790 25900
rect 13846 25844 13894 25900
rect 13686 25834 13950 25844
rect 14140 25844 14196 25854
rect 13580 25620 13636 25630
rect 13580 25526 13636 25564
rect 13132 25442 13188 25452
rect 13692 25508 13748 25518
rect 12908 25330 12964 25340
rect 12460 25284 12516 25294
rect 12460 25190 12516 25228
rect 13468 25282 13524 25294
rect 13468 25230 13470 25282
rect 13522 25230 13524 25282
rect 13468 25172 13524 25230
rect 13356 25116 13524 25172
rect 13356 25060 13412 25116
rect 13692 25060 13748 25452
rect 14140 25506 14196 25788
rect 14476 25618 14532 26124
rect 15036 26114 15092 26124
rect 14476 25566 14478 25618
rect 14530 25566 14532 25618
rect 14476 25554 14532 25566
rect 15372 25618 15428 26348
rect 15372 25566 15374 25618
rect 15426 25566 15428 25618
rect 15372 25554 15428 25566
rect 14140 25454 14142 25506
rect 14194 25454 14196 25506
rect 14140 25442 14196 25454
rect 14252 25506 14308 25518
rect 14252 25454 14254 25506
rect 14306 25454 14308 25506
rect 13356 24994 13412 25004
rect 13468 25004 13748 25060
rect 14028 25396 14084 25406
rect 12124 24882 12180 24892
rect 12460 24948 12516 24986
rect 12460 24882 12516 24892
rect 11788 24770 11844 24780
rect 12348 24834 12404 24846
rect 12348 24782 12350 24834
rect 12402 24782 12404 24834
rect 11676 24722 11732 24734
rect 11676 24670 11678 24722
rect 11730 24670 11732 24722
rect 11564 24164 11620 24174
rect 10892 22484 10948 22876
rect 10892 22418 10948 22428
rect 11228 23100 11396 23156
rect 11452 23268 11508 23278
rect 11452 23154 11508 23212
rect 11452 23102 11454 23154
rect 11506 23102 11508 23154
rect 11004 21812 11060 21822
rect 10668 21410 10724 21420
rect 10780 21698 10836 21710
rect 10780 21646 10782 21698
rect 10834 21646 10836 21698
rect 10556 20638 10558 20690
rect 10610 20638 10612 20690
rect 10556 20626 10612 20638
rect 10668 21252 10724 21262
rect 10668 20690 10724 21196
rect 10668 20638 10670 20690
rect 10722 20638 10724 20690
rect 10444 20580 10500 20590
rect 10444 20486 10500 20524
rect 10332 20300 10500 20356
rect 10220 20066 10276 20076
rect 10332 20130 10388 20142
rect 10332 20078 10334 20130
rect 10386 20078 10388 20130
rect 9660 19908 9716 19918
rect 9660 19814 9716 19852
rect 9772 19572 9828 19964
rect 9996 19954 10052 19964
rect 10332 19908 10388 20078
rect 10332 19842 10388 19852
rect 9772 19516 9940 19572
rect 9548 19404 9828 19460
rect 9436 19348 9492 19358
rect 9212 19346 9492 19348
rect 9212 19294 9438 19346
rect 9490 19294 9492 19346
rect 9212 19292 9492 19294
rect 9212 19234 9268 19292
rect 9436 19282 9492 19292
rect 9772 19346 9828 19404
rect 9772 19294 9774 19346
rect 9826 19294 9828 19346
rect 9212 19182 9214 19234
rect 9266 19182 9268 19234
rect 9212 19170 9268 19182
rect 9772 19236 9828 19294
rect 9772 19170 9828 19180
rect 8876 19068 9044 19124
rect 8988 18676 9044 19068
rect 9100 18788 9156 19068
rect 9528 18844 9792 18854
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9100 18732 9380 18788
rect 9528 18778 9792 18788
rect 8988 18620 9268 18676
rect 8764 18564 8820 18574
rect 8428 17778 8484 17836
rect 8428 17726 8430 17778
rect 8482 17726 8484 17778
rect 8428 17332 8484 17726
rect 8204 17276 8372 17332
rect 7588 16828 7924 16884
rect 7980 16996 8036 17006
rect 7532 16790 7588 16828
rect 6076 16770 6356 16772
rect 6076 16718 6078 16770
rect 6130 16718 6356 16770
rect 6076 16716 6356 16718
rect 6076 16706 6132 16716
rect 7644 16660 7700 16670
rect 7980 16660 8036 16940
rect 8092 16994 8148 17276
rect 8204 17108 8260 17118
rect 8204 17014 8260 17052
rect 8092 16942 8094 16994
rect 8146 16942 8148 16994
rect 8092 16930 8148 16942
rect 8316 16772 8372 17276
rect 8428 17266 8484 17276
rect 8540 18562 8820 18564
rect 8540 18510 8766 18562
rect 8818 18510 8820 18562
rect 8540 18508 8820 18510
rect 8540 17668 8596 18508
rect 8764 18498 8820 18508
rect 8876 18564 8932 18574
rect 8932 18508 9156 18564
rect 8876 18470 8932 18508
rect 8876 18228 8932 18238
rect 8876 18134 8932 18172
rect 9100 17668 9156 18508
rect 8428 17108 8484 17118
rect 8540 17108 8596 17612
rect 8428 17106 8596 17108
rect 8428 17054 8430 17106
rect 8482 17054 8596 17106
rect 8428 17052 8596 17054
rect 8652 17666 9156 17668
rect 8652 17614 9102 17666
rect 9154 17614 9156 17666
rect 8652 17612 9156 17614
rect 8652 17106 8708 17612
rect 9100 17556 9156 17612
rect 9100 17490 9156 17500
rect 9212 18340 9268 18620
rect 9324 18564 9380 18732
rect 9884 18676 9940 19516
rect 10332 19236 10388 19246
rect 9772 18620 9940 18676
rect 9996 19122 10052 19134
rect 9996 19070 9998 19122
rect 10050 19070 10052 19122
rect 9996 19012 10052 19070
rect 9548 18564 9604 18574
rect 9324 18562 9604 18564
rect 9324 18510 9550 18562
rect 9602 18510 9604 18562
rect 9324 18508 9604 18510
rect 9548 18498 9604 18508
rect 9660 18564 9716 18574
rect 9660 18470 9716 18508
rect 9772 18340 9828 18620
rect 9212 18284 9828 18340
rect 9884 18450 9940 18462
rect 9884 18398 9886 18450
rect 9938 18398 9940 18450
rect 9884 18340 9940 18398
rect 8876 17444 8932 17454
rect 8876 17442 9044 17444
rect 8876 17390 8878 17442
rect 8930 17390 9044 17442
rect 8876 17388 9044 17390
rect 8876 17378 8932 17388
rect 8988 17332 9044 17388
rect 9212 17332 9268 18284
rect 9884 18274 9940 18284
rect 9996 18116 10052 18956
rect 10332 18900 10388 19180
rect 10332 18834 10388 18844
rect 10332 18340 10388 18350
rect 10220 18338 10388 18340
rect 10220 18286 10334 18338
rect 10386 18286 10388 18338
rect 10220 18284 10388 18286
rect 10108 18228 10164 18238
rect 10108 18134 10164 18172
rect 9772 18060 10052 18116
rect 9548 17892 9604 17902
rect 9548 17798 9604 17836
rect 9772 17554 9828 18060
rect 10220 18004 10276 18284
rect 10332 18274 10388 18284
rect 9884 17948 10276 18004
rect 10444 18228 10500 20300
rect 10556 20018 10612 20030
rect 10556 19966 10558 20018
rect 10610 19966 10612 20018
rect 10556 19348 10612 19966
rect 10668 20020 10724 20638
rect 10780 20580 10836 21646
rect 10892 21588 10948 21598
rect 10892 21494 10948 21532
rect 11004 20914 11060 21756
rect 11228 21810 11284 23100
rect 11452 23090 11508 23102
rect 11564 23044 11620 24108
rect 11676 23938 11732 24670
rect 12236 24724 12292 24734
rect 12348 24724 12404 24782
rect 12684 24836 12740 24874
rect 12684 24770 12740 24780
rect 13132 24836 13188 24846
rect 12460 24724 12516 24734
rect 12348 24668 12460 24724
rect 12236 24630 12292 24668
rect 12460 24658 12516 24668
rect 12572 24722 12628 24734
rect 12572 24670 12574 24722
rect 12626 24670 12628 24722
rect 12124 24164 12180 24174
rect 11900 24162 12180 24164
rect 11900 24110 12126 24162
rect 12178 24110 12180 24162
rect 11900 24108 12180 24110
rect 11676 23886 11678 23938
rect 11730 23886 11732 23938
rect 11676 23604 11732 23886
rect 11676 23538 11732 23548
rect 11788 23940 11844 23950
rect 11788 23266 11844 23884
rect 11788 23214 11790 23266
rect 11842 23214 11844 23266
rect 11788 23202 11844 23214
rect 11676 23044 11732 23054
rect 11564 23042 11732 23044
rect 11564 22990 11678 23042
rect 11730 22990 11732 23042
rect 11564 22988 11732 22990
rect 11340 22930 11396 22942
rect 11340 22878 11342 22930
rect 11394 22878 11396 22930
rect 11340 22820 11396 22878
rect 11340 22754 11396 22764
rect 11228 21758 11230 21810
rect 11282 21758 11284 21810
rect 11228 21746 11284 21758
rect 11340 22484 11396 22494
rect 11340 21810 11396 22428
rect 11564 22036 11620 22988
rect 11676 22978 11732 22988
rect 11564 21970 11620 21980
rect 11340 21758 11342 21810
rect 11394 21758 11396 21810
rect 11340 21746 11396 21758
rect 11564 21588 11620 21598
rect 11452 21586 11620 21588
rect 11452 21534 11566 21586
rect 11618 21534 11620 21586
rect 11452 21532 11620 21534
rect 11452 21026 11508 21532
rect 11564 21522 11620 21532
rect 11900 21586 11956 24108
rect 12124 24098 12180 24108
rect 12012 23828 12068 23838
rect 12012 23734 12068 23772
rect 12236 23828 12292 23838
rect 12124 23714 12180 23726
rect 12124 23662 12126 23714
rect 12178 23662 12180 23714
rect 12124 23380 12180 23662
rect 12124 23314 12180 23324
rect 12124 23156 12180 23166
rect 12124 23062 12180 23100
rect 11900 21534 11902 21586
rect 11954 21534 11956 21586
rect 11900 21522 11956 21534
rect 11452 20974 11454 21026
rect 11506 20974 11508 21026
rect 11452 20962 11508 20974
rect 12012 21476 12068 21486
rect 11004 20862 11006 20914
rect 11058 20862 11060 20914
rect 11004 20850 11060 20862
rect 11340 20692 11396 20702
rect 10780 20514 10836 20524
rect 10892 20690 11396 20692
rect 10892 20638 11342 20690
rect 11394 20638 11396 20690
rect 10892 20636 11396 20638
rect 10780 20020 10836 20030
rect 10668 20018 10836 20020
rect 10668 19966 10782 20018
rect 10834 19966 10836 20018
rect 10668 19964 10836 19966
rect 10780 19954 10836 19964
rect 10892 19460 10948 20636
rect 11340 20626 11396 20636
rect 11452 20580 11508 20590
rect 11340 20244 11396 20254
rect 10556 19282 10612 19292
rect 10668 19404 10948 19460
rect 11004 19796 11060 19806
rect 10556 19124 10612 19134
rect 10556 19030 10612 19068
rect 9884 17890 9940 17948
rect 9884 17838 9886 17890
rect 9938 17838 9940 17890
rect 9884 17826 9940 17838
rect 10220 17668 10276 17678
rect 10220 17574 10276 17612
rect 9772 17502 9774 17554
rect 9826 17502 9828 17554
rect 9772 17444 9828 17502
rect 9772 17378 9828 17388
rect 10444 17442 10500 18172
rect 10444 17390 10446 17442
rect 10498 17390 10500 17442
rect 8988 17276 9268 17332
rect 9528 17276 9792 17286
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9528 17210 9792 17220
rect 8652 17054 8654 17106
rect 8706 17054 8708 17106
rect 8428 17042 8484 17052
rect 8652 17042 8708 17054
rect 9884 17108 9940 17118
rect 9884 17014 9940 17052
rect 10444 16996 10500 17390
rect 10556 18452 10612 18462
rect 10556 17108 10612 18396
rect 10668 18450 10724 19404
rect 10780 19236 10836 19246
rect 11004 19236 11060 19740
rect 11340 19346 11396 20188
rect 11452 20018 11508 20524
rect 12012 20130 12068 21420
rect 12124 20244 12180 20254
rect 12236 20244 12292 23772
rect 12572 23828 12628 24670
rect 13132 24722 13188 24780
rect 13468 24834 13524 25004
rect 13468 24782 13470 24834
rect 13522 24782 13524 24834
rect 13468 24770 13524 24782
rect 14028 24948 14084 25340
rect 14252 25284 14308 25454
rect 14252 25218 14308 25228
rect 14700 25508 14756 25518
rect 13132 24670 13134 24722
rect 13186 24670 13188 24722
rect 13132 24658 13188 24670
rect 13244 24724 13300 24734
rect 13020 23940 13076 23950
rect 13020 23846 13076 23884
rect 12572 23762 12628 23772
rect 12348 23604 12404 23614
rect 12572 23604 12628 23614
rect 12348 21924 12404 23548
rect 12460 23548 12572 23604
rect 12460 23380 12516 23548
rect 12572 23538 12628 23548
rect 12460 23314 12516 23324
rect 12908 23380 12964 23390
rect 12908 23286 12964 23324
rect 12684 23268 12740 23278
rect 12684 23174 12740 23212
rect 12460 23154 12516 23166
rect 12460 23102 12462 23154
rect 12514 23102 12516 23154
rect 12460 22596 12516 23102
rect 13020 23156 13076 23166
rect 13076 23100 13188 23156
rect 13020 23090 13076 23100
rect 12572 23044 12628 23054
rect 12572 22950 12628 22988
rect 12460 22540 13076 22596
rect 12908 22372 12964 22382
rect 12348 21858 12404 21868
rect 12460 22316 12908 22372
rect 12348 21700 12404 21710
rect 12348 21252 12404 21644
rect 12348 21186 12404 21196
rect 12348 20916 12404 20926
rect 12460 20916 12516 22316
rect 12908 22278 12964 22316
rect 12684 21812 12740 21822
rect 12684 21718 12740 21756
rect 13020 21476 13076 22540
rect 13020 21410 13076 21420
rect 13132 21586 13188 23100
rect 13244 21700 13300 24668
rect 13356 24610 13412 24622
rect 13356 24558 13358 24610
rect 13410 24558 13412 24610
rect 13356 23940 13412 24558
rect 13686 24332 13950 24342
rect 13742 24276 13790 24332
rect 13846 24276 13894 24332
rect 13686 24266 13950 24276
rect 13580 24164 13636 24174
rect 13580 24162 13860 24164
rect 13580 24110 13582 24162
rect 13634 24110 13860 24162
rect 13580 24108 13860 24110
rect 13580 24098 13636 24108
rect 13468 23940 13524 23950
rect 13692 23940 13748 23950
rect 13356 23938 13524 23940
rect 13356 23886 13470 23938
rect 13522 23886 13524 23938
rect 13356 23884 13524 23886
rect 13468 23874 13524 23884
rect 13580 23884 13692 23940
rect 13580 23380 13636 23884
rect 13692 23874 13748 23884
rect 13692 23716 13748 23726
rect 13692 23622 13748 23660
rect 13692 23380 13748 23390
rect 13580 23378 13748 23380
rect 13580 23326 13694 23378
rect 13746 23326 13748 23378
rect 13580 23324 13748 23326
rect 13692 23314 13748 23324
rect 13804 23266 13860 24108
rect 14028 23940 14084 24892
rect 14364 25060 14420 25070
rect 14252 24834 14308 24846
rect 14252 24782 14254 24834
rect 14306 24782 14308 24834
rect 14140 24722 14196 24734
rect 14140 24670 14142 24722
rect 14194 24670 14196 24722
rect 14140 24164 14196 24670
rect 14140 24098 14196 24108
rect 14140 23940 14196 23950
rect 14028 23938 14196 23940
rect 14028 23886 14142 23938
rect 14194 23886 14196 23938
rect 14028 23884 14196 23886
rect 14140 23874 14196 23884
rect 13916 23828 13972 23838
rect 13916 23734 13972 23772
rect 14140 23716 14196 23726
rect 13916 23380 13972 23390
rect 13972 23324 14084 23380
rect 13916 23314 13972 23324
rect 13804 23214 13806 23266
rect 13858 23214 13860 23266
rect 13804 23202 13860 23214
rect 13468 23154 13524 23166
rect 13468 23102 13470 23154
rect 13522 23102 13524 23154
rect 13468 21924 13524 23102
rect 13686 22764 13950 22774
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13686 22698 13950 22708
rect 14028 22596 14084 23324
rect 14140 23378 14196 23660
rect 14140 23326 14142 23378
rect 14194 23326 14196 23378
rect 14140 23314 14196 23326
rect 14252 23156 14308 24782
rect 14364 23380 14420 25004
rect 14476 24722 14532 24734
rect 14476 24670 14478 24722
rect 14530 24670 14532 24722
rect 14476 24388 14532 24670
rect 14588 24724 14644 24734
rect 14588 24630 14644 24668
rect 14476 24322 14532 24332
rect 14700 24164 14756 25452
rect 15148 25506 15204 25518
rect 15148 25454 15150 25506
rect 15202 25454 15204 25506
rect 14924 25396 14980 25406
rect 14924 25302 14980 25340
rect 15148 24946 15204 25454
rect 15484 25508 15540 25518
rect 15484 25414 15540 25452
rect 15596 25172 15652 26460
rect 15484 25116 15652 25172
rect 15708 26292 15764 26302
rect 15148 24894 15150 24946
rect 15202 24894 15204 24946
rect 15148 24882 15204 24894
rect 15260 24948 15316 24958
rect 15260 24854 15316 24892
rect 15036 24722 15092 24734
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 15036 24388 15092 24670
rect 14476 24108 14756 24164
rect 14924 24332 15092 24388
rect 14476 23716 14532 24108
rect 14924 24052 14980 24332
rect 14700 24050 14980 24052
rect 14700 23998 14926 24050
rect 14978 23998 14980 24050
rect 14700 23996 14980 23998
rect 14476 23650 14532 23660
rect 14588 23940 14644 23950
rect 14364 23314 14420 23324
rect 14364 23156 14420 23166
rect 14252 23100 14364 23156
rect 14364 23090 14420 23100
rect 14476 23154 14532 23166
rect 14476 23102 14478 23154
rect 14530 23102 14532 23154
rect 13804 22540 14084 22596
rect 13580 22260 13636 22270
rect 13636 22204 13748 22260
rect 13580 22194 13636 22204
rect 13244 21634 13300 21644
rect 13356 21868 13524 21924
rect 13580 22036 13636 22046
rect 13356 21812 13412 21868
rect 13132 21534 13134 21586
rect 13186 21534 13188 21586
rect 12796 21028 12852 21038
rect 12796 20934 12852 20972
rect 12348 20914 12516 20916
rect 12348 20862 12350 20914
rect 12402 20862 12516 20914
rect 12348 20860 12516 20862
rect 12348 20850 12404 20860
rect 12180 20188 12292 20244
rect 12684 20690 12740 20702
rect 12684 20638 12686 20690
rect 12738 20638 12740 20690
rect 12684 20244 12740 20638
rect 12796 20580 12852 20590
rect 12796 20486 12852 20524
rect 12796 20244 12852 20254
rect 12684 20242 12852 20244
rect 12684 20190 12798 20242
rect 12850 20190 12852 20242
rect 12684 20188 12852 20190
rect 12124 20178 12180 20188
rect 12796 20178 12852 20188
rect 12012 20078 12014 20130
rect 12066 20078 12068 20130
rect 12012 20066 12068 20078
rect 12460 20132 12516 20142
rect 12460 20038 12516 20076
rect 12572 20130 12628 20142
rect 12572 20078 12574 20130
rect 12626 20078 12628 20130
rect 11900 20020 11956 20030
rect 11452 19966 11454 20018
rect 11506 19966 11508 20018
rect 11452 19954 11508 19966
rect 11564 20018 11956 20020
rect 11564 19966 11902 20018
rect 11954 19966 11956 20018
rect 11564 19964 11956 19966
rect 11340 19294 11342 19346
rect 11394 19294 11396 19346
rect 11340 19282 11396 19294
rect 10780 19234 11172 19236
rect 10780 19182 10782 19234
rect 10834 19182 11172 19234
rect 10780 19180 11172 19182
rect 10780 19170 10836 19180
rect 10892 19012 10948 19022
rect 10780 18900 10836 18910
rect 10780 18674 10836 18844
rect 10780 18622 10782 18674
rect 10834 18622 10836 18674
rect 10780 18610 10836 18622
rect 10668 18398 10670 18450
rect 10722 18398 10724 18450
rect 10668 18386 10724 18398
rect 10780 17892 10836 17902
rect 10892 17892 10948 18956
rect 11004 19010 11060 19022
rect 11004 18958 11006 19010
rect 11058 18958 11060 19010
rect 11004 18228 11060 18958
rect 11116 18788 11172 19180
rect 11116 18722 11172 18732
rect 11228 19122 11284 19134
rect 11228 19070 11230 19122
rect 11282 19070 11284 19122
rect 11228 18676 11284 19070
rect 11452 18676 11508 18686
rect 11564 18676 11620 19964
rect 11900 19954 11956 19964
rect 12124 20018 12180 20030
rect 12124 19966 12126 20018
rect 12178 19966 12180 20018
rect 12124 19572 12180 19966
rect 12572 19796 12628 20078
rect 13132 20132 13188 21534
rect 13356 21028 13412 21756
rect 13580 21810 13636 21980
rect 13580 21758 13582 21810
rect 13634 21758 13636 21810
rect 13580 21746 13636 21758
rect 13692 21810 13748 22204
rect 13692 21758 13694 21810
rect 13746 21758 13748 21810
rect 13692 21746 13748 21758
rect 13804 21810 13860 22540
rect 13804 21758 13806 21810
rect 13858 21758 13860 21810
rect 13804 21746 13860 21758
rect 14476 21812 14532 23102
rect 13468 21700 13524 21738
rect 13468 21634 13524 21644
rect 14140 21588 14196 21598
rect 14028 21586 14196 21588
rect 14028 21534 14142 21586
rect 14194 21534 14196 21586
rect 14028 21532 14196 21534
rect 13686 21196 13950 21206
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13686 21130 13950 21140
rect 13356 20972 13636 21028
rect 13580 20804 13636 20972
rect 14028 20916 14084 21532
rect 14140 21522 14196 21532
rect 14476 21586 14532 21756
rect 14476 21534 14478 21586
rect 14530 21534 14532 21586
rect 14476 21522 14532 21534
rect 13468 20692 13524 20702
rect 13132 20066 13188 20076
rect 13356 20690 13524 20692
rect 13356 20638 13470 20690
rect 13522 20638 13524 20690
rect 13356 20636 13524 20638
rect 12572 19730 12628 19740
rect 12124 19516 12740 19572
rect 12684 19458 12740 19516
rect 12684 19406 12686 19458
rect 12738 19406 12740 19458
rect 12684 19394 12740 19406
rect 12348 19348 12404 19358
rect 12236 19292 12348 19348
rect 12236 19234 12292 19292
rect 12348 19282 12404 19292
rect 13356 19348 13412 20636
rect 13468 20626 13524 20636
rect 13580 20690 13636 20748
rect 13804 20860 14084 20916
rect 13804 20802 13860 20860
rect 13804 20750 13806 20802
rect 13858 20750 13860 20802
rect 13804 20738 13860 20750
rect 14140 20804 14196 20814
rect 14140 20710 14196 20748
rect 14364 20804 14420 20814
rect 13580 20638 13582 20690
rect 13634 20638 13636 20690
rect 13580 20626 13636 20638
rect 14364 20690 14420 20748
rect 14364 20638 14366 20690
rect 14418 20638 14420 20690
rect 14364 20580 14420 20638
rect 14364 20514 14420 20524
rect 13580 20132 13636 20142
rect 13356 19282 13412 19292
rect 13468 20076 13580 20132
rect 12236 19182 12238 19234
rect 12290 19182 12292 19234
rect 12236 19170 12292 19182
rect 12796 19122 12852 19134
rect 12796 19070 12798 19122
rect 12850 19070 12852 19122
rect 11900 19012 11956 19022
rect 12124 19012 12180 19022
rect 11900 18918 11956 18956
rect 12012 19010 12180 19012
rect 12012 18958 12126 19010
rect 12178 18958 12180 19010
rect 12012 18956 12180 18958
rect 11284 18620 11396 18676
rect 11228 18610 11284 18620
rect 11228 18450 11284 18462
rect 11228 18398 11230 18450
rect 11282 18398 11284 18450
rect 11116 18228 11172 18238
rect 11228 18228 11284 18398
rect 11340 18452 11396 18620
rect 11452 18674 11620 18676
rect 11452 18622 11454 18674
rect 11506 18622 11620 18674
rect 11452 18620 11620 18622
rect 11452 18610 11508 18620
rect 11452 18452 11508 18462
rect 11788 18452 11844 18462
rect 12012 18452 12068 18956
rect 12124 18946 12180 18956
rect 12348 19012 12404 19022
rect 12348 19010 12628 19012
rect 12348 18958 12350 19010
rect 12402 18958 12628 19010
rect 12348 18956 12628 18958
rect 12348 18946 12404 18956
rect 12572 18676 12628 18956
rect 12684 18676 12740 18686
rect 12572 18674 12740 18676
rect 12572 18622 12686 18674
rect 12738 18622 12740 18674
rect 12572 18620 12740 18622
rect 12684 18610 12740 18620
rect 11340 18450 11732 18452
rect 11340 18398 11454 18450
rect 11506 18398 11732 18450
rect 11340 18396 11732 18398
rect 11452 18386 11508 18396
rect 11004 18172 11116 18228
rect 11172 18172 11284 18228
rect 11676 18228 11732 18396
rect 11844 18396 12068 18452
rect 11788 18358 11844 18396
rect 12124 18338 12180 18350
rect 12124 18286 12126 18338
rect 12178 18286 12180 18338
rect 12124 18228 12180 18286
rect 12348 18340 12404 18350
rect 12348 18246 12404 18284
rect 11676 18172 12180 18228
rect 11116 18162 11172 18172
rect 12796 18116 12852 19070
rect 12796 18050 12852 18060
rect 10780 17890 10948 17892
rect 10780 17838 10782 17890
rect 10834 17838 10948 17890
rect 10780 17836 10948 17838
rect 10780 17826 10836 17836
rect 11004 17780 11060 17790
rect 10892 17668 10948 17678
rect 11004 17668 11060 17724
rect 10892 17666 11060 17668
rect 10892 17614 10894 17666
rect 10946 17614 11060 17666
rect 10892 17612 11060 17614
rect 10892 17602 10948 17612
rect 10668 17556 10724 17566
rect 10668 17462 10724 17500
rect 11228 17554 11284 17566
rect 11228 17502 11230 17554
rect 11282 17502 11284 17554
rect 11116 17444 11172 17454
rect 11116 17350 11172 17388
rect 10556 17042 10612 17052
rect 11228 17108 11284 17502
rect 11228 17042 11284 17052
rect 10444 16930 10500 16940
rect 8316 16706 8372 16716
rect 8876 16884 8932 16894
rect 9548 16884 9604 16894
rect 8876 16882 9604 16884
rect 8876 16830 8878 16882
rect 8930 16830 9550 16882
rect 9602 16830 9604 16882
rect 8876 16828 9604 16830
rect 7644 16658 8036 16660
rect 7644 16606 7646 16658
rect 7698 16606 8036 16658
rect 7644 16604 8036 16606
rect 7644 16594 7700 16604
rect 6300 15874 6356 15886
rect 6300 15822 6302 15874
rect 6354 15822 6356 15874
rect 5852 15092 6132 15148
rect 4620 14642 4676 14654
rect 4620 14590 4622 14642
rect 4674 14590 4676 14642
rect 2940 14242 2996 14252
rect 3724 14308 3780 14318
rect 3724 13074 3780 14252
rect 4620 14308 4676 14590
rect 4620 14242 4676 14252
rect 5068 14306 5124 15036
rect 5740 15026 5796 15036
rect 5370 14924 5634 14934
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5370 14858 5634 14868
rect 5068 14254 5070 14306
rect 5122 14254 5124 14306
rect 5068 13524 5124 14254
rect 5628 14308 5684 14318
rect 5516 13748 5572 13758
rect 5516 13654 5572 13692
rect 5628 13634 5684 14252
rect 5964 14306 6020 14318
rect 5964 14254 5966 14306
rect 6018 14254 6020 14306
rect 5964 14084 6020 14254
rect 5964 14018 6020 14028
rect 5964 13860 6020 13870
rect 5628 13582 5630 13634
rect 5682 13582 5684 13634
rect 5628 13570 5684 13582
rect 5740 13804 5964 13860
rect 5068 13458 5124 13468
rect 5370 13356 5634 13366
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5370 13290 5634 13300
rect 3724 13022 3726 13074
rect 3778 13022 3780 13074
rect 3724 13010 3780 13022
rect 4620 13074 4676 13086
rect 4620 13022 4622 13074
rect 4674 13022 4676 13074
rect 4284 12962 4340 12974
rect 4284 12910 4286 12962
rect 4338 12910 4340 12962
rect 3388 12738 3444 12750
rect 3388 12686 3390 12738
rect 3442 12686 3444 12738
rect 2492 11554 2548 11564
rect 2828 12628 2884 12638
rect 2828 12178 2884 12572
rect 2828 12126 2830 12178
rect 2882 12126 2884 12178
rect 2380 11454 2382 11506
rect 2434 11454 2436 11506
rect 2380 11442 2436 11454
rect 2156 11396 2212 11406
rect 2156 11302 2212 11340
rect 2268 11172 2324 11182
rect 2156 11170 2324 11172
rect 2156 11118 2270 11170
rect 2322 11118 2324 11170
rect 2156 11116 2324 11118
rect 2156 8372 2212 11116
rect 2268 11106 2324 11116
rect 2492 11170 2548 11182
rect 2492 11118 2494 11170
rect 2546 11118 2548 11170
rect 2492 10948 2548 11118
rect 2604 11172 2660 11182
rect 2604 11078 2660 11116
rect 2492 10892 2772 10948
rect 2716 10836 2772 10892
rect 2716 10770 2772 10780
rect 2716 10612 2772 10622
rect 2268 10610 2772 10612
rect 2268 10558 2718 10610
rect 2770 10558 2772 10610
rect 2268 10556 2772 10558
rect 2268 10050 2324 10556
rect 2716 10546 2772 10556
rect 2268 9998 2270 10050
rect 2322 9998 2324 10050
rect 2268 9986 2324 9998
rect 2604 9940 2660 9950
rect 2380 8930 2436 8942
rect 2380 8878 2382 8930
rect 2434 8878 2436 8930
rect 2380 8596 2436 8878
rect 2492 8596 2548 8606
rect 2380 8540 2492 8596
rect 2492 8530 2548 8540
rect 2156 8306 2212 8316
rect 2604 8146 2660 9884
rect 2716 9828 2772 9838
rect 2716 9734 2772 9772
rect 2828 9266 2884 12126
rect 3164 12290 3220 12302
rect 3164 12238 3166 12290
rect 3218 12238 3220 12290
rect 3164 11732 3220 12238
rect 3388 12292 3444 12686
rect 3612 12740 3668 12750
rect 3612 12646 3668 12684
rect 3836 12738 3892 12750
rect 3836 12686 3838 12738
rect 3890 12686 3892 12738
rect 3836 12404 3892 12686
rect 4172 12404 4228 12414
rect 3836 12402 4228 12404
rect 3836 12350 4174 12402
rect 4226 12350 4228 12402
rect 3836 12348 4228 12350
rect 4172 12338 4228 12348
rect 3724 12292 3780 12302
rect 3388 12290 3780 12292
rect 3388 12238 3726 12290
rect 3778 12238 3780 12290
rect 3388 12236 3780 12238
rect 3500 11956 3556 11966
rect 2940 11676 3220 11732
rect 3388 11900 3500 11956
rect 2940 10724 2996 11676
rect 3052 11508 3108 11518
rect 3052 11414 3108 11452
rect 3276 11394 3332 11406
rect 3276 11342 3278 11394
rect 3330 11342 3332 11394
rect 3276 10948 3332 11342
rect 3276 10882 3332 10892
rect 2940 10658 2996 10668
rect 3276 10724 3332 10734
rect 3276 10630 3332 10668
rect 3052 10610 3108 10622
rect 3052 10558 3054 10610
rect 3106 10558 3108 10610
rect 2940 10500 2996 10510
rect 2940 10406 2996 10444
rect 3052 10052 3108 10558
rect 3052 9986 3108 9996
rect 3164 9940 3220 9950
rect 3164 9846 3220 9884
rect 2940 9826 2996 9838
rect 3388 9828 3444 11900
rect 3500 11862 3556 11900
rect 3724 11732 3780 12236
rect 3836 12180 3892 12190
rect 3836 12066 3892 12124
rect 3836 12014 3838 12066
rect 3890 12014 3892 12066
rect 3836 12002 3892 12014
rect 4172 12178 4228 12190
rect 4172 12126 4174 12178
rect 4226 12126 4228 12178
rect 4172 11844 4228 12126
rect 4172 11778 4228 11788
rect 3724 11666 3780 11676
rect 4284 11506 4340 12910
rect 4620 12516 4676 13022
rect 5628 13076 5684 13086
rect 5740 13076 5796 13804
rect 5964 13766 6020 13804
rect 6076 13188 6132 15092
rect 6300 15092 6356 15822
rect 6412 15202 6468 15214
rect 6412 15150 6414 15202
rect 6466 15150 6468 15202
rect 6412 15148 6468 15150
rect 8540 15204 8596 15214
rect 8876 15204 8932 16828
rect 9548 16818 9604 16828
rect 10780 16884 10836 16894
rect 10780 16210 10836 16828
rect 12236 16884 12292 16894
rect 12236 16790 12292 16828
rect 12348 16882 12404 16894
rect 12348 16830 12350 16882
rect 12402 16830 12404 16882
rect 10780 16158 10782 16210
rect 10834 16158 10836 16210
rect 10780 16146 10836 16158
rect 11676 16772 11732 16782
rect 9996 16098 10052 16110
rect 9996 16046 9998 16098
rect 10050 16046 10052 16098
rect 9660 15876 9716 15886
rect 9996 15876 10052 16046
rect 9660 15874 10052 15876
rect 9660 15822 9662 15874
rect 9714 15822 10052 15874
rect 9660 15820 10052 15822
rect 9660 15810 9716 15820
rect 9528 15708 9792 15718
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9528 15642 9792 15652
rect 8540 15202 8932 15204
rect 8540 15150 8542 15202
rect 8594 15150 8932 15202
rect 8540 15148 8932 15150
rect 8988 15314 9044 15326
rect 8988 15262 8990 15314
rect 9042 15262 9044 15314
rect 6412 15092 6804 15148
rect 8540 15138 8596 15148
rect 6300 15026 6356 15036
rect 6748 13970 6804 15092
rect 8988 15092 9044 15262
rect 6748 13918 6750 13970
rect 6802 13918 6804 13970
rect 6748 13906 6804 13918
rect 8428 14420 8484 14430
rect 8988 14420 9044 15036
rect 9996 15092 10052 15820
rect 11228 15316 11284 15326
rect 11228 15222 11284 15260
rect 9996 15026 10052 15036
rect 8428 14418 9044 14420
rect 8428 14366 8430 14418
rect 8482 14366 9044 14418
rect 8428 14364 9044 14366
rect 7308 13860 7364 13870
rect 7308 13766 7364 13804
rect 7420 13860 7476 13870
rect 7644 13860 7700 13870
rect 7420 13858 7644 13860
rect 7420 13806 7422 13858
rect 7474 13806 7644 13858
rect 7420 13804 7644 13806
rect 7420 13794 7476 13804
rect 7644 13794 7700 13804
rect 5628 13074 5796 13076
rect 5628 13022 5630 13074
rect 5682 13022 5796 13074
rect 5628 13020 5796 13022
rect 5964 13132 6132 13188
rect 6300 13746 6356 13758
rect 6524 13748 6580 13758
rect 6860 13748 6916 13758
rect 6300 13694 6302 13746
rect 6354 13694 6356 13746
rect 5628 13010 5684 13020
rect 4956 12964 5012 12974
rect 4676 12460 4788 12516
rect 4620 12450 4676 12460
rect 4508 12180 4564 12190
rect 4508 12086 4564 12124
rect 4620 12178 4676 12190
rect 4620 12126 4622 12178
rect 4674 12126 4676 12178
rect 4396 11956 4452 11966
rect 4620 11956 4676 12126
rect 4452 11900 4676 11956
rect 4396 11890 4452 11900
rect 4284 11454 4286 11506
rect 4338 11454 4340 11506
rect 4284 11442 4340 11454
rect 3500 11396 3556 11406
rect 3500 10724 3556 11340
rect 3612 11396 3668 11406
rect 4172 11396 4228 11406
rect 3612 11394 4228 11396
rect 3612 11342 3614 11394
rect 3666 11342 4174 11394
rect 4226 11342 4228 11394
rect 3612 11340 4228 11342
rect 3612 11330 3668 11340
rect 4172 11330 4228 11340
rect 4620 11394 4676 11406
rect 4620 11342 4622 11394
rect 4674 11342 4676 11394
rect 3612 11172 3668 11182
rect 3612 10836 3668 11116
rect 3724 11172 3780 11182
rect 3724 11170 4228 11172
rect 3724 11118 3726 11170
rect 3778 11118 4228 11170
rect 3724 11116 4228 11118
rect 3724 11106 3780 11116
rect 3724 10836 3780 10846
rect 3612 10834 3780 10836
rect 3612 10782 3726 10834
rect 3778 10782 3780 10834
rect 3612 10780 3780 10782
rect 3724 10770 3780 10780
rect 3500 10668 3668 10724
rect 3612 10612 3668 10668
rect 3836 10722 3892 10734
rect 3836 10670 3838 10722
rect 3890 10670 3892 10722
rect 3836 10612 3892 10670
rect 3612 10556 3892 10612
rect 3612 10388 3668 10398
rect 3612 10386 3892 10388
rect 3612 10334 3614 10386
rect 3666 10334 3892 10386
rect 3612 10332 3892 10334
rect 3612 10322 3668 10332
rect 3612 10052 3668 10062
rect 3612 9938 3668 9996
rect 3612 9886 3614 9938
rect 3666 9886 3668 9938
rect 3612 9874 3668 9886
rect 2940 9774 2942 9826
rect 2994 9774 2996 9826
rect 2940 9492 2996 9774
rect 2940 9426 2996 9436
rect 3276 9772 3444 9828
rect 2828 9214 2830 9266
rect 2882 9214 2884 9266
rect 2828 9202 2884 9214
rect 3276 9268 3332 9772
rect 3500 9602 3556 9614
rect 3500 9550 3502 9602
rect 3554 9550 3556 9602
rect 3500 9492 3556 9550
rect 3724 9604 3780 9614
rect 3724 9510 3780 9548
rect 3500 9426 3556 9436
rect 3836 9268 3892 10332
rect 4060 9828 4116 9838
rect 3948 9268 4004 9278
rect 3276 9212 3556 9268
rect 3836 9266 4004 9268
rect 3836 9214 3950 9266
rect 4002 9214 4004 9266
rect 3836 9212 4004 9214
rect 3164 9042 3220 9054
rect 3164 8990 3166 9042
rect 3218 8990 3220 9042
rect 3164 8428 3220 8990
rect 2716 8372 3220 8428
rect 3500 9042 3556 9212
rect 3948 9202 4004 9212
rect 3724 9044 3780 9054
rect 3500 8990 3502 9042
rect 3554 8990 3556 9042
rect 2716 8370 2772 8372
rect 2716 8318 2718 8370
rect 2770 8318 2772 8370
rect 2716 8306 2772 8318
rect 3164 8260 3220 8270
rect 2940 8258 3220 8260
rect 2940 8206 3166 8258
rect 3218 8206 3220 8258
rect 2940 8204 3220 8206
rect 2604 8094 2606 8146
rect 2658 8094 2660 8146
rect 2268 8036 2324 8046
rect 2268 7474 2324 7980
rect 2492 7700 2548 7710
rect 2604 7700 2660 8094
rect 2828 8148 2884 8158
rect 2828 8054 2884 8092
rect 2492 7698 2660 7700
rect 2492 7646 2494 7698
rect 2546 7646 2660 7698
rect 2492 7644 2660 7646
rect 2492 7634 2548 7644
rect 2268 7422 2270 7474
rect 2322 7422 2324 7474
rect 2268 7410 2324 7422
rect 2604 7140 2660 7644
rect 2940 7698 2996 8204
rect 3164 8194 3220 8204
rect 3388 8258 3444 8270
rect 3388 8206 3390 8258
rect 3442 8206 3444 8258
rect 3388 8148 3444 8206
rect 3388 8082 3444 8092
rect 3500 7812 3556 8990
rect 2940 7646 2942 7698
rect 2994 7646 2996 7698
rect 2940 7634 2996 7646
rect 3388 7756 3556 7812
rect 3612 9042 3780 9044
rect 3612 8990 3726 9042
rect 3778 8990 3780 9042
rect 3612 8988 3780 8990
rect 3612 8596 3668 8988
rect 3724 8978 3780 8988
rect 3948 9044 4004 9054
rect 3612 8258 3668 8540
rect 3612 8206 3614 8258
rect 3666 8206 3668 8258
rect 2828 7474 2884 7486
rect 3052 7476 3108 7486
rect 2828 7422 2830 7474
rect 2882 7422 2884 7474
rect 2828 7252 2884 7422
rect 2828 7186 2884 7196
rect 2940 7474 3108 7476
rect 2940 7422 3054 7474
rect 3106 7422 3108 7474
rect 2940 7420 3108 7422
rect 2604 7074 2660 7084
rect 2828 7028 2884 7038
rect 2604 5908 2660 5918
rect 2604 5814 2660 5852
rect 2156 5796 2212 5806
rect 2156 5794 2548 5796
rect 2156 5742 2158 5794
rect 2210 5742 2548 5794
rect 2156 5740 2548 5742
rect 2156 5730 2212 5740
rect 2492 5124 2548 5740
rect 2828 5236 2884 6972
rect 2940 6132 2996 7420
rect 3052 7410 3108 7420
rect 3388 7252 3444 7756
rect 3500 7588 3556 7598
rect 3500 7474 3556 7532
rect 3500 7422 3502 7474
rect 3554 7422 3556 7474
rect 3500 7410 3556 7422
rect 3612 7476 3668 8206
rect 3612 7410 3668 7420
rect 3724 8818 3780 8830
rect 3724 8766 3726 8818
rect 3778 8766 3780 8818
rect 3388 7196 3668 7252
rect 3500 6916 3556 6926
rect 3500 6802 3556 6860
rect 3500 6750 3502 6802
rect 3554 6750 3556 6802
rect 3500 6738 3556 6750
rect 3388 6468 3444 6478
rect 2940 6066 2996 6076
rect 3052 6466 3444 6468
rect 3052 6414 3390 6466
rect 3442 6414 3444 6466
rect 3052 6412 3444 6414
rect 3052 5908 3108 6412
rect 3276 6132 3332 6142
rect 3276 6038 3332 6076
rect 3052 5814 3108 5852
rect 2940 5236 2996 5246
rect 2492 5030 2548 5068
rect 2604 5234 2996 5236
rect 2604 5182 2942 5234
rect 2994 5182 2996 5234
rect 2604 5180 2996 5182
rect 2492 4452 2548 4462
rect 2604 4452 2660 5180
rect 2940 5170 2996 5180
rect 3388 5234 3444 6412
rect 3612 6468 3668 7196
rect 3724 6580 3780 8766
rect 3836 8372 3892 8410
rect 3836 8306 3892 8316
rect 3836 8148 3892 8158
rect 3948 8148 4004 8988
rect 4060 8820 4116 9772
rect 4060 8754 4116 8764
rect 3836 8146 4004 8148
rect 3836 8094 3838 8146
rect 3890 8094 4004 8146
rect 3836 8092 4004 8094
rect 4172 8372 4228 11116
rect 4396 11170 4452 11182
rect 4396 11118 4398 11170
rect 4450 11118 4452 11170
rect 4396 10612 4452 11118
rect 4620 11060 4676 11342
rect 4732 11396 4788 12460
rect 4956 12290 5012 12908
rect 5852 12964 5908 12974
rect 5852 12870 5908 12908
rect 5068 12738 5124 12750
rect 5068 12686 5070 12738
rect 5122 12686 5124 12738
rect 5068 12404 5124 12686
rect 5068 12338 5124 12348
rect 5404 12740 5460 12750
rect 5404 12402 5460 12684
rect 5404 12350 5406 12402
rect 5458 12350 5460 12402
rect 5404 12338 5460 12350
rect 5516 12516 5572 12526
rect 5516 12402 5572 12460
rect 5516 12350 5518 12402
rect 5570 12350 5572 12402
rect 5516 12338 5572 12350
rect 4956 12238 4958 12290
rect 5010 12238 5012 12290
rect 4956 12226 5012 12238
rect 5852 12292 5908 12302
rect 5292 12178 5348 12190
rect 5292 12126 5294 12178
rect 5346 12126 5348 12178
rect 5292 11956 5348 12126
rect 5852 12178 5908 12236
rect 5852 12126 5854 12178
rect 5906 12126 5908 12178
rect 5852 12114 5908 12126
rect 5292 11890 5348 11900
rect 4956 11844 5012 11854
rect 4732 11330 4788 11340
rect 4844 11394 4900 11406
rect 4844 11342 4846 11394
rect 4898 11342 4900 11394
rect 4844 11172 4900 11342
rect 4620 11004 4788 11060
rect 4732 10834 4788 11004
rect 4732 10782 4734 10834
rect 4786 10782 4788 10834
rect 4732 10770 4788 10782
rect 4396 10546 4452 10556
rect 4732 10388 4788 10398
rect 4284 9492 4340 9502
rect 4284 9042 4340 9436
rect 4620 9268 4676 9278
rect 4620 9174 4676 9212
rect 4284 8990 4286 9042
rect 4338 8990 4340 9042
rect 4284 8932 4340 8990
rect 4284 8866 4340 8876
rect 4396 9154 4452 9166
rect 4396 9102 4398 9154
rect 4450 9102 4452 9154
rect 4396 8596 4452 9102
rect 4396 8530 4452 8540
rect 3836 8082 3892 8092
rect 4060 8034 4116 8046
rect 4060 7982 4062 8034
rect 4114 7982 4116 8034
rect 4060 7924 4116 7982
rect 4060 7858 4116 7868
rect 3836 7812 3892 7822
rect 3836 7474 3892 7756
rect 4172 7700 4228 8316
rect 4396 8260 4452 8270
rect 4172 7634 4228 7644
rect 4284 8148 4340 8158
rect 3836 7422 3838 7474
rect 3890 7422 3892 7474
rect 3836 7410 3892 7422
rect 3948 7476 4004 7486
rect 4284 7476 4340 8092
rect 3948 7474 4340 7476
rect 3948 7422 3950 7474
rect 4002 7422 4340 7474
rect 3948 7420 4340 7422
rect 4396 7474 4452 8204
rect 4508 8036 4564 8046
rect 4508 7942 4564 7980
rect 4508 7700 4564 7710
rect 4508 7586 4564 7644
rect 4508 7534 4510 7586
rect 4562 7534 4564 7586
rect 4508 7522 4564 7534
rect 4396 7422 4398 7474
rect 4450 7422 4452 7474
rect 3948 7410 4004 7420
rect 4396 7410 4452 7422
rect 4732 7474 4788 10332
rect 4844 10052 4900 11116
rect 4956 10834 5012 11788
rect 5370 11788 5634 11798
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5370 11722 5634 11732
rect 5964 11620 6020 13132
rect 6076 12962 6132 12974
rect 6076 12910 6078 12962
rect 6130 12910 6132 12962
rect 6076 12180 6132 12910
rect 6076 12114 6132 12124
rect 6188 12964 6244 12974
rect 5740 11564 6020 11620
rect 4956 10782 4958 10834
rect 5010 10782 5012 10834
rect 4956 10770 5012 10782
rect 5516 11396 5572 11406
rect 5068 10612 5124 10622
rect 5068 10518 5124 10556
rect 5516 10388 5572 11340
rect 5516 10322 5572 10332
rect 5370 10220 5634 10230
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5370 10154 5634 10164
rect 4956 10052 5012 10062
rect 4844 9996 4956 10052
rect 4956 9986 5012 9996
rect 5628 9940 5684 9950
rect 5628 9826 5684 9884
rect 5628 9774 5630 9826
rect 5682 9774 5684 9826
rect 5628 9762 5684 9774
rect 4956 9604 5012 9614
rect 5740 9604 5796 11564
rect 5964 11394 6020 11406
rect 5964 11342 5966 11394
rect 6018 11342 6020 11394
rect 5964 11284 6020 11342
rect 5964 11218 6020 11228
rect 6076 11394 6132 11406
rect 6076 11342 6078 11394
rect 6130 11342 6132 11394
rect 6076 10724 6132 11342
rect 6076 10658 6132 10668
rect 6076 9940 6132 9950
rect 6188 9940 6244 12908
rect 6300 11956 6356 13694
rect 6412 13746 6580 13748
rect 6412 13694 6526 13746
rect 6578 13694 6580 13746
rect 6412 13692 6580 13694
rect 6412 12292 6468 13692
rect 6524 13682 6580 13692
rect 6636 13746 6916 13748
rect 6636 13694 6862 13746
rect 6914 13694 6916 13746
rect 6636 13692 6916 13694
rect 6524 13188 6580 13198
rect 6636 13188 6692 13692
rect 6860 13682 6916 13692
rect 7756 13636 7812 13646
rect 7532 13634 7812 13636
rect 7532 13582 7758 13634
rect 7810 13582 7812 13634
rect 7532 13580 7812 13582
rect 6524 13186 6692 13188
rect 6524 13134 6526 13186
rect 6578 13134 6692 13186
rect 6524 13132 6692 13134
rect 6748 13524 6804 13534
rect 6524 13122 6580 13132
rect 6412 12226 6468 12236
rect 6524 12404 6580 12414
rect 6524 12178 6580 12348
rect 6524 12126 6526 12178
rect 6578 12126 6580 12178
rect 6524 12114 6580 12126
rect 6300 11900 6468 11956
rect 6412 11506 6468 11900
rect 6412 11454 6414 11506
rect 6466 11454 6468 11506
rect 6412 11442 6468 11454
rect 6524 11620 6580 11630
rect 6076 9938 6244 9940
rect 6076 9886 6078 9938
rect 6130 9886 6244 9938
rect 6076 9884 6244 9886
rect 6300 11396 6356 11406
rect 6300 10612 6356 11340
rect 6524 11394 6580 11564
rect 6524 11342 6526 11394
rect 6578 11342 6580 11394
rect 6524 10836 6580 11342
rect 6748 10836 6804 13468
rect 7308 13524 7364 13534
rect 7532 13524 7588 13580
rect 7756 13570 7812 13580
rect 7980 13634 8036 13646
rect 7980 13582 7982 13634
rect 8034 13582 8036 13634
rect 7308 13522 7588 13524
rect 7308 13470 7310 13522
rect 7362 13470 7588 13522
rect 7308 13468 7588 13470
rect 7196 12850 7252 12862
rect 7196 12798 7198 12850
rect 7250 12798 7252 12850
rect 7196 12628 7252 12798
rect 7196 12562 7252 12572
rect 7308 12404 7364 13468
rect 7868 13412 7924 13422
rect 7868 12962 7924 13356
rect 7868 12910 7870 12962
rect 7922 12910 7924 12962
rect 7868 12898 7924 12910
rect 7532 12852 7588 12862
rect 7532 12758 7588 12796
rect 7308 12338 7364 12348
rect 6972 12180 7028 12190
rect 7868 12180 7924 12190
rect 7980 12180 8036 13582
rect 8428 13524 8484 14364
rect 9528 14140 9792 14150
rect 8428 13458 8484 13468
rect 8540 14084 8596 14094
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9528 14074 9792 14084
rect 6972 12178 7588 12180
rect 6972 12126 6974 12178
rect 7026 12126 7588 12178
rect 6972 12124 7588 12126
rect 6972 12114 7028 12124
rect 7084 11956 7140 11966
rect 7140 11900 7252 11956
rect 7084 11890 7140 11900
rect 6860 11620 6916 11630
rect 6860 11526 6916 11564
rect 7084 11396 7140 11406
rect 7084 11302 7140 11340
rect 6524 10770 6580 10780
rect 6636 10780 6804 10836
rect 6076 9874 6132 9884
rect 4844 8820 4900 8830
rect 4844 8726 4900 8764
rect 4956 8484 5012 9548
rect 5404 9548 5796 9604
rect 5964 9826 6020 9838
rect 5964 9774 5966 9826
rect 6018 9774 6020 9826
rect 5292 9268 5348 9278
rect 4956 8418 5012 8428
rect 5068 9266 5348 9268
rect 5068 9214 5294 9266
rect 5346 9214 5348 9266
rect 5068 9212 5348 9214
rect 4732 7422 4734 7474
rect 4786 7422 4788 7474
rect 4172 7250 4228 7262
rect 4172 7198 4174 7250
rect 4226 7198 4228 7250
rect 4172 7140 4228 7198
rect 4172 7074 4228 7084
rect 4732 7028 4788 7422
rect 4732 6962 4788 6972
rect 4844 8146 4900 8158
rect 4844 8094 4846 8146
rect 4898 8094 4900 8146
rect 4844 7364 4900 8094
rect 5068 7700 5124 9212
rect 5292 9202 5348 9212
rect 5404 9266 5460 9548
rect 5404 9214 5406 9266
rect 5458 9214 5460 9266
rect 5404 9202 5460 9214
rect 5852 9268 5908 9278
rect 5516 9156 5572 9166
rect 5516 9062 5572 9100
rect 5180 9042 5236 9054
rect 5180 8990 5182 9042
rect 5234 8990 5236 9042
rect 5180 8036 5236 8990
rect 5370 8652 5634 8662
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5370 8586 5634 8596
rect 5628 8484 5684 8494
rect 5628 8258 5684 8428
rect 5852 8370 5908 9212
rect 5964 8596 6020 9774
rect 6188 9716 6244 9726
rect 5964 8530 6020 8540
rect 6076 9660 6188 9716
rect 6076 8428 6132 9660
rect 6188 9622 6244 9660
rect 6300 9492 6356 10556
rect 6636 10164 6692 10780
rect 6860 10722 6916 10734
rect 6860 10670 6862 10722
rect 6914 10670 6916 10722
rect 6748 10610 6804 10622
rect 6748 10558 6750 10610
rect 6802 10558 6804 10610
rect 6748 10276 6804 10558
rect 6860 10388 6916 10670
rect 7084 10612 7140 10622
rect 7084 10518 7140 10556
rect 6860 10332 7140 10388
rect 6748 10220 7028 10276
rect 6636 10108 6916 10164
rect 5852 8318 5854 8370
rect 5906 8318 5908 8370
rect 5852 8306 5908 8318
rect 5964 8372 6132 8428
rect 6188 9436 6356 9492
rect 5628 8206 5630 8258
rect 5682 8206 5684 8258
rect 5628 8194 5684 8206
rect 5516 8036 5572 8046
rect 5740 8036 5796 8046
rect 5180 8034 5572 8036
rect 5180 7982 5518 8034
rect 5570 7982 5572 8034
rect 5180 7980 5572 7982
rect 5516 7970 5572 7980
rect 5628 7980 5740 8036
rect 5180 7700 5236 7710
rect 5068 7698 5236 7700
rect 5068 7646 5182 7698
rect 5234 7646 5236 7698
rect 5068 7644 5236 7646
rect 5180 7634 5236 7644
rect 5068 7476 5124 7486
rect 4844 6916 4900 7308
rect 4844 6850 4900 6860
rect 4956 7474 5124 7476
rect 4956 7422 5070 7474
rect 5122 7422 5124 7474
rect 4956 7420 5124 7422
rect 4956 6802 5012 7420
rect 5068 7410 5124 7420
rect 5292 7476 5348 7486
rect 5292 7382 5348 7420
rect 5516 7476 5572 7486
rect 5628 7476 5684 7980
rect 5740 7970 5796 7980
rect 5740 7812 5796 7822
rect 5796 7756 5908 7812
rect 5740 7746 5796 7756
rect 5516 7474 5684 7476
rect 5516 7422 5518 7474
rect 5570 7422 5684 7474
rect 5516 7420 5684 7422
rect 5740 7474 5796 7486
rect 5740 7422 5742 7474
rect 5794 7422 5796 7474
rect 5516 7410 5572 7420
rect 5740 7140 5796 7422
rect 5370 7084 5634 7094
rect 4956 6750 4958 6802
rect 5010 6750 5012 6802
rect 4956 6738 5012 6750
rect 5068 7028 5124 7038
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5740 7074 5796 7084
rect 5370 7018 5634 7028
rect 5068 6804 5124 6972
rect 5068 6690 5124 6748
rect 5068 6638 5070 6690
rect 5122 6638 5124 6690
rect 5068 6626 5124 6638
rect 5180 6916 5236 6926
rect 3724 6524 3892 6580
rect 3612 6402 3668 6412
rect 3388 5182 3390 5234
rect 3442 5182 3444 5234
rect 3388 5170 3444 5182
rect 3724 5906 3780 5918
rect 3724 5854 3726 5906
rect 3778 5854 3780 5906
rect 2492 4450 2660 4452
rect 2492 4398 2494 4450
rect 2546 4398 2660 4450
rect 2492 4396 2660 4398
rect 3612 5124 3668 5134
rect 3724 5124 3780 5854
rect 3612 5122 3780 5124
rect 3612 5070 3614 5122
rect 3666 5070 3780 5122
rect 3612 5068 3780 5070
rect 3612 4452 3668 5068
rect 3836 4900 3892 6524
rect 4620 6468 4676 6478
rect 4620 6374 4676 6412
rect 4844 6468 4900 6478
rect 5180 6468 5236 6860
rect 5628 6804 5684 6814
rect 5628 6710 5684 6748
rect 5740 6580 5796 6590
rect 5740 6486 5796 6524
rect 4844 6466 5236 6468
rect 4844 6414 4846 6466
rect 4898 6414 5236 6466
rect 4844 6412 5236 6414
rect 4844 6402 4900 6412
rect 3948 6356 4004 6366
rect 3948 5346 4004 6300
rect 4060 6018 4116 6030
rect 4060 5966 4062 6018
rect 4114 5966 4116 6018
rect 4060 5796 4116 5966
rect 5292 6020 5348 6030
rect 4396 5908 4452 5918
rect 4396 5814 4452 5852
rect 4844 5906 4900 5918
rect 5292 5908 5348 5964
rect 4844 5854 4846 5906
rect 4898 5854 4900 5906
rect 4060 5730 4116 5740
rect 3948 5294 3950 5346
rect 4002 5294 4004 5346
rect 3948 5282 4004 5294
rect 4620 5348 4676 5358
rect 4620 5254 4676 5292
rect 4284 5124 4340 5134
rect 4284 5030 4340 5068
rect 4844 5124 4900 5854
rect 5180 5906 5348 5908
rect 5180 5854 5294 5906
rect 5346 5854 5348 5906
rect 5180 5852 5348 5854
rect 5180 5348 5236 5852
rect 5292 5842 5348 5852
rect 5852 6018 5908 7756
rect 5852 5966 5854 6018
rect 5906 5966 5908 6018
rect 5852 5684 5908 5966
rect 5964 5796 6020 8372
rect 6076 8258 6132 8270
rect 6076 8206 6078 8258
rect 6130 8206 6132 8258
rect 6076 7700 6132 8206
rect 6076 7634 6132 7644
rect 6188 7476 6244 9436
rect 6524 9156 6580 9166
rect 6524 9062 6580 9100
rect 6412 9044 6468 9054
rect 6412 8950 6468 8988
rect 6636 9042 6692 9054
rect 6636 8990 6638 9042
rect 6690 8990 6692 9042
rect 6636 8484 6692 8990
rect 6636 8418 6692 8428
rect 6524 8260 6580 8270
rect 6524 8166 6580 8204
rect 6300 8148 6356 8158
rect 6300 8146 6468 8148
rect 6300 8094 6302 8146
rect 6354 8094 6468 8146
rect 6300 8092 6468 8094
rect 6300 8082 6356 8092
rect 5964 5730 6020 5740
rect 6076 7420 6244 7476
rect 6300 7924 6356 7934
rect 6076 5684 6132 7420
rect 6300 6804 6356 7868
rect 6412 7812 6468 8092
rect 6860 8036 6916 10108
rect 6972 8708 7028 10220
rect 7084 9828 7140 10332
rect 7084 9762 7140 9772
rect 7084 9268 7140 9278
rect 7084 9042 7140 9212
rect 7084 8990 7086 9042
rect 7138 8990 7140 9042
rect 7084 8820 7140 8990
rect 7084 8754 7140 8764
rect 6972 8642 7028 8652
rect 7196 8428 7252 11900
rect 7532 11394 7588 12124
rect 7532 11342 7534 11394
rect 7586 11342 7588 11394
rect 7420 11284 7476 11294
rect 7420 11190 7476 11228
rect 7308 11170 7364 11182
rect 7308 11118 7310 11170
rect 7362 11118 7364 11170
rect 7308 11060 7364 11118
rect 7308 11004 7476 11060
rect 7308 10836 7364 10846
rect 7308 9268 7364 10780
rect 7420 10164 7476 11004
rect 7420 10098 7476 10108
rect 7532 10052 7588 11342
rect 7644 12178 8036 12180
rect 7644 12126 7870 12178
rect 7922 12126 8036 12178
rect 7644 12124 8036 12126
rect 8316 12628 8372 12638
rect 7644 10836 7700 12124
rect 7868 12114 7924 12124
rect 8204 12068 8260 12078
rect 7644 10742 7700 10780
rect 7980 11396 8036 11406
rect 7532 9986 7588 9996
rect 7980 10050 8036 11340
rect 7980 9998 7982 10050
rect 8034 9998 8036 10050
rect 7980 9986 8036 9998
rect 8204 10612 8260 12012
rect 7308 9202 7364 9212
rect 7868 9828 7924 9838
rect 8204 9828 8260 10556
rect 7868 9266 7924 9772
rect 7980 9772 8260 9828
rect 7980 9714 8036 9772
rect 7980 9662 7982 9714
rect 8034 9662 8036 9714
rect 7980 9650 8036 9662
rect 8092 9658 8148 9670
rect 7868 9214 7870 9266
rect 7922 9214 7924 9266
rect 7868 9202 7924 9214
rect 8092 9606 8094 9658
rect 8146 9606 8148 9658
rect 7644 9042 7700 9054
rect 7644 8990 7646 9042
rect 7698 8990 7700 9042
rect 7644 8708 7700 8990
rect 7756 9044 7812 9054
rect 7756 8950 7812 8988
rect 7644 8642 7700 8652
rect 7980 8932 8036 8942
rect 6972 8372 7028 8382
rect 7196 8372 7476 8428
rect 6972 8258 7028 8316
rect 6972 8206 6974 8258
rect 7026 8206 7028 8258
rect 6972 8194 7028 8206
rect 7196 8148 7252 8158
rect 7196 8054 7252 8092
rect 7420 8148 7476 8372
rect 7420 8082 7476 8092
rect 7532 8146 7588 8158
rect 7532 8094 7534 8146
rect 7586 8094 7588 8146
rect 6860 7980 7028 8036
rect 6412 7756 6804 7812
rect 6748 7698 6804 7756
rect 6748 7646 6750 7698
rect 6802 7646 6804 7698
rect 6748 7634 6804 7646
rect 6636 7474 6692 7486
rect 6636 7422 6638 7474
rect 6690 7422 6692 7474
rect 6636 7140 6692 7422
rect 6860 7476 6916 7486
rect 6860 7382 6916 7420
rect 6972 7252 7028 7980
rect 7084 8034 7140 8046
rect 7084 7982 7086 8034
rect 7138 7982 7140 8034
rect 7084 7924 7140 7982
rect 7308 8034 7364 8046
rect 7308 7982 7310 8034
rect 7362 7982 7364 8034
rect 7196 7924 7252 7934
rect 7084 7868 7196 7924
rect 7196 7858 7252 7868
rect 7308 7812 7364 7982
rect 7532 7924 7588 8094
rect 7532 7868 7812 7924
rect 7364 7756 7700 7812
rect 7308 7746 7364 7756
rect 7644 7698 7700 7756
rect 7644 7646 7646 7698
rect 7698 7646 7700 7698
rect 7644 7634 7700 7646
rect 6636 7074 6692 7084
rect 6748 7196 7028 7252
rect 7308 7474 7364 7486
rect 7756 7476 7812 7868
rect 7308 7422 7310 7474
rect 7362 7422 7364 7474
rect 6300 6748 6692 6804
rect 6188 6692 6244 6702
rect 6188 6690 6356 6692
rect 6188 6638 6190 6690
rect 6242 6638 6356 6690
rect 6188 6636 6356 6638
rect 6188 6626 6244 6636
rect 6188 6468 6244 6478
rect 6188 6374 6244 6412
rect 6300 6132 6356 6636
rect 6524 6578 6580 6590
rect 6524 6526 6526 6578
rect 6578 6526 6580 6578
rect 6188 6076 6356 6132
rect 6412 6468 6468 6478
rect 6188 6020 6244 6076
rect 6412 6020 6468 6412
rect 6524 6244 6580 6526
rect 6524 6178 6580 6188
rect 6188 5954 6244 5964
rect 6300 5964 6468 6020
rect 6524 6018 6580 6030
rect 6524 5966 6526 6018
rect 6578 5966 6580 6018
rect 6300 5906 6356 5964
rect 6300 5854 6302 5906
rect 6354 5854 6356 5906
rect 6300 5842 6356 5854
rect 6412 5794 6468 5806
rect 6412 5742 6414 5794
rect 6466 5742 6468 5794
rect 6076 5628 6356 5684
rect 5852 5618 5908 5628
rect 5370 5516 5634 5526
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5370 5450 5634 5460
rect 4844 5030 4900 5068
rect 5068 5236 5124 5246
rect 5068 5010 5124 5180
rect 5068 4958 5070 5010
rect 5122 4958 5124 5010
rect 5068 4946 5124 4958
rect 4284 4900 4340 4910
rect 3836 4898 4340 4900
rect 3836 4846 4286 4898
rect 4338 4846 4340 4898
rect 3836 4844 4340 4846
rect 4284 4834 4340 4844
rect 4732 4564 4788 4574
rect 4732 4470 4788 4508
rect 2492 4386 2548 4396
rect 3612 4386 3668 4396
rect 1820 4340 1876 4350
rect 1820 4246 1876 4284
rect 1596 4162 1652 4172
rect 3612 4228 3668 4238
rect 3612 800 3668 4172
rect 5180 3668 5236 5292
rect 6188 5236 6244 5246
rect 5964 5124 6020 5134
rect 5740 4340 5796 4350
rect 5370 3948 5634 3958
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5370 3882 5634 3892
rect 5180 3602 5236 3612
rect 5740 3666 5796 4284
rect 5852 4116 5908 4126
rect 5964 4116 6020 5068
rect 5852 4114 6020 4116
rect 5852 4062 5854 4114
rect 5906 4062 6020 4114
rect 5852 4060 6020 4062
rect 5852 4050 5908 4060
rect 5740 3614 5742 3666
rect 5794 3614 5796 3666
rect 5740 3602 5796 3614
rect 5964 3332 6020 4060
rect 6076 5012 6132 5022
rect 6076 3554 6132 4956
rect 6188 5010 6244 5180
rect 6188 4958 6190 5010
rect 6242 4958 6244 5010
rect 6188 4946 6244 4958
rect 6300 4898 6356 5628
rect 6300 4846 6302 4898
rect 6354 4846 6356 4898
rect 6300 4834 6356 4846
rect 6412 4450 6468 5742
rect 6412 4398 6414 4450
rect 6466 4398 6468 4450
rect 6412 4116 6468 4398
rect 6412 4050 6468 4060
rect 6524 3892 6580 5966
rect 6076 3502 6078 3554
rect 6130 3502 6132 3554
rect 6076 3490 6132 3502
rect 6412 3836 6580 3892
rect 6300 3444 6356 3454
rect 6188 3442 6356 3444
rect 6188 3390 6302 3442
rect 6354 3390 6356 3442
rect 6188 3388 6356 3390
rect 6188 3332 6244 3388
rect 6300 3378 6356 3388
rect 5964 3276 6244 3332
rect 6412 2996 6468 3836
rect 6636 3556 6692 6748
rect 6748 4340 6804 7196
rect 7084 6244 7140 6254
rect 6860 5012 6916 5022
rect 6860 4562 6916 4956
rect 6860 4510 6862 4562
rect 6914 4510 6916 4562
rect 6860 4498 6916 4510
rect 6972 4452 7028 4462
rect 6972 4358 7028 4396
rect 6748 4274 6804 4284
rect 6860 4228 6916 4238
rect 6860 4114 6916 4172
rect 6860 4062 6862 4114
rect 6914 4062 6916 4114
rect 6860 4050 6916 4062
rect 6972 4116 7028 4126
rect 6524 3500 6692 3556
rect 6748 3668 6804 3678
rect 6748 3554 6804 3612
rect 6748 3502 6750 3554
rect 6802 3502 6804 3554
rect 6524 3442 6580 3500
rect 6748 3490 6804 3502
rect 6972 3554 7028 4060
rect 7084 3778 7140 6188
rect 7308 5012 7364 7422
rect 7644 7420 7812 7476
rect 7868 7476 7924 7486
rect 7308 4918 7364 4956
rect 7420 5906 7476 5918
rect 7420 5854 7422 5906
rect 7474 5854 7476 5906
rect 7420 5122 7476 5854
rect 7644 5908 7700 7420
rect 7868 6692 7924 7420
rect 7644 5814 7700 5852
rect 7756 6636 7924 6692
rect 7420 5070 7422 5122
rect 7474 5070 7476 5122
rect 7084 3726 7086 3778
rect 7138 3726 7140 3778
rect 7084 3714 7140 3726
rect 7420 4338 7476 5070
rect 7756 5012 7812 6636
rect 7868 6468 7924 6478
rect 7868 6374 7924 6412
rect 7980 6466 8036 8876
rect 8092 8484 8148 9606
rect 8316 9042 8372 12572
rect 8540 11620 8596 14028
rect 9772 13972 9828 13982
rect 9548 13748 9604 13758
rect 9548 13524 9604 13692
rect 9548 13458 9604 13468
rect 9772 13076 9828 13916
rect 11676 13972 11732 16716
rect 12348 16772 12404 16830
rect 12908 16884 12964 16894
rect 12348 16706 12404 16716
rect 12796 16770 12852 16782
rect 12796 16718 12798 16770
rect 12850 16718 12852 16770
rect 12684 16660 12740 16670
rect 12460 16658 12740 16660
rect 12460 16606 12686 16658
rect 12738 16606 12740 16658
rect 12460 16604 12740 16606
rect 12460 15876 12516 16604
rect 12684 16594 12740 16604
rect 12796 16212 12852 16718
rect 12796 16146 12852 16156
rect 12908 16210 12964 16828
rect 12908 16158 12910 16210
rect 12962 16158 12964 16210
rect 12908 16146 12964 16158
rect 13468 16884 13524 20076
rect 13580 20066 13636 20076
rect 14028 20132 14084 20142
rect 14028 20038 14084 20076
rect 14252 20020 14308 20030
rect 14588 20020 14644 23884
rect 14700 21810 14756 23996
rect 14924 23986 14980 23996
rect 15036 24164 15092 24174
rect 15036 23940 15092 24108
rect 15036 23884 15204 23940
rect 14924 23828 14980 23838
rect 14812 23492 14868 23502
rect 14812 23378 14868 23436
rect 14812 23326 14814 23378
rect 14866 23326 14868 23378
rect 14812 23314 14868 23326
rect 14700 21758 14702 21810
rect 14754 21758 14756 21810
rect 14700 21588 14756 21758
rect 14924 21810 14980 23772
rect 14924 21758 14926 21810
rect 14978 21758 14980 21810
rect 14924 21746 14980 21758
rect 15036 23156 15092 23166
rect 14812 21700 14868 21710
rect 14812 21606 14868 21644
rect 14700 21522 14756 21532
rect 15036 20132 15092 23100
rect 15148 21586 15204 23884
rect 15372 23604 15428 23614
rect 15372 23268 15428 23548
rect 15372 23154 15428 23212
rect 15372 23102 15374 23154
rect 15426 23102 15428 23154
rect 15372 23090 15428 23102
rect 15484 23156 15540 25116
rect 15708 24834 15764 26236
rect 15820 26290 15876 26460
rect 15820 26238 15822 26290
rect 15874 26238 15876 26290
rect 15820 26226 15876 26238
rect 15932 26514 16324 26516
rect 15932 26462 16270 26514
rect 16322 26462 16324 26514
rect 15932 26460 16324 26462
rect 15820 25508 15876 25518
rect 15932 25508 15988 26460
rect 16268 26450 16324 26460
rect 16156 26292 16212 26302
rect 15820 25506 15988 25508
rect 15820 25454 15822 25506
rect 15874 25454 15988 25506
rect 15820 25452 15988 25454
rect 16044 26290 16212 26292
rect 16044 26238 16158 26290
rect 16210 26238 16212 26290
rect 16044 26236 16212 26238
rect 15820 25442 15876 25452
rect 16044 25396 16100 26236
rect 16156 26226 16212 26236
rect 16380 26292 16436 27132
rect 17164 27188 17220 27198
rect 17164 27094 17220 27132
rect 17612 27074 17668 27086
rect 17612 27022 17614 27074
rect 17666 27022 17668 27074
rect 16380 26198 16436 26236
rect 16604 26402 16660 26414
rect 16604 26350 16606 26402
rect 16658 26350 16660 26402
rect 16604 25844 16660 26350
rect 16156 25396 16212 25406
rect 16044 25340 16156 25396
rect 16156 25302 16212 25340
rect 16604 25396 16660 25788
rect 17612 26180 17668 27022
rect 17724 27076 17780 27086
rect 17724 26852 17780 27020
rect 17724 26292 17780 26796
rect 18284 26962 18340 26974
rect 18284 26910 18286 26962
rect 18338 26910 18340 26962
rect 17844 26684 18108 26694
rect 17900 26628 17948 26684
rect 18004 26628 18052 26684
rect 17844 26618 18108 26628
rect 18060 26516 18116 26526
rect 18284 26516 18340 26910
rect 18060 26514 18340 26516
rect 18060 26462 18062 26514
rect 18114 26462 18340 26514
rect 18060 26460 18340 26462
rect 18956 26628 19012 26638
rect 18956 26514 19012 26572
rect 18956 26462 18958 26514
rect 19010 26462 19012 26514
rect 18060 26450 18116 26460
rect 18956 26450 19012 26462
rect 17836 26292 17892 26302
rect 17724 26290 17892 26292
rect 17724 26238 17838 26290
rect 17890 26238 17892 26290
rect 17724 26236 17892 26238
rect 16604 25394 17332 25396
rect 16604 25342 16606 25394
rect 16658 25342 17332 25394
rect 16604 25340 17332 25342
rect 16604 25330 16660 25340
rect 16268 25284 16324 25294
rect 16268 25190 16324 25228
rect 16380 25282 16436 25294
rect 16380 25230 16382 25282
rect 16434 25230 16436 25282
rect 16380 24948 16436 25230
rect 16380 24882 16436 24892
rect 15708 24782 15710 24834
rect 15762 24782 15764 24834
rect 15708 24770 15764 24782
rect 15596 24498 15652 24510
rect 15596 24446 15598 24498
rect 15650 24446 15652 24498
rect 15596 23940 15652 24446
rect 15596 23874 15652 23884
rect 15932 23828 15988 23838
rect 15820 23492 15876 23502
rect 15820 23378 15876 23436
rect 15820 23326 15822 23378
rect 15874 23326 15876 23378
rect 15820 23314 15876 23326
rect 15932 23378 15988 23772
rect 17164 23828 17220 23838
rect 17164 23734 17220 23772
rect 15932 23326 15934 23378
rect 15986 23326 15988 23378
rect 15932 23314 15988 23326
rect 16044 23380 16100 23390
rect 16044 23286 16100 23324
rect 15596 23156 15652 23166
rect 15484 23100 15596 23156
rect 15596 22258 15652 23100
rect 15596 22206 15598 22258
rect 15650 22206 15652 22258
rect 15148 21534 15150 21586
rect 15202 21534 15204 21586
rect 15148 21522 15204 21534
rect 15484 21586 15540 21598
rect 15484 21534 15486 21586
rect 15538 21534 15540 21586
rect 15372 21476 15428 21486
rect 15372 21382 15428 21420
rect 15484 21028 15540 21534
rect 15484 20962 15540 20972
rect 14924 20130 15092 20132
rect 14924 20078 15038 20130
rect 15090 20078 15092 20130
rect 14924 20076 15092 20078
rect 14812 20020 14868 20030
rect 14588 20018 14868 20020
rect 14588 19966 14814 20018
rect 14866 19966 14868 20018
rect 14588 19964 14868 19966
rect 14252 19926 14308 19964
rect 14812 19908 14868 19964
rect 14812 19842 14868 19852
rect 13686 19628 13950 19638
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13686 19562 13950 19572
rect 14588 19124 14644 19134
rect 14028 18452 14084 18462
rect 14028 18358 14084 18396
rect 13686 18060 13950 18070
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13686 17994 13950 18004
rect 14364 17556 14420 17566
rect 14364 17106 14420 17500
rect 14364 17054 14366 17106
rect 14418 17054 14420 17106
rect 14140 16994 14196 17006
rect 14140 16942 14142 16994
rect 14194 16942 14196 16994
rect 13580 16884 13636 16894
rect 13468 16882 13636 16884
rect 13468 16830 13582 16882
rect 13634 16830 13636 16882
rect 13468 16828 13636 16830
rect 13468 16100 13524 16828
rect 13580 16818 13636 16828
rect 13916 16882 13972 16894
rect 13916 16830 13918 16882
rect 13970 16830 13972 16882
rect 13916 16660 13972 16830
rect 14140 16884 14196 16942
rect 14140 16818 14196 16828
rect 14028 16772 14084 16782
rect 14028 16678 14084 16716
rect 13916 16594 13972 16604
rect 13686 16492 13950 16502
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13686 16426 13950 16436
rect 13692 16212 13748 16222
rect 13692 16118 13748 16156
rect 13468 16044 13636 16100
rect 13580 15988 13636 16044
rect 13804 16098 13860 16110
rect 13804 16046 13806 16098
rect 13858 16046 13860 16098
rect 13804 15988 13860 16046
rect 13580 15932 13860 15988
rect 14140 15988 14196 15998
rect 14140 15894 14196 15932
rect 11900 15820 12516 15876
rect 14252 15874 14308 15886
rect 14252 15822 14254 15874
rect 14306 15822 14308 15874
rect 11900 15426 11956 15820
rect 11900 15374 11902 15426
rect 11954 15374 11956 15426
rect 11900 15362 11956 15374
rect 14028 15428 14084 15438
rect 14252 15428 14308 15822
rect 14364 15876 14420 17054
rect 14476 15876 14532 15886
rect 14364 15874 14532 15876
rect 14364 15822 14478 15874
rect 14530 15822 14532 15874
rect 14364 15820 14532 15822
rect 14476 15810 14532 15820
rect 14084 15372 14308 15428
rect 13468 15316 13524 15326
rect 11676 13906 11732 13916
rect 12684 14530 12740 14542
rect 12684 14478 12686 14530
rect 12738 14478 12740 14530
rect 12684 14420 12740 14478
rect 9996 13858 10052 13870
rect 9996 13806 9998 13858
rect 10050 13806 10052 13858
rect 9996 13636 10052 13806
rect 10108 13860 10164 13870
rect 10108 13766 10164 13804
rect 10892 13858 10948 13870
rect 10892 13806 10894 13858
rect 10946 13806 10948 13858
rect 10892 13748 10948 13806
rect 11116 13860 11172 13870
rect 11116 13766 11172 13804
rect 11340 13748 11396 13758
rect 10892 13682 10948 13692
rect 11228 13746 11396 13748
rect 11228 13694 11342 13746
rect 11394 13694 11396 13746
rect 11228 13692 11396 13694
rect 10220 13636 10276 13646
rect 9996 13570 10052 13580
rect 10108 13634 10276 13636
rect 10108 13582 10222 13634
rect 10274 13582 10276 13634
rect 10108 13580 10276 13582
rect 9772 13010 9828 13020
rect 8652 12852 8708 12862
rect 10108 12852 10164 13580
rect 10220 13570 10276 13580
rect 10780 13636 10836 13646
rect 10780 13074 10836 13580
rect 10780 13022 10782 13074
rect 10834 13022 10836 13074
rect 10780 13010 10836 13022
rect 11228 13074 11284 13692
rect 11340 13682 11396 13692
rect 11900 13636 11956 13646
rect 11900 13542 11956 13580
rect 11788 13524 11844 13534
rect 11228 13022 11230 13074
rect 11282 13022 11284 13074
rect 11228 13010 11284 13022
rect 11676 13522 11844 13524
rect 11676 13470 11790 13522
rect 11842 13470 11844 13522
rect 11676 13468 11844 13470
rect 11676 12962 11732 13468
rect 11788 13458 11844 13468
rect 12572 13412 12628 13422
rect 12124 13076 12180 13086
rect 12124 12982 12180 13020
rect 12572 13074 12628 13356
rect 12572 13022 12574 13074
rect 12626 13022 12628 13074
rect 12572 13010 12628 13022
rect 11676 12910 11678 12962
rect 11730 12910 11732 12962
rect 11676 12898 11732 12910
rect 8652 12850 8820 12852
rect 8652 12798 8654 12850
rect 8706 12798 8820 12850
rect 8652 12796 8820 12798
rect 8652 12786 8708 12796
rect 8652 12628 8708 12638
rect 8652 12290 8708 12572
rect 8652 12238 8654 12290
rect 8706 12238 8708 12290
rect 8652 12226 8708 12238
rect 8764 12292 8820 12796
rect 9528 12572 9792 12582
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9528 12506 9792 12516
rect 8988 12292 9044 12302
rect 10108 12292 10164 12796
rect 11116 12740 11172 12750
rect 11340 12740 11396 12750
rect 11116 12738 11284 12740
rect 11116 12686 11118 12738
rect 11170 12686 11284 12738
rect 11116 12684 11284 12686
rect 11116 12674 11172 12684
rect 8764 12236 8988 12292
rect 8988 12198 9044 12236
rect 9884 12236 10164 12292
rect 10668 12292 10724 12302
rect 8540 11526 8596 11564
rect 9212 11508 9268 11518
rect 9100 11452 9212 11508
rect 8764 11394 8820 11406
rect 8764 11342 8766 11394
rect 8818 11342 8820 11394
rect 8428 11282 8484 11294
rect 8428 11230 8430 11282
rect 8482 11230 8484 11282
rect 8428 10610 8484 11230
rect 8428 10558 8430 10610
rect 8482 10558 8484 10610
rect 8428 10546 8484 10558
rect 8652 10386 8708 10398
rect 8652 10334 8654 10386
rect 8706 10334 8708 10386
rect 8652 9940 8708 10334
rect 8764 10388 8820 11342
rect 8876 11394 8932 11406
rect 8876 11342 8878 11394
rect 8930 11342 8932 11394
rect 8876 10948 8932 11342
rect 8876 10882 8932 10892
rect 8988 11284 9044 11294
rect 8876 10724 8932 10734
rect 8876 10610 8932 10668
rect 8988 10722 9044 11228
rect 8988 10670 8990 10722
rect 9042 10670 9044 10722
rect 8988 10658 9044 10670
rect 8876 10558 8878 10610
rect 8930 10558 8932 10610
rect 8876 10546 8932 10558
rect 8764 10322 8820 10332
rect 8876 9940 8932 9950
rect 8652 9938 8932 9940
rect 8652 9886 8878 9938
rect 8930 9886 8932 9938
rect 8652 9884 8932 9886
rect 8876 9874 8932 9884
rect 8764 9716 8820 9726
rect 8764 9622 8820 9660
rect 8988 9714 9044 9726
rect 8988 9662 8990 9714
rect 9042 9662 9044 9714
rect 8988 9604 9044 9662
rect 8988 9538 9044 9548
rect 8988 9156 9044 9166
rect 8316 8990 8318 9042
rect 8370 8990 8372 9042
rect 8316 8978 8372 8990
rect 8876 9100 8988 9156
rect 8092 8418 8148 8428
rect 7980 6414 7982 6466
rect 8034 6414 8036 6466
rect 7980 6402 8036 6414
rect 8092 8148 8148 8158
rect 7868 6132 7924 6142
rect 7868 6038 7924 6076
rect 7980 6132 8036 6142
rect 8092 6132 8148 8092
rect 8652 8146 8708 8158
rect 8652 8094 8654 8146
rect 8706 8094 8708 8146
rect 8428 8036 8484 8046
rect 8652 8036 8708 8094
rect 8764 8148 8820 8158
rect 8764 8054 8820 8092
rect 8876 8146 8932 9100
rect 8988 9090 9044 9100
rect 8876 8094 8878 8146
rect 8930 8094 8932 8146
rect 8876 8082 8932 8094
rect 8988 8484 9044 8494
rect 8316 8034 8484 8036
rect 8316 7982 8430 8034
rect 8482 7982 8484 8034
rect 8316 7980 8484 7982
rect 8316 7362 8372 7980
rect 8428 7970 8484 7980
rect 8540 7980 8708 8036
rect 8540 7812 8596 7980
rect 8316 7310 8318 7362
rect 8370 7310 8372 7362
rect 8316 7298 8372 7310
rect 8428 7756 8596 7812
rect 8876 7924 8932 7934
rect 7980 6130 8148 6132
rect 7980 6078 7982 6130
rect 8034 6078 8148 6130
rect 7980 6076 8148 6078
rect 8204 6690 8260 6702
rect 8204 6638 8206 6690
rect 8258 6638 8260 6690
rect 8204 6580 8260 6638
rect 8204 6132 8260 6524
rect 7980 6066 8036 6076
rect 8204 6066 8260 6076
rect 8316 6468 8372 6478
rect 8204 5906 8260 5918
rect 8204 5854 8206 5906
rect 8258 5854 8260 5906
rect 8204 5796 8260 5854
rect 8204 5730 8260 5740
rect 8092 5684 8148 5694
rect 7980 5460 8036 5470
rect 7868 5012 7924 5022
rect 7756 5010 7924 5012
rect 7756 4958 7870 5010
rect 7922 4958 7924 5010
rect 7756 4956 7924 4958
rect 7644 4900 7700 4910
rect 7644 4806 7700 4844
rect 7644 4564 7700 4574
rect 7644 4470 7700 4508
rect 7420 4286 7422 4338
rect 7474 4286 7476 4338
rect 7420 3668 7476 4286
rect 7868 4116 7924 4956
rect 7980 4562 8036 5404
rect 8092 5122 8148 5628
rect 8316 5348 8372 6412
rect 8428 6020 8484 7756
rect 8876 7586 8932 7868
rect 8876 7534 8878 7586
rect 8930 7534 8932 7586
rect 8764 7474 8820 7486
rect 8764 7422 8766 7474
rect 8818 7422 8820 7474
rect 8764 7252 8820 7422
rect 8876 7476 8932 7534
rect 8876 7410 8932 7420
rect 8764 7196 8932 7252
rect 8428 5926 8484 5964
rect 8540 6690 8596 6702
rect 8540 6638 8542 6690
rect 8594 6638 8596 6690
rect 8540 6244 8596 6638
rect 8540 5572 8596 6188
rect 8764 6018 8820 6030
rect 8764 5966 8766 6018
rect 8818 5966 8820 6018
rect 8540 5506 8596 5516
rect 8652 5906 8708 5918
rect 8652 5854 8654 5906
rect 8706 5854 8708 5906
rect 8428 5348 8484 5358
rect 8316 5292 8428 5348
rect 8092 5070 8094 5122
rect 8146 5070 8148 5122
rect 8092 5058 8148 5070
rect 7980 4510 7982 4562
rect 8034 4510 8036 4562
rect 7980 4498 8036 4510
rect 8204 5012 8260 5022
rect 7868 4050 7924 4060
rect 8204 4338 8260 4956
rect 8204 4286 8206 4338
rect 8258 4286 8260 4338
rect 8092 3668 8148 3678
rect 7420 3666 8148 3668
rect 7420 3614 8094 3666
rect 8146 3614 8148 3666
rect 7420 3612 8148 3614
rect 8092 3602 8148 3612
rect 6972 3502 6974 3554
rect 7026 3502 7028 3554
rect 6972 3490 7028 3502
rect 6524 3390 6526 3442
rect 6578 3390 6580 3442
rect 6524 3378 6580 3390
rect 8204 3332 8260 4286
rect 8428 3666 8484 5292
rect 8652 5236 8708 5854
rect 8764 5908 8820 5966
rect 8764 5842 8820 5852
rect 8876 5796 8932 7196
rect 8876 5730 8932 5740
rect 8988 5794 9044 8428
rect 9100 8372 9156 11452
rect 9212 11442 9268 11452
rect 9884 11394 9940 12236
rect 10668 12198 10724 12236
rect 10220 12180 10276 12190
rect 9884 11342 9886 11394
rect 9938 11342 9940 11394
rect 9884 11330 9940 11342
rect 10108 12178 10276 12180
rect 10108 12126 10222 12178
rect 10274 12126 10276 12178
rect 10108 12124 10276 12126
rect 9324 11282 9380 11294
rect 9324 11230 9326 11282
rect 9378 11230 9380 11282
rect 9324 11172 9380 11230
rect 9324 11106 9380 11116
rect 9996 11172 10052 11182
rect 9528 11004 9792 11014
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9528 10938 9792 10948
rect 9436 10612 9492 10622
rect 9436 10518 9492 10556
rect 9884 10612 9940 10622
rect 9884 10518 9940 10556
rect 9996 10610 10052 11116
rect 9996 10558 9998 10610
rect 10050 10558 10052 10610
rect 9996 10546 10052 10558
rect 10108 10276 10164 12124
rect 10220 12114 10276 12124
rect 10780 12178 10836 12190
rect 10780 12126 10782 12178
rect 10834 12126 10836 12178
rect 10444 12066 10500 12078
rect 10444 12014 10446 12066
rect 10498 12014 10500 12066
rect 10444 11620 10500 12014
rect 10444 11554 10500 11564
rect 10668 11508 10724 11518
rect 10780 11508 10836 12126
rect 11228 11732 11284 12684
rect 11340 12646 11396 12684
rect 12012 12740 12068 12750
rect 12012 12646 12068 12684
rect 12684 12178 12740 14364
rect 12684 12126 12686 12178
rect 12738 12126 12740 12178
rect 12684 12114 12740 12126
rect 13132 13748 13188 13758
rect 13132 12740 13188 13692
rect 11228 11676 11732 11732
rect 10668 11506 10836 11508
rect 10668 11454 10670 11506
rect 10722 11454 10836 11506
rect 10668 11452 10836 11454
rect 10892 11508 10948 11518
rect 10668 11442 10724 11452
rect 10444 11396 10500 11406
rect 10444 11302 10500 11340
rect 10892 11394 10948 11452
rect 11340 11508 11396 11518
rect 11340 11414 11396 11452
rect 10892 11342 10894 11394
rect 10946 11342 10948 11394
rect 10892 11330 10948 11342
rect 10220 11282 10276 11294
rect 10220 11230 10222 11282
rect 10274 11230 10276 11282
rect 10220 10724 10276 11230
rect 11116 11284 11172 11294
rect 11116 11190 11172 11228
rect 10444 11172 10500 11182
rect 10332 11116 10444 11172
rect 10332 10834 10388 11116
rect 10444 11106 10500 11116
rect 11340 11172 11396 11182
rect 11340 11078 11396 11116
rect 10892 10836 10948 10846
rect 10332 10782 10334 10834
rect 10386 10782 10388 10834
rect 10332 10770 10388 10782
rect 10444 10834 10948 10836
rect 10444 10782 10894 10834
rect 10946 10782 10948 10834
rect 10444 10780 10948 10782
rect 10220 10658 10276 10668
rect 10444 10722 10500 10780
rect 10892 10770 10948 10780
rect 11228 10836 11284 10846
rect 10444 10670 10446 10722
rect 10498 10670 10500 10722
rect 10444 10658 10500 10670
rect 10780 10610 10836 10622
rect 10780 10558 10782 10610
rect 10834 10558 10836 10610
rect 10220 10500 10276 10510
rect 10220 10406 10276 10444
rect 10108 10220 10388 10276
rect 9212 10052 9268 10062
rect 9212 9156 9268 9996
rect 9548 9828 9604 9838
rect 9548 9734 9604 9772
rect 9996 9714 10052 9726
rect 9996 9662 9998 9714
rect 10050 9662 10052 9714
rect 9528 9436 9792 9446
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9528 9370 9792 9380
rect 9996 9380 10052 9662
rect 10332 9714 10388 10220
rect 10556 9940 10612 9950
rect 10332 9662 10334 9714
rect 10386 9662 10388 9714
rect 10332 9650 10388 9662
rect 10444 9938 10612 9940
rect 10444 9886 10558 9938
rect 10610 9886 10612 9938
rect 10444 9884 10612 9886
rect 10108 9602 10164 9614
rect 10108 9550 10110 9602
rect 10162 9550 10164 9602
rect 10108 9492 10164 9550
rect 10444 9492 10500 9884
rect 10556 9874 10612 9884
rect 10668 9714 10724 9726
rect 10668 9662 10670 9714
rect 10722 9662 10724 9714
rect 10556 9604 10612 9614
rect 10668 9604 10724 9662
rect 10612 9548 10724 9604
rect 10556 9538 10612 9548
rect 10108 9436 10500 9492
rect 9996 9324 10388 9380
rect 9772 9212 10164 9268
rect 9212 9090 9268 9100
rect 9548 9154 9604 9166
rect 9548 9102 9550 9154
rect 9602 9102 9604 9154
rect 9548 8708 9604 9102
rect 9772 9154 9828 9212
rect 9772 9102 9774 9154
rect 9826 9102 9828 9154
rect 9772 9090 9828 9102
rect 9996 9044 10052 9054
rect 9996 8950 10052 8988
rect 10108 8820 10164 9212
rect 10220 9156 10276 9166
rect 10220 9042 10276 9100
rect 10220 8990 10222 9042
rect 10274 8990 10276 9042
rect 10220 8978 10276 8990
rect 10332 8930 10388 9324
rect 10668 9266 10724 9548
rect 10668 9214 10670 9266
rect 10722 9214 10724 9266
rect 10668 9202 10724 9214
rect 10332 8878 10334 8930
rect 10386 8878 10388 8930
rect 10332 8866 10388 8878
rect 9548 8642 9604 8652
rect 9996 8764 10164 8820
rect 9212 8372 9268 8382
rect 9100 8370 9268 8372
rect 9100 8318 9214 8370
rect 9266 8318 9268 8370
rect 9100 8316 9268 8318
rect 9212 8306 9268 8316
rect 9884 8260 9940 8270
rect 9884 8166 9940 8204
rect 9548 8146 9604 8158
rect 9548 8094 9550 8146
rect 9602 8094 9604 8146
rect 9548 8036 9604 8094
rect 9548 7970 9604 7980
rect 9884 8036 9940 8046
rect 9884 7942 9940 7980
rect 9528 7868 9792 7878
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9528 7802 9792 7812
rect 9772 7700 9828 7710
rect 9772 7642 9828 7644
rect 9436 7588 9492 7598
rect 9436 7494 9492 7532
rect 9660 7586 9716 7598
rect 9660 7534 9662 7586
rect 9714 7534 9716 7586
rect 9772 7590 9774 7642
rect 9826 7590 9828 7642
rect 9772 7578 9828 7590
rect 9660 7476 9716 7534
rect 9884 7476 9940 7486
rect 9996 7476 10052 8764
rect 10668 8596 10724 8606
rect 10108 8372 10164 8382
rect 10164 8316 10276 8372
rect 10108 8306 10164 8316
rect 10108 8146 10164 8158
rect 10108 8094 10110 8146
rect 10162 8094 10164 8146
rect 10108 7588 10164 8094
rect 10108 7522 10164 7532
rect 9660 7420 9828 7476
rect 9660 6804 9716 6814
rect 9660 6710 9716 6748
rect 9100 6692 9156 6702
rect 9100 6578 9156 6636
rect 9772 6692 9828 7420
rect 9940 7420 10052 7476
rect 9884 7410 9940 7420
rect 9772 6598 9828 6636
rect 9884 7252 9940 7262
rect 9100 6526 9102 6578
rect 9154 6526 9156 6578
rect 9100 6514 9156 6526
rect 9548 6468 9604 6478
rect 9324 6466 9604 6468
rect 9324 6414 9550 6466
rect 9602 6414 9604 6466
rect 9324 6412 9604 6414
rect 9324 5908 9380 6412
rect 9548 6402 9604 6412
rect 9528 6300 9792 6310
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9528 6234 9792 6244
rect 9660 6132 9716 6142
rect 9884 6132 9940 7196
rect 10220 6916 10276 8316
rect 10108 6860 10276 6916
rect 10444 8146 10500 8158
rect 10444 8094 10446 8146
rect 10498 8094 10500 8146
rect 10444 7364 10500 8094
rect 9660 6130 9940 6132
rect 9660 6078 9662 6130
rect 9714 6078 9940 6130
rect 9660 6076 9940 6078
rect 9996 6580 10052 6590
rect 9660 6066 9716 6076
rect 9324 5842 9380 5852
rect 9996 5906 10052 6524
rect 9996 5854 9998 5906
rect 10050 5854 10052 5906
rect 9996 5842 10052 5854
rect 8988 5742 8990 5794
rect 9042 5742 9044 5794
rect 8988 5730 9044 5742
rect 8652 5170 8708 5180
rect 9324 5684 9380 5694
rect 10108 5684 10164 6860
rect 10444 6802 10500 7308
rect 10444 6750 10446 6802
rect 10498 6750 10500 6802
rect 10444 6738 10500 6750
rect 10556 7476 10612 7486
rect 10220 6690 10276 6702
rect 10220 6638 10222 6690
rect 10274 6638 10276 6690
rect 10220 6580 10276 6638
rect 10220 6514 10276 6524
rect 10556 5906 10612 7420
rect 10668 7474 10724 8540
rect 10780 8372 10836 10558
rect 11004 10610 11060 10622
rect 11004 10558 11006 10610
rect 11058 10558 11060 10610
rect 11004 10388 11060 10558
rect 11004 10322 11060 10332
rect 11228 10610 11284 10780
rect 11228 10558 11230 10610
rect 11282 10558 11284 10610
rect 10892 9716 10948 9726
rect 10892 9714 11060 9716
rect 10892 9662 10894 9714
rect 10946 9662 11060 9714
rect 10892 9660 11060 9662
rect 10892 9650 10948 9660
rect 10780 8306 10836 8316
rect 10892 9042 10948 9054
rect 10892 8990 10894 9042
rect 10946 8990 10948 9042
rect 10780 8148 10836 8158
rect 10892 8148 10948 8990
rect 10780 8146 10948 8148
rect 10780 8094 10782 8146
rect 10834 8094 10948 8146
rect 10780 8092 10948 8094
rect 10780 8082 10836 8092
rect 10668 7422 10670 7474
rect 10722 7422 10724 7474
rect 10668 7410 10724 7422
rect 11004 6804 11060 9660
rect 11228 9714 11284 10558
rect 11452 9828 11508 9838
rect 11452 9734 11508 9772
rect 11564 9826 11620 9838
rect 11564 9774 11566 9826
rect 11618 9774 11620 9826
rect 11228 9662 11230 9714
rect 11282 9662 11284 9714
rect 11228 9650 11284 9662
rect 11564 9044 11620 9774
rect 11676 9156 11732 11676
rect 13020 11620 13076 11630
rect 12908 11170 12964 11182
rect 12908 11118 12910 11170
rect 12962 11118 12964 11170
rect 12348 10610 12404 10622
rect 12348 10558 12350 10610
rect 12402 10558 12404 10610
rect 12348 10388 12404 10558
rect 12348 10322 12404 10332
rect 12012 10276 12068 10286
rect 12012 9938 12068 10220
rect 12908 10276 12964 11118
rect 13020 10722 13076 11564
rect 13020 10670 13022 10722
rect 13074 10670 13076 10722
rect 13020 10658 13076 10670
rect 12908 10210 12964 10220
rect 12012 9886 12014 9938
rect 12066 9886 12068 9938
rect 12012 9874 12068 9886
rect 12236 10164 12292 10174
rect 11676 9100 11956 9156
rect 11564 8978 11620 8988
rect 11900 9042 11956 9100
rect 11900 8990 11902 9042
rect 11954 8990 11956 9042
rect 11340 8818 11396 8830
rect 11340 8766 11342 8818
rect 11394 8766 11396 8818
rect 11228 8708 11284 8718
rect 11116 8034 11172 8046
rect 11116 7982 11118 8034
rect 11170 7982 11172 8034
rect 11116 7700 11172 7982
rect 11116 7634 11172 7644
rect 11116 7476 11172 7486
rect 11228 7476 11284 8652
rect 11340 8260 11396 8766
rect 11676 8818 11732 8830
rect 11676 8766 11678 8818
rect 11730 8766 11732 8818
rect 11676 8708 11732 8766
rect 11340 8194 11396 8204
rect 11564 8652 11676 8708
rect 11116 7474 11284 7476
rect 11116 7422 11118 7474
rect 11170 7422 11284 7474
rect 11116 7420 11284 7422
rect 11452 8146 11508 8158
rect 11452 8094 11454 8146
rect 11506 8094 11508 8146
rect 11452 7476 11508 8094
rect 11116 7410 11172 7420
rect 11452 7410 11508 7420
rect 11004 6738 11060 6748
rect 11564 6690 11620 8652
rect 11676 8642 11732 8652
rect 11900 8484 11956 8990
rect 11564 6638 11566 6690
rect 11618 6638 11620 6690
rect 11564 6626 11620 6638
rect 11676 8428 11900 8484
rect 10780 6580 10836 6590
rect 11116 6580 11172 6590
rect 10836 6524 10948 6580
rect 10780 6514 10836 6524
rect 10556 5854 10558 5906
rect 10610 5854 10612 5906
rect 10556 5842 10612 5854
rect 8876 5124 8932 5134
rect 8876 5030 8932 5068
rect 9324 5122 9380 5628
rect 9324 5070 9326 5122
rect 9378 5070 9380 5122
rect 9324 5058 9380 5070
rect 9884 5628 10164 5684
rect 10220 5794 10276 5806
rect 10220 5742 10222 5794
rect 10274 5742 10276 5794
rect 8540 5012 8596 5022
rect 8540 4564 8596 4956
rect 9884 5010 9940 5628
rect 10108 5460 10164 5470
rect 10108 5122 10164 5404
rect 10220 5348 10276 5742
rect 10668 5572 10724 5582
rect 10724 5516 10836 5572
rect 10668 5506 10724 5516
rect 10220 5282 10276 5292
rect 10556 5460 10612 5470
rect 10108 5070 10110 5122
rect 10162 5070 10164 5122
rect 10108 5058 10164 5070
rect 9884 4958 9886 5010
rect 9938 4958 9940 5010
rect 9884 4946 9940 4958
rect 10556 5010 10612 5404
rect 10556 4958 10558 5010
rect 10610 4958 10612 5010
rect 10556 4946 10612 4958
rect 9528 4732 9792 4742
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9528 4666 9792 4676
rect 8540 4498 8596 4508
rect 8988 4564 9044 4574
rect 8988 4470 9044 4508
rect 10780 4450 10836 5516
rect 10892 5122 10948 6524
rect 11116 6578 11284 6580
rect 11116 6526 11118 6578
rect 11170 6526 11284 6578
rect 11116 6524 11284 6526
rect 11116 6514 11172 6524
rect 11116 6244 11172 6254
rect 10892 5070 10894 5122
rect 10946 5070 10948 5122
rect 10892 5058 10948 5070
rect 11004 6188 11116 6244
rect 11004 5124 11060 6188
rect 11116 6178 11172 6188
rect 11116 6020 11172 6030
rect 11116 5926 11172 5964
rect 11004 4564 11060 5068
rect 11228 5122 11284 6524
rect 11452 6578 11508 6590
rect 11452 6526 11454 6578
rect 11506 6526 11508 6578
rect 11452 6468 11508 6526
rect 11676 6468 11732 8428
rect 11900 8418 11956 8428
rect 12236 9154 12292 10108
rect 12236 9102 12238 9154
rect 12290 9102 12292 9154
rect 12124 8260 12180 8270
rect 12124 8166 12180 8204
rect 11900 8148 11956 8158
rect 11452 6412 11732 6468
rect 11788 8034 11844 8046
rect 11788 7982 11790 8034
rect 11842 7982 11844 8034
rect 11788 6692 11844 7982
rect 11900 7364 11956 8092
rect 11900 7298 11956 7308
rect 12236 7140 12292 9102
rect 12460 9938 12516 9950
rect 12460 9886 12462 9938
rect 12514 9886 12516 9938
rect 12460 8708 12516 9886
rect 12908 9828 12964 9838
rect 12908 9734 12964 9772
rect 12460 8260 12516 8652
rect 13020 9044 13076 9054
rect 12460 8204 12852 8260
rect 12460 8146 12516 8204
rect 12460 8094 12462 8146
rect 12514 8094 12516 8146
rect 12460 8082 12516 8094
rect 12236 7074 12292 7084
rect 12348 8034 12404 8046
rect 12684 8036 12740 8046
rect 12348 7982 12350 8034
rect 12402 7982 12404 8034
rect 12124 6804 12180 6814
rect 11564 6132 11620 6142
rect 11788 6132 11844 6636
rect 11564 6130 11844 6132
rect 11564 6078 11566 6130
rect 11618 6078 11844 6130
rect 11564 6076 11844 6078
rect 11900 6690 11956 6702
rect 11900 6638 11902 6690
rect 11954 6638 11956 6690
rect 11564 6066 11620 6076
rect 11900 6020 11956 6638
rect 12124 6690 12180 6748
rect 12124 6638 12126 6690
rect 12178 6638 12180 6690
rect 12124 6626 12180 6638
rect 12236 6690 12292 6702
rect 12236 6638 12238 6690
rect 12290 6638 12292 6690
rect 11788 5964 11956 6020
rect 11452 5906 11508 5918
rect 11452 5854 11454 5906
rect 11506 5854 11508 5906
rect 11452 5572 11508 5854
rect 11564 5684 11620 5694
rect 11564 5590 11620 5628
rect 11452 5506 11508 5516
rect 11788 5460 11844 5964
rect 11676 5404 11844 5460
rect 11900 5796 11956 5806
rect 12236 5796 12292 6638
rect 12348 6580 12404 7982
rect 12572 8034 12740 8036
rect 12572 7982 12686 8034
rect 12738 7982 12740 8034
rect 12572 7980 12740 7982
rect 12572 6804 12628 7980
rect 12684 7970 12740 7980
rect 12348 6514 12404 6524
rect 12460 6748 12628 6804
rect 12684 7364 12740 7374
rect 11900 5794 12292 5796
rect 11900 5742 11902 5794
rect 11954 5742 12292 5794
rect 11900 5740 12292 5742
rect 12348 6356 12404 6366
rect 11228 5070 11230 5122
rect 11282 5070 11284 5122
rect 11116 4564 11172 4574
rect 11004 4562 11172 4564
rect 11004 4510 11118 4562
rect 11170 4510 11172 4562
rect 11004 4508 11172 4510
rect 11116 4498 11172 4508
rect 11228 4564 11284 5070
rect 11228 4498 11284 4508
rect 11340 5124 11396 5134
rect 10780 4398 10782 4450
rect 10834 4398 10836 4450
rect 10780 4386 10836 4398
rect 8764 4340 8820 4350
rect 8764 4246 8820 4284
rect 10668 4340 10724 4350
rect 8428 3614 8430 3666
rect 8482 3614 8484 3666
rect 8428 3602 8484 3614
rect 10220 4116 10276 4126
rect 10220 3666 10276 4060
rect 10220 3614 10222 3666
rect 10274 3614 10276 3666
rect 10220 3602 10276 3614
rect 9548 3556 9604 3566
rect 9548 3462 9604 3500
rect 10668 3388 10724 4284
rect 11228 4340 11284 4350
rect 11340 4340 11396 5068
rect 11676 5012 11732 5404
rect 11788 5236 11844 5246
rect 11788 5142 11844 5180
rect 11788 5012 11844 5022
rect 11676 4956 11788 5012
rect 11788 4946 11844 4956
rect 11228 4338 11396 4340
rect 11228 4286 11230 4338
rect 11282 4286 11396 4338
rect 11228 4284 11396 4286
rect 11228 4274 11284 4284
rect 11788 4226 11844 4238
rect 11788 4174 11790 4226
rect 11842 4174 11844 4226
rect 10780 3444 10836 3454
rect 11788 3388 11844 4174
rect 10668 3332 10836 3388
rect 8204 3266 8260 3276
rect 9528 3164 9792 3174
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9528 3098 9792 3108
rect 6412 2930 6468 2940
rect 10780 800 10836 3332
rect 11676 3332 11844 3388
rect 11900 3332 11956 5740
rect 12124 5234 12180 5246
rect 12124 5182 12126 5234
rect 12178 5182 12180 5234
rect 12124 5124 12180 5182
rect 12124 5058 12180 5068
rect 12124 4564 12180 4574
rect 12124 4338 12180 4508
rect 12124 4286 12126 4338
rect 12178 4286 12180 4338
rect 12124 4274 12180 4286
rect 12348 3666 12404 6300
rect 12460 6020 12516 6748
rect 12572 6580 12628 6590
rect 12684 6580 12740 7308
rect 12796 7362 12852 8204
rect 12796 7310 12798 7362
rect 12850 7310 12852 7362
rect 12796 7298 12852 7310
rect 12908 8146 12964 8158
rect 12908 8094 12910 8146
rect 12962 8094 12964 8146
rect 12572 6578 12740 6580
rect 12572 6526 12574 6578
rect 12626 6526 12740 6578
rect 12572 6524 12740 6526
rect 12796 7140 12852 7150
rect 12572 6514 12628 6524
rect 12460 5236 12516 5964
rect 12796 6018 12852 7084
rect 12908 6692 12964 8094
rect 13020 7474 13076 8988
rect 13132 7924 13188 12684
rect 13468 12068 13524 15260
rect 14028 15202 14084 15372
rect 14028 15150 14030 15202
rect 14082 15150 14084 15202
rect 14028 15138 14084 15150
rect 14588 15148 14644 19068
rect 14700 18340 14756 18350
rect 14700 18246 14756 18284
rect 14924 16772 14980 20076
rect 15036 20066 15092 20076
rect 15372 20132 15428 20142
rect 15372 20038 15428 20076
rect 15036 19124 15092 19134
rect 15036 19030 15092 19068
rect 15596 18452 15652 22206
rect 15708 21812 15764 21822
rect 15708 20916 15764 21756
rect 16380 21812 16436 21822
rect 16380 21718 16436 21756
rect 16716 21812 16772 21822
rect 16716 21698 16772 21756
rect 16716 21646 16718 21698
rect 16770 21646 16772 21698
rect 15932 21588 15988 21598
rect 15820 20916 15876 20926
rect 15708 20914 15876 20916
rect 15708 20862 15822 20914
rect 15874 20862 15876 20914
rect 15708 20860 15876 20862
rect 15820 20850 15876 20860
rect 15708 20020 15764 20030
rect 15708 19926 15764 19964
rect 15596 18386 15652 18396
rect 15820 17666 15876 17678
rect 15820 17614 15822 17666
rect 15874 17614 15876 17666
rect 15260 17108 15316 17118
rect 15260 16996 15316 17052
rect 15820 17106 15876 17614
rect 15932 17220 15988 21532
rect 16716 20916 16772 21646
rect 17276 21362 17332 25340
rect 17500 25060 17556 25070
rect 17500 24946 17556 25004
rect 17500 24894 17502 24946
rect 17554 24894 17556 24946
rect 17500 24882 17556 24894
rect 17612 23940 17668 26124
rect 17836 25284 17892 26236
rect 18172 26290 18228 26302
rect 18172 26238 18174 26290
rect 18226 26238 18228 26290
rect 18172 25844 18228 26238
rect 18284 26292 18340 26302
rect 18284 26198 18340 26236
rect 18732 26290 18788 26302
rect 18732 26238 18734 26290
rect 18786 26238 18788 26290
rect 18172 25788 18564 25844
rect 18508 25730 18564 25788
rect 18508 25678 18510 25730
rect 18562 25678 18564 25730
rect 18508 25666 18564 25678
rect 18620 25508 18676 25518
rect 18620 25414 18676 25452
rect 17836 25218 17892 25228
rect 18172 25396 18228 25406
rect 17844 25116 18108 25126
rect 17900 25060 17948 25116
rect 18004 25060 18052 25116
rect 17844 25050 18108 25060
rect 18172 24946 18228 25340
rect 18732 25396 18788 26238
rect 18844 26292 18900 26302
rect 18844 26198 18900 26236
rect 18956 25732 19012 25742
rect 19068 25732 19124 27804
rect 19964 27858 20020 27870
rect 19964 27806 19966 27858
rect 20018 27806 20020 27858
rect 18956 25730 19124 25732
rect 18956 25678 18958 25730
rect 19010 25678 19124 25730
rect 18956 25676 19124 25678
rect 19180 26402 19236 26414
rect 19180 26350 19182 26402
rect 19234 26350 19236 26402
rect 18956 25666 19012 25676
rect 18732 25330 18788 25340
rect 18172 24894 18174 24946
rect 18226 24894 18228 24946
rect 18172 24882 18228 24894
rect 18620 25284 18676 25294
rect 19180 25284 19236 26350
rect 19628 26290 19684 26302
rect 19628 26238 19630 26290
rect 19682 26238 19684 26290
rect 19628 26180 19684 26238
rect 19628 26114 19684 26124
rect 19292 25732 19348 25742
rect 19292 25638 19348 25676
rect 19964 25618 20020 27806
rect 20188 27860 20244 27870
rect 20188 27766 20244 27804
rect 20300 26404 20356 28030
rect 20524 27858 20580 27870
rect 20524 27806 20526 27858
rect 20578 27806 20580 27858
rect 20412 27186 20468 27198
rect 20412 27134 20414 27186
rect 20466 27134 20468 27186
rect 20412 26628 20468 27134
rect 20524 26852 20580 27806
rect 22002 27468 22266 27478
rect 22058 27412 22106 27468
rect 22162 27412 22210 27468
rect 22002 27402 22266 27412
rect 30318 27468 30582 27478
rect 30374 27412 30422 27468
rect 30478 27412 30526 27468
rect 30318 27402 30582 27412
rect 23772 27074 23828 27086
rect 23772 27022 23774 27074
rect 23826 27022 23828 27074
rect 20524 26786 20580 26796
rect 23436 26850 23492 26862
rect 23436 26798 23438 26850
rect 23490 26798 23492 26850
rect 20412 26562 20468 26572
rect 22652 26628 22708 26638
rect 20412 26404 20468 26414
rect 20300 26402 20468 26404
rect 20300 26350 20414 26402
rect 20466 26350 20468 26402
rect 20300 26348 20468 26350
rect 20412 26338 20468 26348
rect 22540 26180 22596 26190
rect 22002 25900 22266 25910
rect 22058 25844 22106 25900
rect 22162 25844 22210 25900
rect 22002 25834 22266 25844
rect 19964 25566 19966 25618
rect 20018 25566 20020 25618
rect 19964 25554 20020 25566
rect 20076 25508 20132 25518
rect 20076 25414 20132 25452
rect 22540 25508 22596 26124
rect 19516 25394 19572 25406
rect 19516 25342 19518 25394
rect 19570 25342 19572 25394
rect 19292 25284 19348 25294
rect 19180 25228 19292 25284
rect 18620 25172 18676 25228
rect 19292 25218 19348 25228
rect 18620 25116 18900 25172
rect 17836 24724 17892 24734
rect 18396 24724 18452 24734
rect 17836 24722 18452 24724
rect 17836 24670 17838 24722
rect 17890 24670 18398 24722
rect 18450 24670 18452 24722
rect 17836 24668 18452 24670
rect 17836 24658 17892 24668
rect 17836 23940 17892 23950
rect 17612 23938 17892 23940
rect 17612 23886 17838 23938
rect 17890 23886 17892 23938
rect 17612 23884 17892 23886
rect 17612 23268 17668 23278
rect 17388 22930 17444 22942
rect 17388 22878 17390 22930
rect 17442 22878 17444 22930
rect 17388 22596 17444 22878
rect 17388 22530 17444 22540
rect 17500 22372 17556 22382
rect 17500 22278 17556 22316
rect 17612 21812 17668 23212
rect 17724 23156 17780 23884
rect 17836 23874 17892 23884
rect 17844 23548 18108 23558
rect 17900 23492 17948 23548
rect 18004 23492 18052 23548
rect 17844 23482 18108 23492
rect 17724 23090 17780 23100
rect 18284 23268 18340 23278
rect 18396 23268 18452 24668
rect 18284 23266 18452 23268
rect 18284 23214 18286 23266
rect 18338 23214 18452 23266
rect 18284 23212 18452 23214
rect 18508 23714 18564 23726
rect 18508 23662 18510 23714
rect 18562 23662 18564 23714
rect 17948 23044 18004 23082
rect 17948 22978 18004 22988
rect 17724 22930 17780 22942
rect 17724 22878 17726 22930
rect 17778 22878 17780 22930
rect 17724 22820 17780 22878
rect 18284 22820 18340 23212
rect 17724 22764 18340 22820
rect 17844 21980 18108 21990
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 17844 21914 18108 21924
rect 17948 21812 18004 21822
rect 17612 21810 18004 21812
rect 17612 21758 17950 21810
rect 18002 21758 18004 21810
rect 17612 21756 18004 21758
rect 17948 21746 18004 21756
rect 18284 21700 18340 22764
rect 18060 21644 18228 21700
rect 17276 21310 17278 21362
rect 17330 21310 17332 21362
rect 17276 21298 17332 21310
rect 17612 21588 17668 21598
rect 18060 21588 18116 21644
rect 17612 21586 18116 21588
rect 17612 21534 17614 21586
rect 17666 21534 18116 21586
rect 17612 21532 18116 21534
rect 18172 21586 18228 21644
rect 18284 21634 18340 21644
rect 18396 23044 18452 23054
rect 18508 23044 18564 23662
rect 18620 23380 18676 25116
rect 18732 24948 18788 24958
rect 18732 24164 18788 24892
rect 18844 24946 18900 25116
rect 18844 24894 18846 24946
rect 18898 24894 18900 24946
rect 18844 24882 18900 24894
rect 19068 24724 19124 24734
rect 18956 24722 19124 24724
rect 18956 24670 19070 24722
rect 19122 24670 19124 24722
rect 18956 24668 19124 24670
rect 18844 24164 18900 24174
rect 18732 24162 18900 24164
rect 18732 24110 18846 24162
rect 18898 24110 18900 24162
rect 18732 24108 18900 24110
rect 18844 24098 18900 24108
rect 18620 23314 18676 23324
rect 18844 23828 18900 23838
rect 18844 23378 18900 23772
rect 18844 23326 18846 23378
rect 18898 23326 18900 23378
rect 18844 23314 18900 23326
rect 18956 23380 19012 24668
rect 19068 24658 19124 24668
rect 19516 24612 19572 25342
rect 19852 25396 19908 25406
rect 19852 25302 19908 25340
rect 20300 25284 20356 25294
rect 20300 25190 20356 25228
rect 19516 24546 19572 24556
rect 20300 24722 20356 24734
rect 20300 24670 20302 24722
rect 20354 24670 20356 24722
rect 19180 24052 19236 24062
rect 19852 24052 19908 24062
rect 20300 24052 20356 24670
rect 19180 24050 19796 24052
rect 19180 23998 19182 24050
rect 19234 23998 19796 24050
rect 19180 23996 19796 23998
rect 19180 23986 19236 23996
rect 19516 23828 19572 23838
rect 19516 23734 19572 23772
rect 19740 23826 19796 23996
rect 19852 24050 20132 24052
rect 19852 23998 19854 24050
rect 19906 23998 20132 24050
rect 19852 23996 20132 23998
rect 19852 23986 19908 23996
rect 19740 23774 19742 23826
rect 19794 23774 19796 23826
rect 19740 23762 19796 23774
rect 19068 23716 19124 23726
rect 19068 23714 19236 23716
rect 19068 23662 19070 23714
rect 19122 23662 19236 23714
rect 19068 23660 19236 23662
rect 19068 23650 19124 23660
rect 19180 23604 19236 23660
rect 19180 23548 19796 23604
rect 18956 23314 19012 23324
rect 19628 23380 19684 23390
rect 19068 23268 19124 23278
rect 19068 23174 19124 23212
rect 18620 23156 18676 23166
rect 18620 23154 19012 23156
rect 18620 23102 18622 23154
rect 18674 23102 19012 23154
rect 18620 23100 19012 23102
rect 18620 23090 18676 23100
rect 18452 22988 18564 23044
rect 18172 21534 18174 21586
rect 18226 21534 18228 21586
rect 17612 21140 17668 21532
rect 18172 21522 18228 21534
rect 18396 21476 18452 22988
rect 18956 22484 19012 23100
rect 19180 23154 19236 23166
rect 19516 23156 19572 23166
rect 19180 23102 19182 23154
rect 19234 23102 19236 23154
rect 19180 22708 19236 23102
rect 19404 23154 19572 23156
rect 19404 23102 19518 23154
rect 19570 23102 19572 23154
rect 19404 23100 19572 23102
rect 19292 23044 19348 23054
rect 19404 23044 19460 23100
rect 19516 23090 19572 23100
rect 19348 22988 19460 23044
rect 19292 22978 19348 22988
rect 19628 22932 19684 23324
rect 19180 22652 19572 22708
rect 18956 22428 19348 22484
rect 18956 21812 19012 22428
rect 19292 22370 19348 22428
rect 19292 22318 19294 22370
rect 19346 22318 19348 22370
rect 19292 22306 19348 22318
rect 18956 21746 19012 21756
rect 19404 21812 19460 21822
rect 19404 21718 19460 21756
rect 19292 21700 19348 21710
rect 19292 21606 19348 21644
rect 19516 21588 19572 22652
rect 19628 22260 19684 22876
rect 19628 22166 19684 22204
rect 19628 21812 19684 21822
rect 19740 21812 19796 23548
rect 20076 23380 20132 23996
rect 20300 23958 20356 23996
rect 20524 24610 20580 24622
rect 20524 24558 20526 24610
rect 20578 24558 20580 24610
rect 20076 23324 20356 23380
rect 20300 23266 20356 23324
rect 20300 23214 20302 23266
rect 20354 23214 20356 23266
rect 20300 23202 20356 23214
rect 20412 23268 20468 23278
rect 20300 22596 20356 22606
rect 20412 22596 20468 23212
rect 20300 22594 20468 22596
rect 20300 22542 20302 22594
rect 20354 22542 20468 22594
rect 20300 22540 20468 22542
rect 20300 22530 20356 22540
rect 19684 21756 19796 21812
rect 19852 22372 19908 22382
rect 19852 21812 19908 22316
rect 20076 22372 20132 22382
rect 20076 22278 20132 22316
rect 20412 22370 20468 22382
rect 20412 22318 20414 22370
rect 20466 22318 20468 22370
rect 20188 22260 20244 22270
rect 19964 21812 20020 21822
rect 19852 21810 20132 21812
rect 19852 21758 19966 21810
rect 20018 21758 20132 21810
rect 19852 21756 20132 21758
rect 19628 21746 19684 21756
rect 19964 21746 20020 21756
rect 19628 21588 19684 21598
rect 19516 21586 19684 21588
rect 19516 21534 19630 21586
rect 19682 21534 19684 21586
rect 19516 21532 19684 21534
rect 18284 21420 18452 21476
rect 16716 20850 16772 20860
rect 17276 21084 17668 21140
rect 17724 21362 17780 21374
rect 17724 21310 17726 21362
rect 17778 21310 17780 21362
rect 16044 20804 16100 20814
rect 16044 20710 16100 20748
rect 17164 20692 17220 20702
rect 16380 20578 16436 20590
rect 16380 20526 16382 20578
rect 16434 20526 16436 20578
rect 16156 19908 16212 19918
rect 16044 18340 16100 18350
rect 16044 17778 16100 18284
rect 16156 18228 16212 19852
rect 16380 19908 16436 20526
rect 16604 20132 16660 20142
rect 16604 20018 16660 20076
rect 16604 19966 16606 20018
rect 16658 19966 16660 20018
rect 16604 19954 16660 19966
rect 16828 20130 16884 20142
rect 16828 20078 16830 20130
rect 16882 20078 16884 20130
rect 16380 19842 16436 19852
rect 16828 19684 16884 20078
rect 16884 19628 17108 19684
rect 16828 19618 16884 19628
rect 16940 19012 16996 19022
rect 16828 18564 16884 18574
rect 16492 18340 16548 18350
rect 16156 18172 16324 18228
rect 16044 17726 16046 17778
rect 16098 17726 16100 17778
rect 16044 17714 16100 17726
rect 16156 17666 16212 17678
rect 16156 17614 16158 17666
rect 16210 17614 16212 17666
rect 16156 17556 16212 17614
rect 16156 17490 16212 17500
rect 15932 17164 16100 17220
rect 15820 17054 15822 17106
rect 15874 17054 15876 17106
rect 15820 17042 15876 17054
rect 14924 16706 14980 16716
rect 15036 16940 15316 16996
rect 15932 16996 15988 17006
rect 14924 16100 14980 16110
rect 14812 15988 14868 15998
rect 14812 15894 14868 15932
rect 14924 15538 14980 16044
rect 15036 15986 15092 16940
rect 15932 16902 15988 16940
rect 15372 16882 15428 16894
rect 15372 16830 15374 16882
rect 15426 16830 15428 16882
rect 15260 16660 15316 16670
rect 15260 16566 15316 16604
rect 15036 15934 15038 15986
rect 15090 15934 15092 15986
rect 15036 15922 15092 15934
rect 15148 16098 15204 16110
rect 15148 16046 15150 16098
rect 15202 16046 15204 16098
rect 15148 15988 15204 16046
rect 15260 15988 15316 15998
rect 15148 15932 15260 15988
rect 15260 15922 15316 15932
rect 14924 15486 14926 15538
rect 14978 15486 14980 15538
rect 14924 15474 14980 15486
rect 15148 15764 15204 15774
rect 14812 15316 14868 15326
rect 14812 15222 14868 15260
rect 14252 15092 14644 15148
rect 15148 15148 15204 15708
rect 15260 15428 15316 15438
rect 15260 15314 15316 15372
rect 15260 15262 15262 15314
rect 15314 15262 15316 15314
rect 15260 15250 15316 15262
rect 15372 15202 15428 16830
rect 15708 16882 15764 16894
rect 15708 16830 15710 16882
rect 15762 16830 15764 16882
rect 15596 16772 15652 16782
rect 15484 16100 15540 16110
rect 15484 16006 15540 16044
rect 15484 15540 15540 15550
rect 15596 15540 15652 16716
rect 15708 16436 15764 16830
rect 16044 16772 16100 17164
rect 15932 16716 16100 16772
rect 15708 16380 15876 16436
rect 15708 16098 15764 16110
rect 15708 16046 15710 16098
rect 15762 16046 15764 16098
rect 15708 15764 15764 16046
rect 15708 15698 15764 15708
rect 15540 15484 15652 15540
rect 15708 15540 15764 15550
rect 15820 15540 15876 16380
rect 15932 16324 15988 16716
rect 16268 16660 16324 18172
rect 16492 17666 16548 18284
rect 16492 17614 16494 17666
rect 16546 17614 16548 17666
rect 16492 17602 16548 17614
rect 16828 18338 16884 18508
rect 16828 18286 16830 18338
rect 16882 18286 16884 18338
rect 16716 16996 16772 17006
rect 16716 16902 16772 16940
rect 16380 16884 16436 16894
rect 16380 16882 16660 16884
rect 16380 16830 16382 16882
rect 16434 16830 16660 16882
rect 16380 16828 16660 16830
rect 16380 16818 16436 16828
rect 16268 16604 16548 16660
rect 15932 16268 16324 16324
rect 15932 16098 15988 16268
rect 15932 16046 15934 16098
rect 15986 16046 15988 16098
rect 15932 16034 15988 16046
rect 16156 16100 16212 16110
rect 16044 15988 16100 16026
rect 16156 16006 16212 16044
rect 16044 15922 16100 15932
rect 15708 15538 15876 15540
rect 15708 15486 15710 15538
rect 15762 15486 15876 15538
rect 15708 15484 15876 15486
rect 15484 15446 15540 15484
rect 15372 15150 15374 15202
rect 15426 15150 15428 15202
rect 15148 15092 15316 15148
rect 15372 15138 15428 15150
rect 15708 15316 15764 15484
rect 16268 15426 16324 16268
rect 16268 15374 16270 15426
rect 16322 15374 16324 15426
rect 16268 15362 16324 15374
rect 13686 14924 13950 14934
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13686 14858 13950 14868
rect 13580 14420 13636 14430
rect 13580 14326 13636 14364
rect 14140 13972 14196 13982
rect 14140 13878 14196 13916
rect 13686 13356 13950 13366
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13686 13290 13950 13300
rect 14140 12852 14196 12862
rect 14252 12852 14308 15092
rect 14140 12850 14308 12852
rect 14140 12798 14142 12850
rect 14194 12798 14308 12850
rect 14140 12796 14308 12798
rect 15260 13746 15316 15092
rect 15260 13694 15262 13746
rect 15314 13694 15316 13746
rect 14140 12786 14196 12796
rect 13804 12740 13860 12750
rect 13804 12646 13860 12684
rect 14588 12738 14644 12750
rect 14588 12686 14590 12738
rect 14642 12686 14644 12738
rect 13580 12068 13636 12078
rect 13468 12066 13636 12068
rect 13468 12014 13582 12066
rect 13634 12014 13636 12066
rect 13468 12012 13636 12014
rect 13468 11394 13524 12012
rect 13580 12002 13636 12012
rect 13686 11788 13950 11798
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13686 11722 13950 11732
rect 14252 11508 14308 11518
rect 14252 11414 14308 11452
rect 13468 11342 13470 11394
rect 13522 11342 13524 11394
rect 13468 10388 13524 11342
rect 13468 10322 13524 10332
rect 13686 10220 13950 10230
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13686 10154 13950 10164
rect 13692 10052 13748 10062
rect 13692 9826 13748 9996
rect 13692 9774 13694 9826
rect 13746 9774 13748 9826
rect 13692 9762 13748 9774
rect 14140 9714 14196 9726
rect 14140 9662 14142 9714
rect 14194 9662 14196 9714
rect 13580 9604 13636 9614
rect 13468 9548 13580 9604
rect 13244 9042 13300 9054
rect 13244 8990 13246 9042
rect 13298 8990 13300 9042
rect 13244 7924 13300 8990
rect 13468 8596 13524 9548
rect 13580 9510 13636 9548
rect 14140 9604 14196 9662
rect 14140 9538 14196 9548
rect 13804 9044 13860 9054
rect 13804 8950 13860 8988
rect 14140 9044 14196 9054
rect 13686 8652 13950 8662
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13686 8586 13950 8596
rect 13468 8530 13524 8540
rect 13356 8484 13412 8494
rect 13356 8370 13412 8428
rect 13356 8318 13358 8370
rect 13410 8318 13412 8370
rect 13356 8306 13412 8318
rect 13804 8484 13860 8494
rect 13468 8260 13524 8270
rect 13468 8166 13524 8204
rect 13468 7924 13524 7934
rect 13244 7868 13468 7924
rect 13132 7858 13188 7868
rect 13020 7422 13022 7474
rect 13074 7422 13076 7474
rect 13020 7410 13076 7422
rect 13132 6692 13188 6702
rect 12908 6636 13132 6692
rect 12796 5966 12798 6018
rect 12850 5966 12852 6018
rect 12796 5908 12852 5966
rect 12796 5842 12852 5852
rect 13132 5906 13188 6636
rect 13468 6580 13524 7868
rect 13804 7474 13860 8428
rect 13804 7422 13806 7474
rect 13858 7422 13860 7474
rect 13804 7410 13860 7422
rect 13686 7084 13950 7094
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13686 7018 13950 7028
rect 14028 6802 14084 6814
rect 14028 6750 14030 6802
rect 14082 6750 14084 6802
rect 13804 6580 13860 6590
rect 13468 6578 13860 6580
rect 13468 6526 13806 6578
rect 13858 6526 13860 6578
rect 13468 6524 13860 6526
rect 13804 6356 13860 6524
rect 13804 6290 13860 6300
rect 13580 6132 13636 6142
rect 13580 6038 13636 6076
rect 13692 6020 13748 6030
rect 13692 5926 13748 5964
rect 13132 5854 13134 5906
rect 13186 5854 13188 5906
rect 12460 5010 12516 5180
rect 12684 5124 12740 5134
rect 12684 5030 12740 5068
rect 13132 5124 13188 5854
rect 13686 5516 13950 5526
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13686 5450 13950 5460
rect 13692 5348 13748 5358
rect 13132 5058 13188 5068
rect 13468 5122 13524 5134
rect 13468 5070 13470 5122
rect 13522 5070 13524 5122
rect 12460 4958 12462 5010
rect 12514 4958 12516 5010
rect 12460 4946 12516 4958
rect 13356 5012 13412 5022
rect 13356 4450 13412 4956
rect 13468 4564 13524 5070
rect 13580 4900 13636 4910
rect 13580 4806 13636 4844
rect 13468 4498 13524 4508
rect 13356 4398 13358 4450
rect 13410 4398 13412 4450
rect 13356 4386 13412 4398
rect 12348 3614 12350 3666
rect 12402 3614 12404 3666
rect 12348 3602 12404 3614
rect 12572 4340 12628 4350
rect 12572 3556 12628 4284
rect 13692 4116 13748 5292
rect 13916 5124 13972 5134
rect 13916 5030 13972 5068
rect 14028 5012 14084 6750
rect 14140 6690 14196 8988
rect 14588 9044 14644 12686
rect 15148 10500 15204 10510
rect 15260 10500 15316 13694
rect 15708 14420 15764 15260
rect 15932 15316 15988 15326
rect 15932 15314 16100 15316
rect 15932 15262 15934 15314
rect 15986 15262 16100 15314
rect 15932 15260 16100 15262
rect 15932 15250 15988 15260
rect 15820 14420 15876 14430
rect 15708 14418 15876 14420
rect 15708 14366 15822 14418
rect 15874 14366 15876 14418
rect 15708 14364 15876 14366
rect 15708 12852 15764 14364
rect 15820 14354 15876 14364
rect 15932 14306 15988 14318
rect 15932 14254 15934 14306
rect 15986 14254 15988 14306
rect 15932 14084 15988 14254
rect 15820 14028 15988 14084
rect 15820 13746 15876 14028
rect 15932 13860 15988 13870
rect 16044 13860 16100 15260
rect 16380 15092 16436 15102
rect 16380 14998 16436 15036
rect 16492 14980 16548 16604
rect 16492 14914 16548 14924
rect 16604 16098 16660 16828
rect 16828 16882 16884 18286
rect 16940 17556 16996 18956
rect 17052 17780 17108 19628
rect 17052 17686 17108 17724
rect 16940 17500 17108 17556
rect 16828 16830 16830 16882
rect 16882 16830 16884 16882
rect 16716 16660 16772 16670
rect 16716 16566 16772 16604
rect 16828 16324 16884 16830
rect 16940 16324 16996 16334
rect 16828 16268 16940 16324
rect 16940 16258 16996 16268
rect 16604 16046 16606 16098
rect 16658 16046 16660 16098
rect 16604 14644 16660 16046
rect 16716 16100 16772 16110
rect 16716 15426 16772 16044
rect 16940 15988 16996 15998
rect 16940 15894 16996 15932
rect 16828 15874 16884 15886
rect 16828 15822 16830 15874
rect 16882 15822 16884 15874
rect 16828 15764 16884 15822
rect 16828 15698 16884 15708
rect 16716 15374 16718 15426
rect 16770 15374 16772 15426
rect 16716 15362 16772 15374
rect 16828 15428 16884 15438
rect 16828 15334 16884 15372
rect 16940 15092 16996 15102
rect 16156 14588 16660 14644
rect 16716 14980 16772 14990
rect 16156 14530 16212 14588
rect 16156 14478 16158 14530
rect 16210 14478 16212 14530
rect 16156 14466 16212 14478
rect 16492 14420 16548 14430
rect 16716 14420 16772 14924
rect 16940 14532 16996 15036
rect 16940 14438 16996 14476
rect 16492 14418 16772 14420
rect 16492 14366 16494 14418
rect 16546 14366 16772 14418
rect 16492 14364 16772 14366
rect 15932 13858 16100 13860
rect 15932 13806 15934 13858
rect 15986 13806 16100 13858
rect 15932 13804 16100 13806
rect 16268 13972 16324 13982
rect 15932 13794 15988 13804
rect 15820 13694 15822 13746
rect 15874 13694 15876 13746
rect 15820 13412 15876 13694
rect 15820 13356 15988 13412
rect 15708 12786 15764 12796
rect 15820 13188 15876 13198
rect 15148 10498 15316 10500
rect 15148 10446 15150 10498
rect 15202 10446 15316 10498
rect 15148 10444 15316 10446
rect 15148 10434 15204 10444
rect 14588 8978 14644 8988
rect 14700 10388 14756 10398
rect 14700 8932 14756 10332
rect 14924 10052 14980 10062
rect 14980 9996 15092 10052
rect 14924 9986 14980 9996
rect 14812 9156 14868 9166
rect 14812 9154 14980 9156
rect 14812 9102 14814 9154
rect 14866 9102 14980 9154
rect 14812 9100 14980 9102
rect 14812 9090 14868 9100
rect 14924 9044 14980 9100
rect 14700 8876 14868 8932
rect 14700 8260 14756 8270
rect 14476 7364 14532 7374
rect 14476 7270 14532 7308
rect 14140 6638 14142 6690
rect 14194 6638 14196 6690
rect 14140 6244 14196 6638
rect 14140 6178 14196 6188
rect 14700 6690 14756 8204
rect 14700 6638 14702 6690
rect 14754 6638 14756 6690
rect 14252 6018 14308 6030
rect 14252 5966 14254 6018
rect 14306 5966 14308 6018
rect 14252 5908 14308 5966
rect 14700 6020 14756 6638
rect 14812 6692 14868 8876
rect 14924 8596 14980 8988
rect 14924 8530 14980 8540
rect 15036 8428 15092 9996
rect 15820 9938 15876 13132
rect 15932 11508 15988 13356
rect 16044 12964 16100 12974
rect 16044 12870 16100 12908
rect 16268 12740 16324 13916
rect 16492 13524 16548 14364
rect 17052 14084 17108 17500
rect 17164 15148 17220 20636
rect 17276 20020 17332 21084
rect 17388 20916 17444 20926
rect 17388 20692 17444 20860
rect 17612 20802 17668 20814
rect 17612 20750 17614 20802
rect 17666 20750 17668 20802
rect 17612 20692 17668 20750
rect 17388 20690 17556 20692
rect 17388 20638 17390 20690
rect 17442 20638 17556 20690
rect 17388 20636 17556 20638
rect 17388 20626 17444 20636
rect 17276 19124 17332 19964
rect 17500 19460 17556 20636
rect 17612 20626 17668 20636
rect 17724 20580 17780 21310
rect 17724 20018 17780 20524
rect 18172 20802 18228 20814
rect 18172 20750 18174 20802
rect 18226 20750 18228 20802
rect 17844 20412 18108 20422
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 17844 20346 18108 20356
rect 18172 20188 18228 20750
rect 18284 20356 18340 21420
rect 18396 20580 18452 20590
rect 18396 20486 18452 20524
rect 18284 20300 18452 20356
rect 17948 20132 18228 20188
rect 17948 20066 18004 20076
rect 17724 19966 17726 20018
rect 17778 19966 17780 20018
rect 17724 19954 17780 19966
rect 18060 20018 18116 20030
rect 18060 19966 18062 20018
rect 18114 19966 18116 20018
rect 18060 19796 18116 19966
rect 18172 20020 18228 20030
rect 18172 19926 18228 19964
rect 18284 20018 18340 20030
rect 18284 19966 18286 20018
rect 18338 19966 18340 20018
rect 18284 19908 18340 19966
rect 18284 19842 18340 19852
rect 18060 19730 18116 19740
rect 18396 19684 18452 20300
rect 18620 20020 18676 20030
rect 18620 19926 18676 19964
rect 18956 20018 19012 20030
rect 18956 19966 18958 20018
rect 19010 19966 19012 20018
rect 18284 19628 18452 19684
rect 18956 19796 19012 19966
rect 19180 20018 19236 20030
rect 19180 19966 19182 20018
rect 19234 19966 19236 20018
rect 17612 19460 17668 19470
rect 17500 19458 17668 19460
rect 17500 19406 17614 19458
rect 17666 19406 17668 19458
rect 17500 19404 17668 19406
rect 17612 19394 17668 19404
rect 17276 19058 17332 19068
rect 17388 19348 17444 19358
rect 17388 19012 17444 19292
rect 18284 19124 18340 19628
rect 18396 19348 18452 19358
rect 18396 19254 18452 19292
rect 18284 19068 18452 19124
rect 17948 19012 18004 19022
rect 17388 18946 17444 18956
rect 17724 19010 18004 19012
rect 17724 18958 17950 19010
rect 18002 18958 18004 19010
rect 17724 18956 18004 18958
rect 17500 18564 17556 18574
rect 17556 18508 17668 18564
rect 17500 18498 17556 18508
rect 17388 18450 17444 18462
rect 17388 18398 17390 18450
rect 17442 18398 17444 18450
rect 17388 17780 17444 18398
rect 17612 18450 17668 18508
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17612 18386 17668 18398
rect 17500 18340 17556 18350
rect 17500 18246 17556 18284
rect 17276 17724 17556 17780
rect 17276 17108 17332 17724
rect 17276 16098 17332 17052
rect 17388 17556 17444 17566
rect 17388 17106 17444 17500
rect 17500 17554 17556 17724
rect 17500 17502 17502 17554
rect 17554 17502 17556 17554
rect 17500 17490 17556 17502
rect 17724 17444 17780 18956
rect 17948 18946 18004 18956
rect 17844 18844 18108 18854
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 17844 18778 18108 18788
rect 17948 18450 18004 18462
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17948 18228 18004 18398
rect 17948 18162 18004 18172
rect 18172 17556 18228 17566
rect 17836 17444 17892 17482
rect 18172 17462 18228 17500
rect 17724 17388 17836 17444
rect 17836 17378 17892 17388
rect 17844 17276 18108 17286
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 17388 17054 17390 17106
rect 17442 17054 17444 17106
rect 17388 17042 17444 17054
rect 17500 17164 17780 17220
rect 17844 17210 18108 17220
rect 17500 16548 17556 17164
rect 17388 16492 17556 16548
rect 17612 16994 17668 17006
rect 17612 16942 17614 16994
rect 17666 16942 17668 16994
rect 17612 16772 17668 16942
rect 17724 16994 17780 17164
rect 18172 17108 18228 17118
rect 17724 16942 17726 16994
rect 17778 16942 17780 16994
rect 17724 16930 17780 16942
rect 17836 16996 17892 17006
rect 17388 16210 17444 16492
rect 17388 16158 17390 16210
rect 17442 16158 17444 16210
rect 17388 16146 17444 16158
rect 17276 16046 17278 16098
rect 17330 16046 17332 16098
rect 17276 16034 17332 16046
rect 17612 16100 17668 16716
rect 17612 16034 17668 16044
rect 17724 16100 17780 16110
rect 17836 16100 17892 16940
rect 17948 16994 18004 17006
rect 17948 16942 17950 16994
rect 18002 16942 18004 16994
rect 17948 16884 18004 16942
rect 17948 16818 18004 16828
rect 18172 16770 18228 17052
rect 18172 16718 18174 16770
rect 18226 16718 18228 16770
rect 18172 16706 18228 16718
rect 17948 16324 18004 16334
rect 17948 16230 18004 16268
rect 17724 16098 17892 16100
rect 17724 16046 17726 16098
rect 17778 16046 17892 16098
rect 17724 16044 17892 16046
rect 17724 16034 17780 16044
rect 18284 15876 18340 15886
rect 17844 15708 18108 15718
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 17844 15642 18108 15652
rect 17948 15316 18004 15326
rect 18172 15316 18228 15326
rect 17948 15314 18228 15316
rect 17948 15262 17950 15314
rect 18002 15262 18174 15314
rect 18226 15262 18228 15314
rect 17948 15260 18228 15262
rect 17948 15204 18004 15260
rect 18172 15250 18228 15260
rect 17164 15092 17556 15148
rect 17948 15138 18004 15148
rect 18284 15148 18340 15820
rect 18396 15540 18452 19068
rect 18956 18676 19012 19740
rect 19068 19906 19124 19918
rect 19068 19854 19070 19906
rect 19122 19854 19124 19906
rect 19068 19124 19124 19854
rect 19180 19908 19236 19966
rect 19628 20020 19684 21532
rect 19628 19954 19684 19964
rect 19180 19842 19236 19852
rect 19068 19068 19572 19124
rect 18956 18610 19012 18620
rect 19516 18562 19572 19068
rect 19516 18510 19518 18562
rect 19570 18510 19572 18562
rect 19516 18498 19572 18510
rect 18508 18452 18564 18462
rect 18732 18452 18788 18462
rect 18564 18450 18788 18452
rect 18564 18398 18734 18450
rect 18786 18398 18788 18450
rect 18564 18396 18788 18398
rect 18508 18386 18564 18396
rect 18732 18386 18788 18396
rect 18956 17554 19012 17566
rect 18956 17502 18958 17554
rect 19010 17502 19012 17554
rect 18508 17444 18564 17454
rect 18508 17220 18564 17388
rect 18508 17154 18564 17164
rect 18956 17108 19012 17502
rect 19068 17444 19124 17454
rect 19068 17350 19124 17388
rect 18956 17042 19012 17052
rect 19628 17220 19684 17230
rect 18508 16772 18564 16782
rect 18508 16678 18564 16716
rect 19292 16660 19348 16670
rect 19292 16098 19348 16604
rect 19292 16046 19294 16098
rect 19346 16046 19348 16098
rect 19292 16034 19348 16046
rect 18732 15988 18788 15998
rect 18732 15894 18788 15932
rect 18844 15876 18900 15886
rect 19068 15876 19124 15886
rect 18844 15874 19012 15876
rect 18844 15822 18846 15874
rect 18898 15822 19012 15874
rect 18844 15820 19012 15822
rect 18844 15810 18900 15820
rect 18956 15540 19012 15820
rect 19068 15782 19124 15820
rect 18396 15484 18900 15540
rect 18732 15316 18788 15326
rect 18284 15092 18676 15148
rect 17276 14532 17332 14542
rect 17276 14438 17332 14476
rect 16828 14028 17108 14084
rect 17388 14308 17444 14318
rect 16828 13970 16884 14028
rect 16828 13918 16830 13970
rect 16882 13918 16884 13970
rect 16604 13524 16660 13534
rect 16492 13468 16604 13524
rect 16604 13458 16660 13468
rect 16268 12646 16324 12684
rect 16604 12962 16660 12974
rect 16604 12910 16606 12962
rect 16658 12910 16660 12962
rect 16380 11508 16436 11518
rect 15932 11506 16436 11508
rect 15932 11454 16382 11506
rect 16434 11454 16436 11506
rect 15932 11452 16436 11454
rect 16380 11442 16436 11452
rect 15820 9886 15822 9938
rect 15874 9886 15876 9938
rect 15820 9874 15876 9886
rect 15708 9826 15764 9838
rect 15708 9774 15710 9826
rect 15762 9774 15764 9826
rect 15708 9268 15764 9774
rect 15708 9212 15876 9268
rect 14924 8372 15092 8428
rect 15708 9042 15764 9054
rect 15708 8990 15710 9042
rect 15762 8990 15764 9042
rect 15708 8484 15764 8990
rect 15820 8932 15876 9212
rect 16044 8932 16100 8942
rect 15820 8930 16100 8932
rect 15820 8878 16046 8930
rect 16098 8878 16100 8930
rect 15820 8876 16100 8878
rect 16044 8820 16100 8876
rect 16044 8754 16100 8764
rect 16156 8930 16212 8942
rect 16156 8878 16158 8930
rect 16210 8878 16212 8930
rect 14924 8146 14980 8372
rect 15372 8258 15428 8270
rect 15372 8206 15374 8258
rect 15426 8206 15428 8258
rect 14924 8094 14926 8146
rect 14978 8094 14980 8146
rect 14924 8082 14980 8094
rect 15036 8148 15092 8158
rect 15036 7474 15092 8092
rect 15372 7924 15428 8206
rect 15372 7858 15428 7868
rect 15036 7422 15038 7474
rect 15090 7422 15092 7474
rect 15036 7410 15092 7422
rect 15260 6692 15316 6702
rect 14812 6690 15316 6692
rect 14812 6638 15262 6690
rect 15314 6638 15316 6690
rect 14812 6636 15316 6638
rect 14700 5954 14756 5964
rect 14812 6244 14868 6254
rect 14252 5842 14308 5852
rect 14588 5908 14644 5918
rect 14588 5814 14644 5852
rect 14812 5908 14868 6188
rect 14812 5842 14868 5852
rect 14028 5010 14196 5012
rect 14028 4958 14030 5010
rect 14082 4958 14196 5010
rect 14028 4956 14196 4958
rect 14028 4946 14084 4956
rect 13468 4060 13748 4116
rect 13468 3668 13524 4060
rect 13686 3948 13950 3958
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13686 3882 13950 3892
rect 14140 3780 14196 4956
rect 14140 3686 14196 3724
rect 14476 4900 14532 4910
rect 14476 3778 14532 4844
rect 14476 3726 14478 3778
rect 14530 3726 14532 3778
rect 14476 3714 14532 3726
rect 14924 4452 14980 4462
rect 14924 3778 14980 4396
rect 15036 4340 15092 6636
rect 15260 6626 15316 6636
rect 15484 6132 15540 6142
rect 15036 4274 15092 4284
rect 15372 4898 15428 4910
rect 15372 4846 15374 4898
rect 15426 4846 15428 4898
rect 14924 3726 14926 3778
rect 14978 3726 14980 3778
rect 14924 3714 14980 3726
rect 15260 3780 15316 3790
rect 15260 3686 15316 3724
rect 13580 3668 13636 3678
rect 13468 3666 13636 3668
rect 13468 3614 13582 3666
rect 13634 3614 13636 3666
rect 13468 3612 13636 3614
rect 13580 3602 13636 3612
rect 15372 3668 15428 4846
rect 15484 4226 15540 6076
rect 15708 5906 15764 8428
rect 16156 8372 16212 8878
rect 16604 8932 16660 12910
rect 16828 12964 16884 13918
rect 17388 13858 17444 14252
rect 17388 13806 17390 13858
rect 17442 13806 17444 13858
rect 17388 13794 17444 13806
rect 16828 12898 16884 12908
rect 16940 12964 16996 12974
rect 16940 12962 17108 12964
rect 16940 12910 16942 12962
rect 16994 12910 17108 12962
rect 16940 12908 17108 12910
rect 16940 12898 16996 12908
rect 16940 12740 16996 12750
rect 16604 8866 16660 8876
rect 16716 11282 16772 11294
rect 16716 11230 16718 11282
rect 16770 11230 16772 11282
rect 15708 5854 15710 5906
rect 15762 5854 15764 5906
rect 15708 5842 15764 5854
rect 15932 8316 16212 8372
rect 15932 5124 15988 8316
rect 16156 8146 16212 8158
rect 16156 8094 16158 8146
rect 16210 8094 16212 8146
rect 16044 6578 16100 6590
rect 16044 6526 16046 6578
rect 16098 6526 16100 6578
rect 16044 6244 16100 6526
rect 16044 6178 16100 6188
rect 16156 5908 16212 8094
rect 16716 7924 16772 11230
rect 16828 11170 16884 11182
rect 16828 11118 16830 11170
rect 16882 11118 16884 11170
rect 16828 9828 16884 11118
rect 16940 10836 16996 12684
rect 17052 11732 17108 12908
rect 17388 12852 17444 12862
rect 17388 12758 17444 12796
rect 17500 12404 17556 15092
rect 18620 14754 18676 15092
rect 18620 14702 18622 14754
rect 18674 14702 18676 14754
rect 18620 14690 18676 14702
rect 18732 14642 18788 15260
rect 18732 14590 18734 14642
rect 18786 14590 18788 14642
rect 18732 14578 18788 14590
rect 17724 14420 17780 14430
rect 17612 14418 18228 14420
rect 17612 14366 17726 14418
rect 17778 14366 18228 14418
rect 17612 14364 18228 14366
rect 17612 12964 17668 14364
rect 17724 14354 17780 14364
rect 17844 14140 18108 14150
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 17844 14074 18108 14084
rect 17724 13860 17780 13870
rect 17724 13766 17780 13804
rect 18172 13746 18228 14364
rect 18844 14308 18900 15484
rect 18956 15474 19012 15484
rect 19068 15428 19124 15438
rect 19068 14418 19124 15372
rect 19068 14366 19070 14418
rect 19122 14366 19124 14418
rect 19068 14354 19124 14366
rect 19180 14420 19236 14430
rect 18396 13972 18452 13982
rect 18396 13878 18452 13916
rect 18844 13972 18900 14252
rect 18844 13970 19124 13972
rect 18844 13918 18846 13970
rect 18898 13918 19124 13970
rect 18844 13916 19124 13918
rect 18844 13906 18900 13916
rect 18172 13694 18174 13746
rect 18226 13694 18228 13746
rect 18172 13682 18228 13694
rect 18732 13748 18788 13758
rect 17612 12962 17780 12964
rect 17612 12910 17614 12962
rect 17666 12910 17780 12962
rect 17612 12908 17780 12910
rect 17612 12898 17668 12908
rect 17388 12348 17556 12404
rect 17052 11676 17332 11732
rect 17276 11620 17332 11676
rect 17276 11526 17332 11564
rect 17388 11060 17444 12348
rect 17612 12292 17668 12302
rect 17500 12178 17556 12190
rect 17500 12126 17502 12178
rect 17554 12126 17556 12178
rect 17500 11284 17556 12126
rect 17612 11618 17668 12236
rect 17612 11566 17614 11618
rect 17666 11566 17668 11618
rect 17612 11554 17668 11566
rect 17724 11396 17780 12908
rect 18284 12962 18340 12974
rect 18284 12910 18286 12962
rect 18338 12910 18340 12962
rect 18172 12740 18228 12750
rect 17844 12572 18108 12582
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 17844 12506 18108 12516
rect 18172 12290 18228 12684
rect 18172 12238 18174 12290
rect 18226 12238 18228 12290
rect 18172 12226 18228 12238
rect 18284 12292 18340 12910
rect 18284 12226 18340 12236
rect 18396 12964 18452 12974
rect 18396 11844 18452 12908
rect 18620 12850 18676 12862
rect 18620 12798 18622 12850
rect 18674 12798 18676 12850
rect 18508 12738 18564 12750
rect 18508 12686 18510 12738
rect 18562 12686 18564 12738
rect 18508 12404 18564 12686
rect 18620 12740 18676 12798
rect 18732 12740 18788 13692
rect 18956 13524 19012 13534
rect 18956 12962 19012 13468
rect 18956 12910 18958 12962
rect 19010 12910 19012 12962
rect 18620 12684 18900 12740
rect 18508 12338 18564 12348
rect 18396 11788 18676 11844
rect 18172 11620 18228 11630
rect 17836 11396 17892 11406
rect 17724 11394 17892 11396
rect 17724 11342 17838 11394
rect 17890 11342 17892 11394
rect 17724 11340 17892 11342
rect 17836 11330 17892 11340
rect 17500 11218 17556 11228
rect 17388 11004 17780 11060
rect 17388 10836 17444 10846
rect 16940 10834 17444 10836
rect 16940 10782 16942 10834
rect 16994 10782 17390 10834
rect 17442 10782 17444 10834
rect 16940 10780 17444 10782
rect 16940 10770 16996 10780
rect 17388 10770 17444 10780
rect 17724 10500 17780 11004
rect 17844 11004 18108 11014
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 17844 10938 18108 10948
rect 17836 10500 17892 10510
rect 16828 9762 16884 9772
rect 17612 10498 17892 10500
rect 17612 10446 17838 10498
rect 17890 10446 17892 10498
rect 17612 10444 17892 10446
rect 17612 9716 17668 10444
rect 17836 10434 17892 10444
rect 17836 9828 17892 9838
rect 17836 9734 17892 9772
rect 18172 9826 18228 11564
rect 18508 11284 18564 11294
rect 18508 10610 18564 11228
rect 18508 10558 18510 10610
rect 18562 10558 18564 10610
rect 18508 10164 18564 10558
rect 18508 10098 18564 10108
rect 18172 9774 18174 9826
rect 18226 9774 18228 9826
rect 17612 9042 17668 9660
rect 17612 8990 17614 9042
rect 17666 8990 17668 9042
rect 17612 8978 17668 8990
rect 17724 9714 17780 9726
rect 17724 9662 17726 9714
rect 17778 9662 17780 9714
rect 17724 9044 17780 9662
rect 17844 9436 18108 9446
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 17844 9370 18108 9380
rect 18172 9154 18228 9774
rect 18620 9828 18676 11788
rect 18732 11618 18788 11630
rect 18732 11566 18734 11618
rect 18786 11566 18788 11618
rect 18732 11506 18788 11566
rect 18732 11454 18734 11506
rect 18786 11454 18788 11506
rect 18732 11442 18788 11454
rect 18620 9714 18676 9772
rect 18620 9662 18622 9714
rect 18674 9662 18676 9714
rect 18620 9650 18676 9662
rect 18732 11284 18788 11294
rect 18844 11284 18900 12684
rect 18956 11618 19012 12910
rect 19068 11732 19124 13916
rect 19068 11666 19124 11676
rect 18956 11566 18958 11618
rect 19010 11566 19012 11618
rect 18956 11554 19012 11566
rect 19068 11508 19124 11518
rect 19180 11508 19236 14364
rect 19516 14418 19572 14430
rect 19516 14366 19518 14418
rect 19570 14366 19572 14418
rect 19516 13972 19572 14366
rect 19628 14418 19684 17164
rect 20076 16772 20132 21756
rect 20188 21586 20244 22204
rect 20188 21534 20190 21586
rect 20242 21534 20244 21586
rect 20188 21522 20244 21534
rect 20412 21028 20468 22318
rect 20524 21924 20580 24558
rect 22428 24612 22484 24622
rect 22002 24332 22266 24342
rect 22058 24276 22106 24332
rect 22162 24276 22210 24332
rect 22002 24266 22266 24276
rect 22428 24050 22484 24556
rect 22428 23998 22430 24050
rect 22482 23998 22484 24050
rect 22428 23986 22484 23998
rect 22204 23938 22260 23950
rect 22204 23886 22206 23938
rect 22258 23886 22260 23938
rect 22204 23828 22260 23886
rect 22540 23828 22596 25452
rect 22652 24722 22708 26572
rect 23436 25732 23492 26798
rect 22988 25618 23044 25630
rect 22988 25566 22990 25618
rect 23042 25566 23044 25618
rect 22988 24948 23044 25566
rect 22988 24882 23044 24892
rect 23212 25284 23268 25294
rect 22652 24670 22654 24722
rect 22706 24670 22708 24722
rect 22652 24658 22708 24670
rect 22204 23772 22596 23828
rect 22764 23940 22820 23950
rect 20972 23268 21028 23278
rect 20636 22260 20692 22270
rect 20636 22166 20692 22204
rect 20748 22260 20804 22270
rect 20748 22258 20916 22260
rect 20748 22206 20750 22258
rect 20802 22206 20916 22258
rect 20748 22204 20916 22206
rect 20748 22194 20804 22204
rect 20524 21868 20692 21924
rect 20524 21700 20580 21710
rect 20524 21606 20580 21644
rect 20412 20962 20468 20972
rect 20636 20188 20692 21868
rect 20860 21810 20916 22204
rect 20860 21758 20862 21810
rect 20914 21758 20916 21810
rect 20860 21746 20916 21758
rect 20972 21810 21028 23212
rect 22002 22764 22266 22774
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22002 22698 22266 22708
rect 20972 21758 20974 21810
rect 21026 21758 21028 21810
rect 20972 21746 21028 21758
rect 21420 22372 21476 22382
rect 20524 20132 20692 20188
rect 20748 21698 20804 21710
rect 20748 21646 20750 21698
rect 20802 21646 20804 21698
rect 20524 19348 20580 20132
rect 20636 20020 20692 20030
rect 20748 20020 20804 21646
rect 21196 21586 21252 21598
rect 21196 21534 21198 21586
rect 21250 21534 21252 21586
rect 21196 20692 21252 21534
rect 21196 20626 21252 20636
rect 21420 20578 21476 22316
rect 21532 22370 21588 22382
rect 21532 22318 21534 22370
rect 21586 22318 21588 22370
rect 21532 20804 21588 22318
rect 22204 22260 22260 22270
rect 22204 22166 22260 22204
rect 21980 21812 22036 21822
rect 21644 21700 21700 21710
rect 21644 21606 21700 21644
rect 21756 21586 21812 21598
rect 21756 21534 21758 21586
rect 21810 21534 21812 21586
rect 21756 21476 21812 21534
rect 21980 21586 22036 21756
rect 21980 21534 21982 21586
rect 22034 21534 22036 21586
rect 21980 21522 22036 21534
rect 22652 21812 22708 21822
rect 21756 21410 21812 21420
rect 22002 21196 22266 21206
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22002 21130 22266 21140
rect 22540 21028 22596 21038
rect 22540 20934 22596 20972
rect 22652 20914 22708 21756
rect 22764 21474 22820 23884
rect 22988 23380 23044 23390
rect 22988 23286 23044 23324
rect 22764 21422 22766 21474
rect 22818 21422 22820 21474
rect 22764 21410 22820 21422
rect 22652 20862 22654 20914
rect 22706 20862 22708 20914
rect 22652 20850 22708 20862
rect 22876 20804 22932 20814
rect 21588 20748 21700 20804
rect 21532 20738 21588 20748
rect 21420 20526 21422 20578
rect 21474 20526 21476 20578
rect 21084 20020 21140 20030
rect 20748 19964 21084 20020
rect 20636 19926 20692 19964
rect 21084 19926 21140 19964
rect 20524 19282 20580 19292
rect 21308 17780 21364 17790
rect 20636 17444 20692 17454
rect 20636 16994 20692 17388
rect 20636 16942 20638 16994
rect 20690 16942 20692 16994
rect 20636 16930 20692 16942
rect 21308 16882 21364 17724
rect 21308 16830 21310 16882
rect 21362 16830 21364 16882
rect 21308 16818 21364 16830
rect 20076 15428 20132 16716
rect 21420 16660 21476 20526
rect 21532 19908 21588 19918
rect 21532 19814 21588 19852
rect 21644 19236 21700 20748
rect 22876 20710 22932 20748
rect 22204 20132 22260 20142
rect 22204 20018 22260 20076
rect 22204 19966 22206 20018
rect 22258 19966 22260 20018
rect 22204 19954 22260 19966
rect 22988 20020 23044 20030
rect 22988 19926 23044 19964
rect 21868 19908 21924 19918
rect 21868 19814 21924 19852
rect 22204 19796 22260 19806
rect 22204 19794 22484 19796
rect 22204 19742 22206 19794
rect 22258 19742 22484 19794
rect 22204 19740 22484 19742
rect 22204 19730 22260 19740
rect 22002 19628 22266 19638
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22002 19562 22266 19572
rect 22316 19348 22372 19358
rect 22428 19348 22484 19740
rect 22316 19346 22484 19348
rect 22316 19294 22318 19346
rect 22370 19294 22484 19346
rect 22316 19292 22484 19294
rect 22316 19282 22372 19292
rect 21644 19234 21812 19236
rect 21644 19182 21646 19234
rect 21698 19182 21812 19234
rect 21644 19180 21812 19182
rect 21644 19170 21700 19180
rect 21308 16604 21476 16660
rect 21644 18676 21700 18686
rect 21644 18338 21700 18620
rect 21644 18286 21646 18338
rect 21698 18286 21700 18338
rect 20972 15988 21028 15998
rect 20636 15932 20972 15988
rect 20188 15428 20244 15438
rect 20076 15426 20244 15428
rect 20076 15374 20190 15426
rect 20242 15374 20244 15426
rect 20076 15372 20244 15374
rect 20076 15148 20132 15372
rect 20188 15362 20244 15372
rect 19628 14366 19630 14418
rect 19682 14366 19684 14418
rect 19628 14354 19684 14366
rect 19964 15092 20132 15148
rect 19964 14420 20020 15092
rect 20636 14642 20692 15932
rect 20972 15922 21028 15932
rect 21308 15148 21364 16604
rect 21644 16212 21700 18286
rect 21756 17780 21812 19180
rect 22876 19124 22932 19134
rect 22876 18452 22932 19068
rect 22876 18358 22932 18396
rect 23212 18562 23268 25228
rect 23436 24722 23492 25676
rect 23436 24670 23438 24722
rect 23490 24670 23492 24722
rect 23436 24658 23492 24670
rect 23436 23938 23492 23950
rect 23436 23886 23438 23938
rect 23490 23886 23492 23938
rect 23436 23828 23492 23886
rect 23772 23940 23828 27022
rect 24220 27074 24276 27086
rect 24220 27022 24222 27074
rect 24274 27022 24276 27074
rect 24108 26962 24164 26974
rect 24108 26910 24110 26962
rect 24162 26910 24164 26962
rect 24108 26180 24164 26910
rect 24108 26114 24164 26124
rect 24220 24724 24276 27022
rect 26160 26684 26424 26694
rect 26216 26628 26264 26684
rect 26320 26628 26368 26684
rect 26160 26618 26424 26628
rect 34476 26684 34740 26694
rect 34532 26628 34580 26684
rect 34636 26628 34684 26684
rect 34476 26618 34740 26628
rect 25676 26516 25732 26526
rect 25676 26514 26404 26516
rect 25676 26462 25678 26514
rect 25730 26462 26404 26514
rect 25676 26460 26404 26462
rect 25676 26450 25732 26460
rect 25340 26402 25396 26414
rect 25340 26350 25342 26402
rect 25394 26350 25396 26402
rect 25228 25394 25284 25406
rect 25228 25342 25230 25394
rect 25282 25342 25284 25394
rect 25228 25284 25284 25342
rect 25340 25396 25396 26350
rect 25340 25330 25396 25340
rect 25564 26290 25620 26302
rect 25564 26238 25566 26290
rect 25618 26238 25620 26290
rect 25228 25218 25284 25228
rect 24332 24948 24388 24958
rect 24388 24892 24612 24948
rect 24332 24854 24388 24892
rect 24220 24668 24388 24724
rect 24220 23940 24276 23950
rect 23772 23874 23828 23884
rect 23884 23938 24276 23940
rect 23884 23886 24222 23938
rect 24274 23886 24276 23938
rect 23884 23884 24276 23886
rect 23436 23762 23492 23772
rect 23884 23380 23940 23884
rect 24220 23874 24276 23884
rect 24332 23828 24388 24668
rect 24556 23938 24612 24892
rect 24668 24834 24724 24846
rect 24668 24782 24670 24834
rect 24722 24782 24724 24834
rect 24668 24724 24724 24782
rect 24668 24658 24724 24668
rect 25564 24724 25620 26238
rect 25788 26290 25844 26302
rect 25788 26238 25790 26290
rect 25842 26238 25844 26290
rect 25788 25396 25844 26238
rect 25564 24658 25620 24668
rect 25676 25340 25788 25396
rect 24556 23886 24558 23938
rect 24610 23886 24612 23938
rect 24556 23874 24612 23886
rect 25564 23940 25620 23950
rect 25564 23846 25620 23884
rect 24332 23762 24388 23772
rect 24780 23716 24836 23726
rect 24780 23622 24836 23660
rect 25228 23716 25284 23726
rect 23884 23286 23940 23324
rect 24668 23380 24724 23390
rect 24668 23286 24724 23324
rect 23548 23266 23604 23278
rect 23548 23214 23550 23266
rect 23602 23214 23604 23266
rect 23548 21700 23604 23214
rect 24444 23156 24500 23166
rect 24444 23062 24500 23100
rect 25228 23154 25284 23660
rect 25676 23380 25732 25340
rect 25788 25330 25844 25340
rect 25900 25506 25956 25518
rect 25900 25454 25902 25506
rect 25954 25454 25956 25506
rect 25900 24836 25956 25454
rect 26348 25506 26404 26460
rect 30318 25900 30582 25910
rect 30374 25844 30422 25900
rect 30478 25844 30526 25900
rect 30318 25834 30582 25844
rect 26348 25454 26350 25506
rect 26402 25454 26404 25506
rect 26348 25442 26404 25454
rect 26572 25394 26628 25406
rect 26572 25342 26574 25394
rect 26626 25342 26628 25394
rect 26160 25116 26424 25126
rect 26216 25060 26264 25116
rect 26320 25060 26368 25116
rect 26160 25050 26424 25060
rect 26572 24836 26628 25342
rect 26908 25396 26964 25406
rect 26908 25302 26964 25340
rect 27356 25396 27412 25406
rect 27356 25302 27412 25340
rect 27580 25396 27636 25406
rect 27580 25394 28084 25396
rect 27580 25342 27582 25394
rect 27634 25342 28084 25394
rect 27580 25340 28084 25342
rect 27580 25330 27636 25340
rect 26684 25284 26740 25294
rect 26684 25190 26740 25228
rect 27468 25282 27524 25294
rect 27468 25230 27470 25282
rect 27522 25230 27524 25282
rect 27468 24948 27524 25230
rect 27468 24882 27524 24892
rect 25900 24770 25956 24780
rect 26012 24780 26628 24836
rect 26012 24724 26068 24780
rect 25228 23102 25230 23154
rect 25282 23102 25284 23154
rect 25228 23090 25284 23102
rect 25452 23268 25508 23278
rect 25452 23154 25508 23212
rect 25452 23102 25454 23154
rect 25506 23102 25508 23154
rect 25452 23090 25508 23102
rect 24444 22482 24500 22494
rect 24444 22430 24446 22482
rect 24498 22430 24500 22482
rect 24444 21812 24500 22430
rect 25564 22372 25620 22382
rect 25676 22372 25732 23324
rect 25788 24052 25844 24062
rect 25788 23378 25844 23996
rect 25788 23326 25790 23378
rect 25842 23326 25844 23378
rect 25788 23314 25844 23326
rect 25564 22370 25732 22372
rect 25564 22318 25566 22370
rect 25618 22318 25732 22370
rect 25564 22316 25732 22318
rect 25788 22484 25844 22494
rect 25564 22306 25620 22316
rect 25676 22148 25732 22158
rect 25676 22054 25732 22092
rect 24444 21718 24500 21756
rect 25452 21812 25508 21822
rect 25452 21718 25508 21756
rect 23548 21634 23604 21644
rect 25564 21700 25620 21710
rect 25788 21700 25844 22428
rect 25564 21698 25844 21700
rect 25564 21646 25566 21698
rect 25618 21646 25844 21698
rect 25564 21644 25844 21646
rect 25900 22146 25956 22158
rect 25900 22094 25902 22146
rect 25954 22094 25956 22146
rect 25564 21634 25620 21644
rect 23884 21588 23940 21598
rect 23884 21494 23940 21532
rect 24444 21586 24500 21598
rect 24444 21534 24446 21586
rect 24498 21534 24500 21586
rect 24444 20916 24500 21534
rect 24444 20850 24500 20860
rect 24556 21476 24612 21486
rect 24668 21476 24724 21486
rect 24612 21474 24724 21476
rect 24612 21422 24670 21474
rect 24722 21422 24724 21474
rect 24612 21420 24724 21422
rect 23772 20692 23828 20702
rect 23772 20690 24388 20692
rect 23772 20638 23774 20690
rect 23826 20638 24388 20690
rect 23772 20636 24388 20638
rect 23772 20626 23828 20636
rect 23212 18510 23214 18562
rect 23266 18510 23268 18562
rect 22540 18340 22596 18350
rect 22002 18060 22266 18070
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22002 17994 22266 18004
rect 21756 17714 21812 17724
rect 22540 17442 22596 18284
rect 23212 18228 23268 18510
rect 23212 18162 23268 18172
rect 23436 20132 23492 20142
rect 22540 17390 22542 17442
rect 22594 17390 22596 17442
rect 21644 16146 21700 16156
rect 21756 16770 21812 16782
rect 21756 16718 21758 16770
rect 21810 16718 21812 16770
rect 21756 16100 21812 16718
rect 22540 16772 22596 17390
rect 22540 16706 22596 16716
rect 21756 16034 21812 16044
rect 21868 16660 21924 16670
rect 21868 16098 21924 16604
rect 22876 16660 22932 16670
rect 22002 16492 22266 16502
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22002 16426 22266 16436
rect 21868 16046 21870 16098
rect 21922 16046 21924 16098
rect 21868 16034 21924 16046
rect 22428 16100 22484 16110
rect 22428 16006 22484 16044
rect 21532 15988 21588 15998
rect 21532 15894 21588 15932
rect 22204 15986 22260 15998
rect 22204 15934 22206 15986
rect 22258 15934 22260 15986
rect 20636 14590 20638 14642
rect 20690 14590 20692 14642
rect 20636 14578 20692 14590
rect 21196 15092 21364 15148
rect 21644 15874 21700 15886
rect 21644 15822 21646 15874
rect 21698 15822 21700 15874
rect 20748 14530 20804 14542
rect 20748 14478 20750 14530
rect 20802 14478 20804 14530
rect 19964 14354 20020 14364
rect 20076 14418 20132 14430
rect 20076 14366 20078 14418
rect 20130 14366 20132 14418
rect 19852 14308 19908 14318
rect 19516 13906 19572 13916
rect 19740 14306 19908 14308
rect 19740 14254 19854 14306
rect 19906 14254 19908 14306
rect 19740 14252 19908 14254
rect 19628 13860 19684 13870
rect 19628 13746 19684 13804
rect 19628 13694 19630 13746
rect 19682 13694 19684 13746
rect 19628 13682 19684 13694
rect 19740 13748 19796 14252
rect 19852 14242 19908 14252
rect 19852 14084 19908 14094
rect 19852 13970 19908 14028
rect 20076 13972 20132 14366
rect 20300 14308 20356 14318
rect 20524 14308 20580 14318
rect 20300 14306 20468 14308
rect 20300 14254 20302 14306
rect 20354 14254 20468 14306
rect 20300 14252 20468 14254
rect 20300 14242 20356 14252
rect 19852 13918 19854 13970
rect 19906 13918 19908 13970
rect 19852 13906 19908 13918
rect 19964 13916 20076 13972
rect 19740 13682 19796 13692
rect 19516 13524 19572 13534
rect 19516 12962 19572 13468
rect 19516 12910 19518 12962
rect 19570 12910 19572 12962
rect 19516 12898 19572 12910
rect 19852 12850 19908 12862
rect 19852 12798 19854 12850
rect 19906 12798 19908 12850
rect 19292 12738 19348 12750
rect 19292 12686 19294 12738
rect 19346 12686 19348 12738
rect 19292 12068 19348 12686
rect 19404 12738 19460 12750
rect 19404 12686 19406 12738
rect 19458 12686 19460 12738
rect 19404 12292 19460 12686
rect 19740 12740 19796 12750
rect 19740 12646 19796 12684
rect 19404 12226 19460 12236
rect 19852 12068 19908 12798
rect 19964 12628 20020 13916
rect 20076 13906 20132 13916
rect 20300 13860 20356 13870
rect 20188 13748 20244 13758
rect 20188 13654 20244 13692
rect 20300 13188 20356 13804
rect 20300 13094 20356 13132
rect 20076 13076 20132 13086
rect 20076 12982 20132 13020
rect 20412 12964 20468 14252
rect 20524 14214 20580 14252
rect 20524 13860 20580 13870
rect 20748 13860 20804 14478
rect 20524 13858 20804 13860
rect 20524 13806 20526 13858
rect 20578 13806 20804 13858
rect 20524 13804 20804 13806
rect 20524 13794 20580 13804
rect 20748 13076 20804 13804
rect 20524 12964 20580 12974
rect 20412 12908 20524 12964
rect 20524 12870 20580 12908
rect 20748 12628 20804 13020
rect 21196 14084 21252 15092
rect 21308 14644 21364 14654
rect 21644 14644 21700 15822
rect 22204 15148 22260 15934
rect 22652 15988 22708 15998
rect 22652 15894 22708 15932
rect 22764 15986 22820 15998
rect 22764 15934 22766 15986
rect 22818 15934 22820 15986
rect 21308 14642 21476 14644
rect 21308 14590 21310 14642
rect 21362 14590 21476 14642
rect 21308 14588 21476 14590
rect 21308 14578 21364 14588
rect 19964 12572 20132 12628
rect 19292 12012 19908 12068
rect 19068 11506 19180 11508
rect 19068 11454 19070 11506
rect 19122 11454 19180 11506
rect 19068 11452 19180 11454
rect 19068 11442 19124 11452
rect 19180 11414 19236 11452
rect 19628 11732 19684 11742
rect 19404 11396 19460 11406
rect 19292 11394 19460 11396
rect 19292 11342 19406 11394
rect 19458 11342 19460 11394
rect 19292 11340 19460 11342
rect 19292 11284 19348 11340
rect 19404 11330 19460 11340
rect 19628 11394 19684 11676
rect 19852 11620 19908 12012
rect 19852 11554 19908 11564
rect 19964 12404 20020 12414
rect 19628 11342 19630 11394
rect 19682 11342 19684 11394
rect 19628 11330 19684 11342
rect 19852 11396 19908 11406
rect 19964 11396 20020 12348
rect 20076 11732 20132 12572
rect 20748 12562 20804 12572
rect 20860 12962 20916 12974
rect 20860 12910 20862 12962
rect 20914 12910 20916 12962
rect 20636 12404 20692 12414
rect 20636 12310 20692 12348
rect 20860 12180 20916 12910
rect 20972 12740 21028 12750
rect 20972 12402 21028 12684
rect 21196 12516 21252 14028
rect 21420 14308 21476 14588
rect 21644 14578 21700 14588
rect 21868 15092 22260 15148
rect 21308 13524 21364 13534
rect 21420 13524 21476 14252
rect 21644 13524 21700 13534
rect 21420 13468 21644 13524
rect 21308 13430 21364 13468
rect 21644 13458 21700 13468
rect 21756 13522 21812 13534
rect 21756 13470 21758 13522
rect 21810 13470 21812 13522
rect 21756 13076 21812 13470
rect 21756 13010 21812 13020
rect 21868 12964 21924 15092
rect 22002 14924 22266 14934
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22002 14858 22266 14868
rect 22204 13972 22260 13982
rect 22204 13746 22260 13916
rect 22204 13694 22206 13746
rect 22258 13694 22260 13746
rect 22204 13682 22260 13694
rect 22652 13746 22708 13758
rect 22652 13694 22654 13746
rect 22706 13694 22708 13746
rect 21980 13524 22036 13562
rect 21980 13458 22036 13468
rect 22002 13356 22266 13366
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22002 13290 22266 13300
rect 22092 13188 22148 13198
rect 22092 13094 22148 13132
rect 22652 13188 22708 13694
rect 22652 13122 22708 13132
rect 22428 13076 22484 13086
rect 21868 12870 21924 12908
rect 22316 12964 22372 12974
rect 21644 12852 21700 12862
rect 21700 12796 21812 12852
rect 21644 12758 21700 12796
rect 21196 12460 21700 12516
rect 20972 12350 20974 12402
rect 21026 12350 21028 12402
rect 20972 12338 21028 12350
rect 21308 12348 21588 12404
rect 21308 12180 21364 12348
rect 20860 12124 21364 12180
rect 21420 12178 21476 12190
rect 21420 12126 21422 12178
rect 21474 12126 21476 12178
rect 20300 12068 20356 12078
rect 20076 11666 20132 11676
rect 20188 12066 20580 12068
rect 20188 12014 20302 12066
rect 20354 12014 20580 12066
rect 20188 12012 20580 12014
rect 19852 11394 20020 11396
rect 19852 11342 19854 11394
rect 19906 11342 20020 11394
rect 19852 11340 20020 11342
rect 20076 11396 20132 11406
rect 20188 11396 20244 12012
rect 20300 12002 20356 12012
rect 20412 11620 20468 11630
rect 20412 11526 20468 11564
rect 20524 11506 20580 12012
rect 20524 11454 20526 11506
rect 20578 11454 20580 11506
rect 20524 11442 20580 11454
rect 21308 11732 21364 11742
rect 20076 11394 20244 11396
rect 20076 11342 20078 11394
rect 20130 11342 20244 11394
rect 20076 11340 20244 11342
rect 19852 11330 19908 11340
rect 20076 11330 20132 11340
rect 18844 11228 19348 11284
rect 18172 9102 18174 9154
rect 18226 9102 18228 9154
rect 18172 9090 18228 9102
rect 18284 9602 18340 9614
rect 18284 9550 18286 9602
rect 18338 9550 18340 9602
rect 17724 8930 17780 8988
rect 17724 8878 17726 8930
rect 17778 8878 17780 8930
rect 17724 8866 17780 8878
rect 17948 8932 18004 8942
rect 17948 8372 18004 8876
rect 17948 8370 18228 8372
rect 17948 8318 17950 8370
rect 18002 8318 18228 8370
rect 17948 8316 18228 8318
rect 17948 8306 18004 8316
rect 16716 7858 16772 7868
rect 17164 8034 17220 8046
rect 17164 7982 17166 8034
rect 17218 7982 17220 8034
rect 16268 7588 16324 7598
rect 16268 7586 16436 7588
rect 16268 7534 16270 7586
rect 16322 7534 16436 7586
rect 16268 7532 16436 7534
rect 16268 7522 16324 7532
rect 16156 5814 16212 5852
rect 16380 5796 16436 7532
rect 16828 7476 16884 7486
rect 16828 7382 16884 7420
rect 17164 6692 17220 7982
rect 17844 7868 18108 7878
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 17844 7802 18108 7812
rect 18060 7476 18116 7486
rect 18172 7476 18228 8316
rect 18060 7474 18228 7476
rect 18060 7422 18062 7474
rect 18114 7422 18228 7474
rect 18060 7420 18228 7422
rect 18060 7410 18116 7420
rect 17388 7364 17444 7374
rect 17388 7362 17556 7364
rect 17388 7310 17390 7362
rect 17442 7310 17556 7362
rect 17388 7308 17556 7310
rect 17388 7298 17444 7308
rect 17164 6626 17220 6636
rect 17388 6020 17444 6030
rect 17388 5926 17444 5964
rect 16716 5796 16772 5806
rect 16380 5794 16772 5796
rect 16380 5742 16718 5794
rect 16770 5742 16772 5794
rect 16380 5740 16772 5742
rect 15484 4174 15486 4226
rect 15538 4174 15540 4226
rect 15484 4162 15540 4174
rect 15596 5122 15988 5124
rect 15596 5070 15934 5122
rect 15986 5070 15988 5122
rect 15596 5068 15988 5070
rect 15372 3602 15428 3612
rect 15484 3668 15540 3678
rect 15596 3668 15652 5068
rect 15932 5058 15988 5068
rect 16268 5684 16324 5694
rect 16268 4564 16324 5628
rect 16268 4498 16324 4508
rect 16716 4340 16772 5740
rect 17500 5796 17556 7308
rect 18172 6802 18228 7420
rect 18284 8258 18340 9550
rect 18284 8206 18286 8258
rect 18338 8206 18340 8258
rect 18284 7474 18340 8206
rect 18284 7422 18286 7474
rect 18338 7422 18340 7474
rect 18284 7410 18340 7422
rect 18732 7476 18788 11228
rect 19740 11170 19796 11182
rect 19740 11118 19742 11170
rect 19794 11118 19796 11170
rect 19180 10498 19236 10510
rect 19180 10446 19182 10498
rect 19234 10446 19236 10498
rect 18732 7410 18788 7420
rect 18844 10164 18900 10174
rect 18844 7474 18900 10108
rect 19180 9940 19236 10446
rect 19740 10052 19796 11118
rect 21308 10498 21364 11676
rect 21308 10446 21310 10498
rect 21362 10446 21364 10498
rect 21308 10434 21364 10446
rect 19740 9986 19796 9996
rect 20972 10164 21028 10174
rect 19180 9874 19236 9884
rect 20076 9828 20132 9838
rect 20076 9734 20132 9772
rect 20636 9828 20692 9838
rect 20636 9734 20692 9772
rect 18956 9716 19012 9726
rect 18956 9622 19012 9660
rect 19628 9714 19684 9726
rect 19628 9662 19630 9714
rect 19682 9662 19684 9714
rect 18956 9154 19012 9166
rect 18956 9102 18958 9154
rect 19010 9102 19012 9154
rect 18956 8932 19012 9102
rect 19068 9044 19124 9054
rect 19628 9044 19684 9662
rect 19068 9042 19684 9044
rect 19068 8990 19070 9042
rect 19122 8990 19684 9042
rect 19068 8988 19684 8990
rect 20972 9042 21028 10108
rect 21420 10164 21476 12126
rect 21532 11506 21588 12348
rect 21532 11454 21534 11506
rect 21586 11454 21588 11506
rect 21532 11442 21588 11454
rect 21644 10612 21700 12460
rect 21756 11844 21812 12796
rect 22092 12738 22148 12750
rect 22092 12686 22094 12738
rect 22146 12686 22148 12738
rect 22092 12290 22148 12686
rect 22316 12628 22372 12908
rect 22316 12562 22372 12572
rect 22092 12238 22094 12290
rect 22146 12238 22148 12290
rect 22092 12226 22148 12238
rect 22428 12068 22484 13020
rect 22764 13076 22820 15934
rect 22876 13970 22932 16604
rect 23436 16660 23492 20076
rect 23996 20130 24052 20142
rect 23996 20078 23998 20130
rect 24050 20078 24052 20130
rect 23996 19348 24052 20078
rect 24332 19906 24388 20636
rect 24444 20132 24500 20142
rect 24444 20038 24500 20076
rect 24332 19854 24334 19906
rect 24386 19854 24388 19906
rect 24332 19842 24388 19854
rect 24556 19348 24612 21420
rect 24668 21410 24724 21420
rect 25452 21364 25508 21374
rect 25452 21270 25508 21308
rect 24668 20020 24724 20030
rect 24668 19926 24724 19964
rect 25228 20020 25284 20030
rect 25228 19926 25284 19964
rect 25676 19906 25732 21644
rect 25900 21252 25956 22094
rect 26012 22148 26068 24668
rect 26460 24612 26516 24622
rect 26460 24610 26740 24612
rect 26460 24558 26462 24610
rect 26514 24558 26740 24610
rect 26460 24556 26740 24558
rect 26460 24546 26516 24556
rect 26460 24052 26516 24062
rect 26516 23996 26628 24052
rect 26460 23986 26516 23996
rect 26124 23828 26180 23838
rect 26124 23714 26180 23772
rect 26124 23662 26126 23714
rect 26178 23662 26180 23714
rect 26124 23650 26180 23662
rect 26160 23548 26424 23558
rect 26216 23492 26264 23548
rect 26320 23492 26368 23548
rect 26160 23482 26424 23492
rect 26124 23156 26180 23166
rect 26124 22596 26180 23100
rect 26124 22502 26180 22540
rect 26460 22596 26516 22606
rect 26572 22596 26628 23996
rect 26460 22594 26628 22596
rect 26460 22542 26462 22594
rect 26514 22542 26628 22594
rect 26460 22540 26628 22542
rect 26684 23940 26740 24556
rect 26460 22530 26516 22540
rect 26684 22482 26740 23884
rect 27916 24052 27972 24062
rect 27916 23938 27972 23996
rect 28028 24050 28084 25340
rect 28140 25284 28196 25294
rect 28140 25282 28308 25284
rect 28140 25230 28142 25282
rect 28194 25230 28308 25282
rect 28140 25228 28308 25230
rect 28140 25218 28196 25228
rect 28028 23998 28030 24050
rect 28082 23998 28084 24050
rect 28028 23986 28084 23998
rect 27916 23886 27918 23938
rect 27970 23886 27972 23938
rect 27916 23874 27972 23886
rect 28140 23940 28196 23950
rect 28140 23846 28196 23884
rect 27132 23828 27188 23838
rect 27132 23734 27188 23772
rect 26796 23716 26852 23726
rect 26796 23042 26852 23660
rect 27020 23714 27076 23726
rect 27020 23662 27022 23714
rect 27074 23662 27076 23714
rect 27020 23268 27076 23662
rect 27244 23716 27300 23726
rect 27244 23622 27300 23660
rect 27468 23716 27524 23726
rect 28252 23716 28308 25228
rect 34476 25116 34740 25126
rect 34532 25060 34580 25116
rect 34636 25060 34684 25116
rect 34476 25050 34740 25060
rect 28700 24948 28756 24958
rect 28700 24834 28756 24892
rect 28700 24782 28702 24834
rect 28754 24782 28756 24834
rect 28700 24770 28756 24782
rect 29372 24836 29428 24846
rect 29372 24722 29428 24780
rect 29372 24670 29374 24722
rect 29426 24670 29428 24722
rect 29372 24658 29428 24670
rect 30044 24836 30100 24846
rect 29372 24052 29428 24062
rect 29148 23828 29204 23838
rect 29148 23734 29204 23772
rect 29372 23826 29428 23996
rect 29372 23774 29374 23826
rect 29426 23774 29428 23826
rect 29372 23762 29428 23774
rect 28364 23716 28420 23726
rect 28252 23660 28364 23716
rect 27020 23202 27076 23212
rect 27468 23044 27524 23660
rect 28364 23622 28420 23660
rect 29260 23714 29316 23726
rect 29260 23662 29262 23714
rect 29314 23662 29316 23714
rect 29148 23268 29204 23278
rect 29260 23268 29316 23662
rect 29932 23716 29988 23726
rect 29932 23622 29988 23660
rect 29148 23266 29316 23268
rect 29148 23214 29150 23266
rect 29202 23214 29316 23266
rect 29148 23212 29316 23214
rect 29148 23202 29204 23212
rect 30044 23156 30100 24780
rect 30318 24332 30582 24342
rect 30374 24276 30422 24332
rect 30478 24276 30526 24332
rect 30318 24266 30582 24276
rect 34476 23548 34740 23558
rect 34532 23492 34580 23548
rect 34636 23492 34684 23548
rect 34476 23482 34740 23492
rect 26796 22990 26798 23042
rect 26850 22990 26852 23042
rect 26796 22978 26852 22990
rect 27020 22988 27524 23044
rect 29708 23154 30100 23156
rect 29708 23102 30046 23154
rect 30098 23102 30100 23154
rect 29708 23100 30100 23102
rect 26684 22430 26686 22482
rect 26738 22430 26740 22482
rect 26684 22418 26740 22430
rect 26908 22596 26964 22606
rect 26908 22370 26964 22540
rect 26908 22318 26910 22370
rect 26962 22318 26964 22370
rect 26908 22306 26964 22318
rect 26124 22148 26180 22158
rect 26012 22092 26124 22148
rect 26124 22082 26180 22092
rect 26160 21980 26424 21990
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26160 21914 26424 21924
rect 26684 21812 26740 21822
rect 26124 21588 26180 21598
rect 26124 21474 26180 21532
rect 26124 21422 26126 21474
rect 26178 21422 26180 21474
rect 26124 21410 26180 21422
rect 25900 21186 25956 21196
rect 26012 20916 26068 20926
rect 25900 20860 26012 20916
rect 25900 20018 25956 20860
rect 26012 20822 26068 20860
rect 26160 20412 26424 20422
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26160 20346 26424 20356
rect 25900 19966 25902 20018
rect 25954 19966 25956 20018
rect 25900 19954 25956 19966
rect 26684 20242 26740 21756
rect 27020 21812 27076 22988
rect 27132 22484 27188 22494
rect 27132 22390 27188 22428
rect 27916 22372 27972 22382
rect 27468 22370 27972 22372
rect 27468 22318 27918 22370
rect 27970 22318 27972 22370
rect 27468 22316 27972 22318
rect 27244 22148 27300 22158
rect 27244 22054 27300 22092
rect 27468 22146 27524 22316
rect 27916 22306 27972 22316
rect 27804 22148 27860 22158
rect 27468 22094 27470 22146
rect 27522 22094 27524 22146
rect 27468 21924 27524 22094
rect 27020 21746 27076 21756
rect 27244 21868 27524 21924
rect 27580 22146 27860 22148
rect 27580 22094 27806 22146
rect 27858 22094 27860 22146
rect 27580 22092 27860 22094
rect 27244 21588 27300 21868
rect 27580 21700 27636 22092
rect 27804 22082 27860 22092
rect 27244 21522 27300 21532
rect 27356 21644 27636 21700
rect 27020 21364 27076 21374
rect 27020 20802 27076 21308
rect 27020 20750 27022 20802
rect 27074 20750 27076 20802
rect 27020 20738 27076 20750
rect 27356 20802 27412 21644
rect 29708 21586 29764 23100
rect 30044 23090 30100 23100
rect 30318 22764 30582 22774
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30318 22698 30582 22708
rect 34476 21980 34740 21990
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34476 21914 34740 21924
rect 29708 21534 29710 21586
rect 29762 21534 29764 21586
rect 27468 21476 27524 21486
rect 27468 20914 27524 21420
rect 28812 21476 28868 21486
rect 28812 21382 28868 21420
rect 27468 20862 27470 20914
rect 27522 20862 27524 20914
rect 27468 20850 27524 20862
rect 27580 21252 27636 21262
rect 27356 20750 27358 20802
rect 27410 20750 27412 20802
rect 27356 20738 27412 20750
rect 27580 20802 27636 21196
rect 27580 20750 27582 20802
rect 27634 20750 27636 20802
rect 27580 20738 27636 20750
rect 26684 20190 26686 20242
rect 26738 20190 26740 20242
rect 25676 19854 25678 19906
rect 25730 19854 25732 19906
rect 25676 19842 25732 19854
rect 26684 19796 26740 20190
rect 29708 20132 29764 21534
rect 30318 21196 30582 21206
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30318 21130 30582 21140
rect 34476 20412 34740 20422
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34476 20346 34740 20356
rect 29708 20066 29764 20076
rect 30604 20132 30660 20142
rect 27132 20020 27188 20030
rect 27132 19926 27188 19964
rect 29148 20020 29204 20030
rect 27804 19906 27860 19918
rect 27804 19854 27806 19906
rect 27858 19854 27860 19906
rect 26684 19730 26740 19740
rect 27132 19794 27188 19806
rect 27132 19742 27134 19794
rect 27186 19742 27188 19794
rect 23996 19346 24612 19348
rect 23996 19294 24558 19346
rect 24610 19294 24612 19346
rect 23996 19292 24612 19294
rect 24556 19282 24612 19292
rect 26460 19348 26516 19358
rect 26460 19254 26516 19292
rect 27132 19348 27188 19742
rect 27132 19282 27188 19292
rect 27468 19794 27524 19806
rect 27468 19742 27470 19794
rect 27522 19742 27524 19794
rect 25676 19234 25732 19246
rect 25676 19182 25678 19234
rect 25730 19182 25732 19234
rect 23548 18452 23604 18462
rect 25676 18452 25732 19182
rect 26160 18844 26424 18854
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26160 18778 26424 18788
rect 26684 18508 26852 18564
rect 26124 18452 26180 18462
rect 26684 18452 26740 18508
rect 23604 18396 23716 18452
rect 23548 18358 23604 18396
rect 23548 17780 23604 17790
rect 23548 17686 23604 17724
rect 23660 17556 23716 18396
rect 25452 18340 25508 18350
rect 25452 18246 25508 18284
rect 23436 16594 23492 16604
rect 23548 17500 23716 17556
rect 24556 17780 24612 17790
rect 23436 16212 23492 16222
rect 23436 16118 23492 16156
rect 23436 14644 23492 14654
rect 23436 14550 23492 14588
rect 22876 13918 22878 13970
rect 22930 13918 22932 13970
rect 22876 13906 22932 13918
rect 23548 13972 23604 17500
rect 24556 16884 24612 17724
rect 25340 16884 25396 16894
rect 25676 16884 25732 18396
rect 26012 18450 26180 18452
rect 26012 18398 26126 18450
rect 26178 18398 26180 18450
rect 26012 18396 26180 18398
rect 25900 18340 25956 18350
rect 24556 16882 24724 16884
rect 24556 16830 24558 16882
rect 24610 16830 24724 16882
rect 24556 16828 24724 16830
rect 24556 16818 24612 16828
rect 23884 16772 23940 16782
rect 23884 16770 24500 16772
rect 23884 16718 23886 16770
rect 23938 16718 24500 16770
rect 23884 16716 24500 16718
rect 23884 16706 23940 16716
rect 24444 16210 24500 16716
rect 24444 16158 24446 16210
rect 24498 16158 24500 16210
rect 24444 16146 24500 16158
rect 24556 16660 24612 16670
rect 23660 16100 23716 16110
rect 23660 16006 23716 16044
rect 24332 15988 24388 15998
rect 24332 15894 24388 15932
rect 24556 15986 24612 16604
rect 24556 15934 24558 15986
rect 24610 15934 24612 15986
rect 24556 15922 24612 15934
rect 23996 15874 24052 15886
rect 23996 15822 23998 15874
rect 24050 15822 24052 15874
rect 23996 15316 24052 15822
rect 23996 15250 24052 15260
rect 24668 15148 24724 16828
rect 25340 16882 25732 16884
rect 25340 16830 25342 16882
rect 25394 16830 25732 16882
rect 25340 16828 25732 16830
rect 25788 18338 25956 18340
rect 25788 18286 25902 18338
rect 25954 18286 25956 18338
rect 25788 18284 25956 18286
rect 25340 16818 25396 16828
rect 25788 16324 25844 18284
rect 25900 18274 25956 18284
rect 26012 17108 26068 18396
rect 26124 18386 26180 18396
rect 26572 18396 26740 18452
rect 26796 18450 26852 18508
rect 27132 18452 27188 18462
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26160 17276 26424 17286
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26160 17210 26424 17220
rect 26012 17052 26180 17108
rect 26012 16772 26068 16782
rect 25788 16258 25844 16268
rect 25900 16770 26068 16772
rect 25900 16718 26014 16770
rect 26066 16718 26068 16770
rect 25900 16716 26068 16718
rect 25900 15204 25956 16716
rect 26012 16706 26068 16716
rect 26124 16772 26180 17052
rect 26124 16706 26180 16716
rect 26236 16100 26292 16110
rect 26236 16006 26292 16044
rect 26124 15988 26180 15998
rect 26124 15894 26180 15932
rect 26012 15876 26068 15886
rect 26012 15782 26068 15820
rect 26160 15708 26424 15718
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26160 15642 26424 15652
rect 26124 15426 26180 15438
rect 26124 15374 26126 15426
rect 26178 15374 26180 15426
rect 26012 15204 26068 15214
rect 25900 15202 26068 15204
rect 25900 15150 26014 15202
rect 26066 15150 26068 15202
rect 25900 15148 26068 15150
rect 24220 15092 24724 15148
rect 26012 15138 26068 15148
rect 24220 14530 24276 15092
rect 24220 14478 24222 14530
rect 24274 14478 24276 14530
rect 24220 14466 24276 14478
rect 25452 14420 25508 14430
rect 23660 13972 23716 13982
rect 24220 13972 24276 13982
rect 23548 13970 24276 13972
rect 23548 13918 23662 13970
rect 23714 13918 24222 13970
rect 24274 13918 24276 13970
rect 23548 13916 24276 13918
rect 23660 13906 23716 13916
rect 24220 13906 24276 13916
rect 23548 13746 23604 13758
rect 23548 13694 23550 13746
rect 23602 13694 23604 13746
rect 22764 13010 22820 13020
rect 22988 13524 23044 13534
rect 22988 13074 23044 13468
rect 22988 13022 22990 13074
rect 23042 13022 23044 13074
rect 22988 13010 23044 13022
rect 22540 12852 22596 12862
rect 22876 12852 22932 12862
rect 22540 12850 22820 12852
rect 22540 12798 22542 12850
rect 22594 12798 22820 12850
rect 22540 12796 22820 12798
rect 22540 12786 22596 12796
rect 21756 11788 21924 11844
rect 21868 11396 21924 11788
rect 22002 11788 22266 11798
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22002 11722 22266 11732
rect 22428 11732 22484 12012
rect 22428 11676 22708 11732
rect 22428 11506 22484 11676
rect 22428 11454 22430 11506
rect 22482 11454 22484 11506
rect 22428 11442 22484 11454
rect 22540 11508 22596 11518
rect 21980 11396 22036 11406
rect 21868 11394 22036 11396
rect 21868 11342 21982 11394
rect 22034 11342 22036 11394
rect 21868 11340 22036 11342
rect 21980 11330 22036 11340
rect 22540 10836 22596 11452
rect 22652 11396 22708 11676
rect 22764 11620 22820 12796
rect 22876 12758 22932 12796
rect 22876 11620 22932 11630
rect 22764 11618 22932 11620
rect 22764 11566 22878 11618
rect 22930 11566 22932 11618
rect 22764 11564 22932 11566
rect 22876 11554 22932 11564
rect 22988 11396 23044 11406
rect 22652 11394 23044 11396
rect 22652 11342 22990 11394
rect 23042 11342 23044 11394
rect 22652 11340 23044 11342
rect 22988 11330 23044 11340
rect 22540 10742 22596 10780
rect 22092 10724 22148 10734
rect 22092 10630 22148 10668
rect 21420 10098 21476 10108
rect 21532 10556 21700 10612
rect 21756 10612 21812 10622
rect 21756 10610 21924 10612
rect 21756 10558 21758 10610
rect 21810 10558 21924 10610
rect 21756 10556 21924 10558
rect 21308 10052 21364 10062
rect 21308 9958 21364 9996
rect 21420 9940 21476 9950
rect 21420 9846 21476 9884
rect 21532 9716 21588 10556
rect 21756 10546 21812 10556
rect 20972 8990 20974 9042
rect 21026 8990 21028 9042
rect 19068 8978 19124 8988
rect 20972 8978 21028 8990
rect 21420 9714 21588 9716
rect 21420 9662 21534 9714
rect 21586 9662 21588 9714
rect 21420 9660 21588 9662
rect 18956 8866 19012 8876
rect 19068 8820 19124 8830
rect 19068 8370 19124 8764
rect 19068 8318 19070 8370
rect 19122 8318 19124 8370
rect 19068 8306 19124 8318
rect 21420 8370 21476 9660
rect 21532 9650 21588 9660
rect 21756 10386 21812 10398
rect 21756 10334 21758 10386
rect 21810 10334 21812 10386
rect 21756 9154 21812 10334
rect 21756 9102 21758 9154
rect 21810 9102 21812 9154
rect 21756 9090 21812 9102
rect 21868 9268 21924 10556
rect 23548 10276 23604 13694
rect 23884 13748 23940 13758
rect 23884 13654 23940 13692
rect 25452 13748 25508 14364
rect 26124 14308 26180 15374
rect 26348 15428 26404 15438
rect 26572 15428 26628 18396
rect 26796 18386 26852 18398
rect 26908 18450 27188 18452
rect 26908 18398 27134 18450
rect 27186 18398 27188 18450
rect 26908 18396 27188 18398
rect 26684 18228 26740 18238
rect 26684 17668 26740 18172
rect 26908 17668 26964 18396
rect 27132 18386 27188 18396
rect 27468 17780 27524 19742
rect 27804 19012 27860 19854
rect 28588 19346 28644 19358
rect 28588 19294 28590 19346
rect 28642 19294 28644 19346
rect 28028 19012 28084 19022
rect 27804 18956 28028 19012
rect 27468 17714 27524 17724
rect 26684 17666 26964 17668
rect 26684 17614 26686 17666
rect 26738 17614 26964 17666
rect 26684 17612 26964 17614
rect 26684 17602 26740 17612
rect 28028 16996 28084 18956
rect 28588 18004 28644 19294
rect 29148 19236 29204 19964
rect 30604 20020 30660 20076
rect 30604 20018 30772 20020
rect 30604 19966 30606 20018
rect 30658 19966 30772 20018
rect 30604 19964 30772 19966
rect 30604 19954 30660 19964
rect 29932 19908 29988 19918
rect 29708 19906 29988 19908
rect 29708 19854 29934 19906
rect 29986 19854 29988 19906
rect 29708 19852 29988 19854
rect 29148 19234 29652 19236
rect 29148 19182 29150 19234
rect 29202 19182 29652 19234
rect 29148 19180 29652 19182
rect 29148 19170 29204 19180
rect 29260 19010 29316 19022
rect 29260 18958 29262 19010
rect 29314 18958 29316 19010
rect 28588 17948 29204 18004
rect 29036 17780 29092 17790
rect 27580 16884 27636 16894
rect 27468 16324 27524 16334
rect 27468 16230 27524 16268
rect 27580 16098 27636 16828
rect 27580 16046 27582 16098
rect 27634 16046 27636 16098
rect 27580 16034 27636 16046
rect 27916 15988 27972 15998
rect 27916 15894 27972 15932
rect 27468 15876 27524 15886
rect 27468 15782 27524 15820
rect 28028 15876 28084 16940
rect 28924 17668 28980 17678
rect 28140 16772 28196 16782
rect 28196 16716 28420 16772
rect 28140 16678 28196 16716
rect 28252 15988 28308 15998
rect 28028 15810 28084 15820
rect 28140 15874 28196 15886
rect 28140 15822 28142 15874
rect 28194 15822 28196 15874
rect 26348 15426 26628 15428
rect 26348 15374 26350 15426
rect 26402 15374 26628 15426
rect 26348 15372 26628 15374
rect 28140 15428 28196 15822
rect 26348 15362 26404 15372
rect 28140 15362 28196 15372
rect 28028 15316 28084 15326
rect 27356 15204 27412 15214
rect 27244 14532 27300 14542
rect 27244 14438 27300 14476
rect 25788 14252 26180 14308
rect 25676 13860 25732 13870
rect 25676 13766 25732 13804
rect 25452 13654 25508 13692
rect 24780 13524 24836 13534
rect 24780 13074 24836 13468
rect 24780 13022 24782 13074
rect 24834 13022 24836 13074
rect 24780 13010 24836 13022
rect 24108 12964 24164 12974
rect 24108 12962 24500 12964
rect 24108 12910 24110 12962
rect 24162 12910 24500 12962
rect 24108 12908 24500 12910
rect 24108 12898 24164 12908
rect 24220 12068 24276 12078
rect 24220 11974 24276 12012
rect 24444 11394 24500 12908
rect 24444 11342 24446 11394
rect 24498 11342 24500 11394
rect 22002 10220 22266 10230
rect 23548 10220 23940 10276
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22002 10154 22266 10164
rect 23100 10052 23156 10062
rect 22092 9828 22148 9838
rect 22092 9734 22148 9772
rect 21868 8484 21924 9212
rect 23100 9716 23156 9996
rect 22002 8652 22266 8662
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22002 8586 22266 8596
rect 21868 8428 22372 8484
rect 21420 8318 21422 8370
rect 21474 8318 21476 8370
rect 18844 7422 18846 7474
rect 18898 7422 18900 7474
rect 18172 6750 18174 6802
rect 18226 6750 18228 6802
rect 18172 6738 18228 6750
rect 18732 6468 18788 6478
rect 18620 6466 18788 6468
rect 18620 6414 18734 6466
rect 18786 6414 18788 6466
rect 18620 6412 18788 6414
rect 17844 6300 18108 6310
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 17844 6234 18108 6244
rect 17948 6132 18004 6142
rect 17948 6038 18004 6076
rect 16940 5124 16996 5134
rect 16828 4340 16884 4350
rect 16716 4284 16828 4340
rect 16828 4274 16884 4284
rect 15484 3666 15652 3668
rect 15484 3614 15486 3666
rect 15538 3614 15652 3666
rect 15484 3612 15652 3614
rect 16940 3666 16996 5068
rect 17500 4788 17556 5740
rect 18284 5236 18340 5246
rect 18172 5124 18228 5134
rect 18172 5030 18228 5068
rect 17724 5012 17780 5022
rect 17724 4918 17780 4956
rect 17500 4732 17780 4788
rect 17276 4564 17332 4574
rect 17276 4470 17332 4508
rect 17612 4340 17668 4350
rect 17612 4246 17668 4284
rect 17724 4226 17780 4732
rect 17844 4732 18108 4742
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 17844 4666 18108 4676
rect 18060 4564 18116 4574
rect 18060 4338 18116 4508
rect 18060 4286 18062 4338
rect 18114 4286 18116 4338
rect 18060 4274 18116 4286
rect 17724 4174 17726 4226
rect 17778 4174 17780 4226
rect 17724 4162 17780 4174
rect 16940 3614 16942 3666
rect 16994 3614 16996 3666
rect 12572 3490 12628 3500
rect 14364 3556 14420 3566
rect 13244 3444 13300 3482
rect 14364 3462 14420 3500
rect 15484 3556 15540 3612
rect 16940 3602 16996 3614
rect 15484 3490 15540 3500
rect 13244 3378 13300 3388
rect 11676 3108 11732 3332
rect 11900 3266 11956 3276
rect 17844 3164 18108 3174
rect 11788 3108 11844 3118
rect 11676 3052 11788 3108
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 17844 3098 18108 3108
rect 11788 3042 11844 3052
rect 18284 2548 18340 5180
rect 18620 5012 18676 6412
rect 18732 6402 18788 6412
rect 18732 5906 18788 5918
rect 18732 5854 18734 5906
rect 18786 5854 18788 5906
rect 18732 5124 18788 5854
rect 18732 5058 18788 5068
rect 18620 4946 18676 4956
rect 18844 5012 18900 7422
rect 18956 8258 19012 8270
rect 18956 8206 18958 8258
rect 19010 8206 19012 8258
rect 18956 6132 19012 8206
rect 19180 7476 19236 7486
rect 19180 6804 19236 7420
rect 18956 6066 19012 6076
rect 19068 6748 19180 6804
rect 18844 4946 18900 4956
rect 19068 4564 19124 6748
rect 19180 6710 19236 6748
rect 19516 7362 19572 7374
rect 19516 7310 19518 7362
rect 19570 7310 19572 7362
rect 19516 6132 19572 7310
rect 19740 6804 19796 6814
rect 19740 6690 19796 6748
rect 19740 6638 19742 6690
rect 19794 6638 19796 6690
rect 19740 6626 19796 6638
rect 19516 6066 19572 6076
rect 21308 6132 21364 6142
rect 20076 6020 20132 6030
rect 19292 5908 19348 5918
rect 19292 5814 19348 5852
rect 20076 5906 20132 5964
rect 20524 6020 20580 6030
rect 20524 5926 20580 5964
rect 20972 6020 21028 6030
rect 20972 5926 21028 5964
rect 21308 6018 21364 6076
rect 21308 5966 21310 6018
rect 21362 5966 21364 6018
rect 21308 5954 21364 5966
rect 21420 6020 21476 8318
rect 21756 8036 21812 8046
rect 21644 7476 21700 7486
rect 21644 7362 21700 7420
rect 21644 7310 21646 7362
rect 21698 7310 21700 7362
rect 21644 7298 21700 7310
rect 20076 5854 20078 5906
rect 20130 5854 20132 5906
rect 20076 5842 20132 5854
rect 21420 5906 21476 5964
rect 21420 5854 21422 5906
rect 21474 5854 21476 5906
rect 21420 5842 21476 5854
rect 21532 7252 21588 7262
rect 21532 5908 21588 7196
rect 21756 6916 21812 7980
rect 21980 7474 22036 8428
rect 22316 8372 22372 8428
rect 22316 8370 22708 8372
rect 22316 8318 22318 8370
rect 22370 8318 22708 8370
rect 22316 8316 22708 8318
rect 22316 8306 22372 8316
rect 21980 7422 21982 7474
rect 22034 7422 22036 7474
rect 21980 7410 22036 7422
rect 22092 8258 22148 8270
rect 22092 8206 22094 8258
rect 22146 8206 22148 8258
rect 22092 7476 22148 8206
rect 22428 7586 22484 7598
rect 22428 7534 22430 7586
rect 22482 7534 22484 7586
rect 22204 7476 22260 7486
rect 22092 7420 22204 7476
rect 22204 7382 22260 7420
rect 22002 7084 22266 7094
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22002 7018 22266 7028
rect 21644 6860 21812 6916
rect 22092 6916 22148 6926
rect 21644 6244 21700 6860
rect 21868 6804 21924 6814
rect 21644 6188 21812 6244
rect 21532 5842 21588 5852
rect 21644 6020 21700 6030
rect 21644 5906 21700 5964
rect 21644 5854 21646 5906
rect 21698 5854 21700 5906
rect 21644 5842 21700 5854
rect 21756 5906 21812 6188
rect 21756 5854 21758 5906
rect 21810 5854 21812 5906
rect 19404 5796 19460 5806
rect 19740 5796 19796 5806
rect 19404 5794 19796 5796
rect 19404 5742 19406 5794
rect 19458 5742 19742 5794
rect 19794 5742 19796 5794
rect 19404 5740 19796 5742
rect 19404 5730 19460 5740
rect 19740 5730 19796 5740
rect 19852 5794 19908 5806
rect 19852 5742 19854 5794
rect 19906 5742 19908 5794
rect 19180 5236 19236 5246
rect 19180 5142 19236 5180
rect 19068 4470 19124 4508
rect 19516 5012 19572 5022
rect 19516 4340 19572 4956
rect 19516 4338 19796 4340
rect 19516 4286 19518 4338
rect 19570 4286 19796 4338
rect 19516 4284 19796 4286
rect 19516 4274 19572 4284
rect 19740 3556 19796 4284
rect 19740 3462 19796 3500
rect 19068 3442 19124 3454
rect 19068 3390 19070 3442
rect 19122 3390 19124 3442
rect 19068 3388 19124 3390
rect 19068 3332 19684 3388
rect 19852 3332 19908 5742
rect 21644 5236 21700 5246
rect 21644 5142 21700 5180
rect 21532 5010 21588 5022
rect 21532 4958 21534 5010
rect 21586 4958 21588 5010
rect 20300 4228 20356 4238
rect 20300 4134 20356 4172
rect 21532 3666 21588 4958
rect 21756 4340 21812 5854
rect 21868 5348 21924 6748
rect 22092 6690 22148 6860
rect 22092 6638 22094 6690
rect 22146 6638 22148 6690
rect 22092 6626 22148 6638
rect 22204 6802 22260 6814
rect 22204 6750 22206 6802
rect 22258 6750 22260 6802
rect 22204 6692 22260 6750
rect 22204 6626 22260 6636
rect 22316 6692 22372 6702
rect 22428 6692 22484 7534
rect 22316 6690 22484 6692
rect 22316 6638 22318 6690
rect 22370 6638 22484 6690
rect 22316 6636 22484 6638
rect 22316 6626 22372 6636
rect 22002 5516 22266 5526
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22002 5450 22266 5460
rect 21980 5348 22036 5358
rect 21868 5346 22036 5348
rect 21868 5294 21982 5346
rect 22034 5294 22036 5346
rect 21868 5292 22036 5294
rect 21980 5282 22036 5292
rect 21868 5122 21924 5134
rect 21868 5070 21870 5122
rect 21922 5070 21924 5122
rect 21868 4564 21924 5070
rect 21868 4498 21924 4508
rect 21756 4274 21812 4284
rect 22428 4226 22484 6636
rect 22540 7476 22596 7486
rect 22540 5794 22596 7420
rect 22652 5906 22708 8316
rect 23100 8258 23156 9660
rect 23100 8206 23102 8258
rect 23154 8206 23156 8258
rect 23100 8194 23156 8206
rect 23660 10052 23716 10062
rect 23324 8036 23380 8046
rect 23324 7586 23380 7980
rect 23324 7534 23326 7586
rect 23378 7534 23380 7586
rect 23324 7522 23380 7534
rect 23548 7586 23604 7598
rect 23548 7534 23550 7586
rect 23602 7534 23604 7586
rect 22652 5854 22654 5906
rect 22706 5854 22708 5906
rect 22652 5842 22708 5854
rect 22764 7474 22820 7486
rect 22764 7422 22766 7474
rect 22818 7422 22820 7474
rect 22540 5742 22542 5794
rect 22594 5742 22596 5794
rect 22540 5730 22596 5742
rect 22764 5122 22820 7422
rect 22988 7476 23044 7486
rect 22988 7382 23044 7420
rect 23436 7362 23492 7374
rect 23436 7310 23438 7362
rect 23490 7310 23492 7362
rect 23324 6916 23380 6926
rect 23212 6692 23268 6702
rect 23100 6690 23268 6692
rect 23100 6638 23214 6690
rect 23266 6638 23268 6690
rect 23100 6636 23268 6638
rect 22988 6580 23044 6590
rect 22988 6486 23044 6524
rect 22988 6020 23044 6030
rect 23100 6020 23156 6636
rect 23212 6626 23268 6636
rect 23044 5964 23156 6020
rect 22988 5926 23044 5964
rect 22764 5070 22766 5122
rect 22818 5070 22820 5122
rect 22764 5012 22820 5070
rect 22764 4946 22820 4956
rect 23324 5122 23380 6860
rect 23436 6804 23492 7310
rect 23548 6916 23604 7534
rect 23548 6850 23604 6860
rect 23436 6738 23492 6748
rect 23660 6692 23716 9996
rect 23772 8932 23828 8942
rect 23772 8370 23828 8876
rect 23772 8318 23774 8370
rect 23826 8318 23828 8370
rect 23772 8306 23828 8318
rect 23772 7252 23828 7262
rect 23884 7252 23940 10220
rect 24444 9716 24500 11342
rect 25228 11284 25284 11294
rect 25228 11282 25732 11284
rect 25228 11230 25230 11282
rect 25282 11230 25732 11282
rect 25228 11228 25732 11230
rect 25228 11218 25284 11228
rect 24444 9622 24500 9660
rect 24668 10836 24724 10846
rect 24668 9828 24724 10780
rect 25676 10498 25732 11228
rect 25788 10836 25844 14252
rect 26160 14140 26424 14150
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26160 14074 26424 14084
rect 26796 13860 26852 13870
rect 26124 13748 26180 13758
rect 26124 13654 26180 13692
rect 26348 13746 26404 13758
rect 26348 13694 26350 13746
rect 26402 13694 26404 13746
rect 26348 13412 26404 13694
rect 26684 13746 26740 13758
rect 26684 13694 26686 13746
rect 26738 13694 26740 13746
rect 26460 13636 26516 13646
rect 26460 13542 26516 13580
rect 26348 13076 26404 13356
rect 26348 13020 26628 13076
rect 26160 12572 26424 12582
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26160 12506 26424 12516
rect 26012 12178 26068 12190
rect 26012 12126 26014 12178
rect 26066 12126 26068 12178
rect 25788 10834 25956 10836
rect 25788 10782 25790 10834
rect 25842 10782 25956 10834
rect 25788 10780 25956 10782
rect 25788 10770 25844 10780
rect 25676 10446 25678 10498
rect 25730 10446 25732 10498
rect 25676 10434 25732 10446
rect 25900 10724 25956 10780
rect 23996 9268 24052 9278
rect 23996 9174 24052 9212
rect 24668 9266 24724 9772
rect 25900 9380 25956 10668
rect 26012 10722 26068 12126
rect 26572 12178 26628 13020
rect 26572 12126 26574 12178
rect 26626 12126 26628 12178
rect 26572 12114 26628 12126
rect 26684 12852 26740 13694
rect 26684 12066 26740 12796
rect 26684 12014 26686 12066
rect 26738 12014 26740 12066
rect 26684 12002 26740 12014
rect 26160 11004 26424 11014
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26160 10938 26424 10948
rect 26012 10670 26014 10722
rect 26066 10670 26068 10722
rect 26012 10658 26068 10670
rect 26796 9716 26852 13804
rect 27020 13860 27076 13870
rect 27020 13746 27076 13804
rect 27020 13694 27022 13746
rect 27074 13694 27076 13746
rect 27020 13682 27076 13694
rect 27356 13746 27412 15148
rect 27916 14756 27972 14766
rect 27804 14700 27916 14756
rect 27580 14530 27636 14542
rect 27580 14478 27582 14530
rect 27634 14478 27636 14530
rect 27356 13694 27358 13746
rect 27410 13694 27412 13746
rect 27356 13682 27412 13694
rect 27468 14418 27524 14430
rect 27468 14366 27470 14418
rect 27522 14366 27524 14418
rect 27468 13748 27524 14366
rect 27244 13636 27300 13646
rect 27244 13542 27300 13580
rect 26908 13524 26964 13534
rect 27468 13524 27524 13692
rect 26908 13430 26964 13468
rect 27356 13468 27524 13524
rect 26908 13076 26964 13086
rect 27356 13076 27412 13468
rect 26908 13074 27412 13076
rect 26908 13022 26910 13074
rect 26962 13022 27412 13074
rect 26908 13020 27412 13022
rect 26908 13010 26964 13020
rect 27356 12850 27412 13020
rect 27580 13412 27636 14478
rect 27804 14530 27860 14700
rect 27916 14690 27972 14700
rect 27804 14478 27806 14530
rect 27858 14478 27860 14530
rect 27804 14466 27860 14478
rect 27916 14532 27972 14542
rect 27804 13636 27860 13646
rect 27916 13636 27972 14476
rect 27804 13634 27972 13636
rect 27804 13582 27806 13634
rect 27858 13582 27972 13634
rect 27804 13580 27972 13582
rect 28028 13636 28084 15260
rect 28252 15204 28308 15932
rect 28364 15986 28420 16716
rect 28364 15934 28366 15986
rect 28418 15934 28420 15986
rect 28364 15922 28420 15934
rect 28924 15988 28980 17612
rect 29036 16212 29092 17724
rect 29148 17554 29204 17948
rect 29148 17502 29150 17554
rect 29202 17502 29204 17554
rect 29148 16660 29204 17502
rect 29260 16882 29316 18958
rect 29372 19012 29428 19022
rect 29372 18918 29428 18956
rect 29596 17892 29652 19180
rect 29708 18340 29764 19852
rect 29932 19842 29988 19852
rect 30318 19628 30582 19638
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30318 19562 30582 19572
rect 29820 19236 29876 19246
rect 29820 19234 30100 19236
rect 29820 19182 29822 19234
rect 29874 19182 30100 19234
rect 29820 19180 30100 19182
rect 29820 19170 29876 19180
rect 29708 18284 29876 18340
rect 29708 17892 29764 17902
rect 29484 17890 29764 17892
rect 29484 17838 29710 17890
rect 29762 17838 29764 17890
rect 29484 17836 29764 17838
rect 29372 17668 29428 17678
rect 29372 17574 29428 17612
rect 29372 16996 29428 17006
rect 29372 16902 29428 16940
rect 29260 16830 29262 16882
rect 29314 16830 29316 16882
rect 29260 16818 29316 16830
rect 29484 16884 29540 17836
rect 29708 17826 29764 17836
rect 29820 17668 29876 18284
rect 29596 17612 29876 17668
rect 29596 17106 29652 17612
rect 29596 17054 29598 17106
rect 29650 17054 29652 17106
rect 29596 17042 29652 17054
rect 30044 17108 30100 19180
rect 30716 18564 30772 19964
rect 34476 18844 34740 18854
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34476 18778 34740 18788
rect 30318 18060 30582 18070
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30318 17994 30582 18004
rect 30716 17780 30772 18508
rect 31948 17780 32004 17790
rect 30492 17724 31332 17780
rect 30492 17666 30548 17724
rect 30492 17614 30494 17666
rect 30546 17614 30548 17666
rect 30492 17602 30548 17614
rect 31164 17554 31220 17566
rect 31164 17502 31166 17554
rect 31218 17502 31220 17554
rect 30044 17106 30212 17108
rect 30044 17054 30046 17106
rect 30098 17054 30212 17106
rect 30044 17052 30212 17054
rect 30044 17042 30100 17052
rect 29708 16884 29764 16894
rect 29540 16882 29764 16884
rect 29540 16830 29710 16882
rect 29762 16830 29764 16882
rect 29540 16828 29764 16830
rect 29484 16790 29540 16828
rect 29708 16818 29764 16828
rect 29820 16772 29876 16782
rect 29148 16604 29428 16660
rect 29260 16212 29316 16222
rect 29036 16210 29316 16212
rect 29036 16158 29262 16210
rect 29314 16158 29316 16210
rect 29036 16156 29316 16158
rect 29260 16146 29316 16156
rect 29372 16100 29428 16604
rect 29372 16006 29428 16044
rect 29820 16098 29876 16716
rect 30156 16322 30212 17052
rect 30380 16994 30436 17006
rect 30380 16942 30382 16994
rect 30434 16942 30436 16994
rect 30380 16772 30436 16942
rect 30380 16706 30436 16716
rect 30318 16492 30582 16502
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30318 16426 30582 16436
rect 30156 16270 30158 16322
rect 30210 16270 30212 16322
rect 30156 16258 30212 16270
rect 29820 16046 29822 16098
rect 29874 16046 29876 16098
rect 29148 15988 29204 15998
rect 28980 15986 29204 15988
rect 28980 15934 29150 15986
rect 29202 15934 29204 15986
rect 28980 15932 29204 15934
rect 28924 15894 28980 15932
rect 29148 15922 29204 15932
rect 28476 15874 28532 15886
rect 28476 15822 28478 15874
rect 28530 15822 28532 15874
rect 28476 15540 28532 15822
rect 28252 14754 28308 15148
rect 28252 14702 28254 14754
rect 28306 14702 28308 14754
rect 28252 14690 28308 14702
rect 28364 15484 28532 15540
rect 27804 13570 27860 13580
rect 28028 13570 28084 13580
rect 27356 12798 27358 12850
rect 27410 12798 27412 12850
rect 27356 12786 27412 12798
rect 27468 12964 27524 12974
rect 27580 12964 27636 13356
rect 28364 13188 28420 15484
rect 28812 15316 28868 15326
rect 28700 15260 28812 15316
rect 28252 13132 28420 13188
rect 28476 15090 28532 15102
rect 28476 15038 28478 15090
rect 28530 15038 28532 15090
rect 28476 14756 28532 15038
rect 27468 12962 27636 12964
rect 27468 12910 27470 12962
rect 27522 12910 27636 12962
rect 27468 12908 27636 12910
rect 28028 12964 28084 12974
rect 27132 12740 27188 12750
rect 26908 12738 27188 12740
rect 26908 12686 27134 12738
rect 27186 12686 27188 12738
rect 26908 12684 27188 12686
rect 26908 10052 26964 12684
rect 27132 12674 27188 12684
rect 27356 11508 27412 11518
rect 27468 11508 27524 12908
rect 28028 12870 28084 12908
rect 27356 11506 27524 11508
rect 27356 11454 27358 11506
rect 27410 11454 27524 11506
rect 27356 11452 27524 11454
rect 27356 11442 27412 11452
rect 28252 11172 28308 13132
rect 28364 12964 28420 12974
rect 28476 12964 28532 14700
rect 28700 14532 28756 15260
rect 28812 15222 28868 15260
rect 28588 14476 28700 14532
rect 28588 13074 28644 14476
rect 28700 14466 28756 14476
rect 28812 15090 28868 15102
rect 28812 15038 28814 15090
rect 28866 15038 28868 15090
rect 28588 13022 28590 13074
rect 28642 13022 28644 13074
rect 28588 13010 28644 13022
rect 28364 12962 28532 12964
rect 28364 12910 28366 12962
rect 28418 12910 28532 12962
rect 28364 12908 28532 12910
rect 28812 12964 28868 15038
rect 29148 14420 29204 14430
rect 29148 14326 29204 14364
rect 29484 14308 29540 14318
rect 29484 14306 29652 14308
rect 29484 14254 29486 14306
rect 29538 14254 29652 14306
rect 29484 14252 29652 14254
rect 29484 14242 29540 14252
rect 29596 13188 29652 14252
rect 29820 13860 29876 16046
rect 30044 15986 30100 15998
rect 30044 15934 30046 15986
rect 30098 15934 30100 15986
rect 30044 14420 30100 15934
rect 31164 15764 31220 17502
rect 31276 16098 31332 17724
rect 31948 17108 32004 17724
rect 33292 17780 33348 17790
rect 33292 17686 33348 17724
rect 34476 17276 34740 17286
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34476 17210 34740 17220
rect 31724 17106 32004 17108
rect 31724 17054 31950 17106
rect 32002 17054 32004 17106
rect 31724 17052 32004 17054
rect 31500 16882 31556 16894
rect 31500 16830 31502 16882
rect 31554 16830 31556 16882
rect 31500 16772 31556 16830
rect 31500 16706 31556 16716
rect 31276 16046 31278 16098
rect 31330 16046 31332 16098
rect 31276 16034 31332 16046
rect 31164 15698 31220 15708
rect 30380 15540 30436 15550
rect 30380 15446 30436 15484
rect 30940 15428 30996 15438
rect 30940 15334 30996 15372
rect 31388 15428 31444 15438
rect 31052 15316 31108 15326
rect 31388 15316 31444 15372
rect 31052 15314 31444 15316
rect 31052 15262 31054 15314
rect 31106 15262 31444 15314
rect 31052 15260 31444 15262
rect 31052 15250 31108 15260
rect 30492 15202 30548 15214
rect 30492 15150 30494 15202
rect 30546 15150 30548 15202
rect 30492 15092 30548 15150
rect 30604 15204 30660 15242
rect 30604 15138 30660 15148
rect 31276 15092 31332 15102
rect 30492 15026 30548 15036
rect 30828 15090 31332 15092
rect 30828 15038 31278 15090
rect 31330 15038 31332 15090
rect 30828 15036 31332 15038
rect 30318 14924 30582 14934
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30318 14858 30582 14868
rect 30828 14754 30884 15036
rect 31276 15026 31332 15036
rect 31388 14756 31444 15260
rect 31500 15316 31556 15326
rect 31500 15222 31556 15260
rect 31724 15314 31780 17052
rect 31948 17042 32004 17052
rect 32172 16884 32228 16894
rect 32172 16882 32900 16884
rect 32172 16830 32174 16882
rect 32226 16830 32900 16882
rect 32172 16828 32900 16830
rect 32172 16818 32228 16828
rect 32060 16772 32116 16782
rect 31948 16770 32116 16772
rect 31948 16718 32062 16770
rect 32114 16718 32116 16770
rect 31948 16716 32116 16718
rect 31948 15428 32004 16716
rect 32060 16706 32116 16716
rect 32060 15988 32116 15998
rect 32060 15986 32788 15988
rect 32060 15934 32062 15986
rect 32114 15934 32788 15986
rect 32060 15932 32788 15934
rect 32060 15922 32116 15932
rect 32284 15764 32340 15774
rect 32340 15708 32452 15764
rect 32284 15698 32340 15708
rect 32060 15428 32116 15438
rect 31948 15426 32116 15428
rect 31948 15374 32062 15426
rect 32114 15374 32116 15426
rect 31948 15372 32116 15374
rect 32060 15362 32116 15372
rect 32284 15426 32340 15438
rect 32284 15374 32286 15426
rect 32338 15374 32340 15426
rect 31724 15262 31726 15314
rect 31778 15262 31780 15314
rect 31724 15148 31780 15262
rect 30828 14702 30830 14754
rect 30882 14702 30884 14754
rect 30828 14690 30884 14702
rect 31164 14700 31444 14756
rect 31612 15092 31780 15148
rect 31164 14530 31220 14700
rect 31164 14478 31166 14530
rect 31218 14478 31220 14530
rect 31164 14466 31220 14478
rect 31276 14530 31332 14542
rect 31276 14478 31278 14530
rect 31330 14478 31332 14530
rect 30044 14354 30100 14364
rect 30716 14418 30772 14430
rect 30716 14366 30718 14418
rect 30770 14366 30772 14418
rect 30716 14308 30772 14366
rect 31276 14308 31332 14478
rect 31612 14530 31668 15092
rect 32172 14756 32228 14766
rect 32284 14756 32340 15374
rect 32396 15202 32452 15708
rect 32396 15150 32398 15202
rect 32450 15150 32452 15202
rect 32396 15138 32452 15150
rect 32508 15204 32564 15214
rect 32732 15148 32788 15932
rect 32228 14700 32340 14756
rect 32172 14662 32228 14700
rect 31612 14478 31614 14530
rect 31666 14478 31668 14530
rect 31612 14466 31668 14478
rect 31836 14530 31892 14542
rect 31836 14478 31838 14530
rect 31890 14478 31892 14530
rect 30716 14252 31780 14308
rect 31164 13970 31220 14252
rect 31164 13918 31166 13970
rect 31218 13918 31220 13970
rect 29820 13804 30100 13860
rect 29932 13636 29988 13646
rect 29596 13094 29652 13132
rect 29708 13634 29988 13636
rect 29708 13582 29934 13634
rect 29986 13582 29988 13634
rect 29708 13580 29988 13582
rect 29708 13186 29764 13580
rect 29932 13570 29988 13580
rect 29708 13134 29710 13186
rect 29762 13134 29764 13186
rect 29708 13122 29764 13134
rect 29148 12964 29204 12974
rect 28812 12962 29204 12964
rect 28812 12910 29150 12962
rect 29202 12910 29204 12962
rect 28812 12908 29204 12910
rect 28364 12898 28420 12908
rect 29148 12898 29204 12908
rect 29372 12964 29428 12974
rect 29372 12870 29428 12908
rect 29820 11396 29876 11406
rect 30044 11396 30100 13804
rect 30716 13746 30772 13758
rect 30716 13694 30718 13746
rect 30770 13694 30772 13746
rect 30318 13356 30582 13366
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30318 13290 30582 13300
rect 30318 11788 30582 11798
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30318 11722 30582 11732
rect 29820 11394 30100 11396
rect 29820 11342 29822 11394
rect 29874 11342 30100 11394
rect 29820 11340 30100 11342
rect 30268 11394 30324 11406
rect 30268 11342 30270 11394
rect 30322 11342 30324 11394
rect 28252 11116 28420 11172
rect 26908 9986 26964 9996
rect 27132 10610 27188 10622
rect 27132 10558 27134 10610
rect 27186 10558 27188 10610
rect 27132 10052 27188 10558
rect 27132 9986 27188 9996
rect 27804 10498 27860 10510
rect 27804 10446 27806 10498
rect 27858 10446 27860 10498
rect 27804 9940 27860 10446
rect 27804 9874 27860 9884
rect 26572 9660 26796 9716
rect 26160 9436 26424 9446
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 24668 9214 24670 9266
rect 24722 9214 24724 9266
rect 24668 9202 24724 9214
rect 25564 9324 26068 9380
rect 26160 9370 26424 9380
rect 25564 9042 25620 9324
rect 26012 9268 26068 9324
rect 26236 9268 26292 9278
rect 26012 9266 26292 9268
rect 26012 9214 26238 9266
rect 26290 9214 26292 9266
rect 26012 9212 26292 9214
rect 26236 9202 26292 9212
rect 26572 9266 26628 9660
rect 26796 9650 26852 9660
rect 27244 9828 27300 9838
rect 26572 9214 26574 9266
rect 26626 9214 26628 9266
rect 26572 9202 26628 9214
rect 25564 8990 25566 9042
rect 25618 8990 25620 9042
rect 25564 8978 25620 8990
rect 27244 9042 27300 9772
rect 27244 8990 27246 9042
rect 27298 8990 27300 9042
rect 27244 8978 27300 8990
rect 27916 9604 27972 9614
rect 28140 9604 28196 9614
rect 27972 9602 28196 9604
rect 27972 9550 28142 9602
rect 28194 9550 28196 9602
rect 27972 9548 28196 9550
rect 25340 8932 25396 8942
rect 25340 8838 25396 8876
rect 25228 8818 25284 8830
rect 25228 8766 25230 8818
rect 25282 8766 25284 8818
rect 23828 7196 23940 7252
rect 24108 7252 24164 7262
rect 25228 7252 25284 8766
rect 25900 8370 25956 8382
rect 25900 8318 25902 8370
rect 25954 8318 25956 8370
rect 25900 8260 25956 8318
rect 25900 7586 25956 8204
rect 26908 8260 26964 8270
rect 27692 8260 27748 8270
rect 26908 8166 26964 8204
rect 27580 8258 27748 8260
rect 27580 8206 27694 8258
rect 27746 8206 27748 8258
rect 27580 8204 27748 8206
rect 26236 8036 26292 8046
rect 26012 8034 26292 8036
rect 26012 7982 26238 8034
rect 26290 7982 26292 8034
rect 26012 7980 26292 7982
rect 26012 7700 26068 7980
rect 26236 7970 26292 7980
rect 26572 8034 26628 8046
rect 26572 7982 26574 8034
rect 26626 7982 26628 8034
rect 26160 7868 26424 7878
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26160 7802 26424 7812
rect 26012 7644 26292 7700
rect 25900 7534 25902 7586
rect 25954 7534 25956 7586
rect 25900 7522 25956 7534
rect 25564 7476 25620 7486
rect 23772 6802 23828 7196
rect 23772 6750 23774 6802
rect 23826 6750 23828 6802
rect 23772 6738 23828 6750
rect 23660 6626 23716 6636
rect 24108 6578 24164 7196
rect 25116 7196 25284 7252
rect 25340 7474 25620 7476
rect 25340 7422 25566 7474
rect 25618 7422 25620 7474
rect 25340 7420 25620 7422
rect 24108 6526 24110 6578
rect 24162 6526 24164 6578
rect 24108 6514 24164 6526
rect 24780 6580 24836 6590
rect 24780 6486 24836 6524
rect 24220 6020 24276 6030
rect 24108 5908 24164 5918
rect 23324 5070 23326 5122
rect 23378 5070 23380 5122
rect 22428 4174 22430 4226
rect 22482 4174 22484 4226
rect 22002 3948 22266 3958
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22002 3882 22266 3892
rect 21532 3614 21534 3666
rect 21586 3614 21588 3666
rect 21532 3602 21588 3614
rect 20748 3556 20804 3566
rect 20748 3462 20804 3500
rect 22428 3556 22484 4174
rect 22764 4564 22820 4574
rect 22764 3668 22820 4508
rect 23100 4340 23156 4350
rect 23100 4246 23156 4284
rect 23324 4226 23380 5070
rect 23772 5236 23828 5246
rect 23436 5012 23492 5022
rect 23492 4956 23604 5012
rect 23436 4946 23492 4956
rect 23324 4174 23326 4226
rect 23378 4174 23380 4226
rect 23324 4116 23380 4174
rect 23324 4050 23380 4060
rect 23548 3668 23604 4956
rect 23772 4338 23828 5180
rect 24108 5234 24164 5852
rect 24220 5906 24276 5964
rect 24668 6020 24724 6030
rect 25116 6020 25172 7196
rect 24668 6018 25172 6020
rect 24668 5966 24670 6018
rect 24722 5966 25172 6018
rect 24668 5964 25172 5966
rect 25340 6580 25396 7420
rect 25564 7410 25620 7420
rect 26012 7474 26068 7486
rect 26012 7422 26014 7474
rect 26066 7422 26068 7474
rect 24668 5954 24724 5964
rect 24220 5854 24222 5906
rect 24274 5854 24276 5906
rect 24220 5842 24276 5854
rect 25228 5908 25284 5918
rect 25340 5908 25396 6524
rect 26012 6916 26068 7422
rect 26236 7476 26292 7644
rect 26572 7476 26628 7982
rect 27244 8034 27300 8046
rect 27244 7982 27246 8034
rect 27298 7982 27300 8034
rect 27244 7476 27300 7982
rect 27580 7698 27636 8204
rect 27692 8194 27748 8204
rect 27580 7646 27582 7698
rect 27634 7646 27636 7698
rect 27580 7634 27636 7646
rect 27468 7476 27524 7486
rect 26572 7420 26852 7476
rect 26236 7382 26292 7420
rect 26012 6244 26068 6860
rect 26684 7250 26740 7262
rect 26684 7198 26686 7250
rect 26738 7198 26740 7250
rect 26684 6804 26740 7198
rect 26460 6692 26516 6702
rect 26460 6598 26516 6636
rect 25900 6188 26068 6244
rect 26160 6300 26424 6310
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26160 6234 26424 6244
rect 25452 6020 25508 6030
rect 25452 5926 25508 5964
rect 25284 5852 25396 5908
rect 25564 5906 25620 5918
rect 25564 5854 25566 5906
rect 25618 5854 25620 5906
rect 25228 5814 25284 5852
rect 24108 5182 24110 5234
rect 24162 5182 24164 5234
rect 24108 5170 24164 5182
rect 24332 5796 24388 5806
rect 23772 4286 23774 4338
rect 23826 4286 23828 4338
rect 23772 4274 23828 4286
rect 24220 4340 24276 4350
rect 24332 4340 24388 5740
rect 25564 5796 25620 5854
rect 25564 5730 25620 5740
rect 24220 4338 24388 4340
rect 24220 4286 24222 4338
rect 24274 4286 24388 4338
rect 24220 4284 24388 4286
rect 24220 4274 24276 4284
rect 23660 4228 23716 4238
rect 23660 4134 23716 4172
rect 25788 4228 25844 4238
rect 25900 4228 25956 6188
rect 26684 5906 26740 6748
rect 26684 5854 26686 5906
rect 26738 5854 26740 5906
rect 26684 5842 26740 5854
rect 26796 6578 26852 7420
rect 27132 7474 27524 7476
rect 27132 7422 27470 7474
rect 27522 7422 27524 7474
rect 27132 7420 27524 7422
rect 27020 6692 27076 6702
rect 27132 6692 27188 7420
rect 27468 7410 27524 7420
rect 27692 7474 27748 7486
rect 27692 7422 27694 7474
rect 27746 7422 27748 7474
rect 27692 7364 27748 7422
rect 27692 7298 27748 7308
rect 26796 6526 26798 6578
rect 26850 6526 26852 6578
rect 26796 5908 26852 6526
rect 26908 6690 27188 6692
rect 26908 6638 27022 6690
rect 27074 6638 27188 6690
rect 26908 6636 27188 6638
rect 27244 7250 27300 7262
rect 27244 7198 27246 7250
rect 27298 7198 27300 7250
rect 27244 6690 27300 7198
rect 27692 7140 27748 7150
rect 27244 6638 27246 6690
rect 27298 6638 27300 6690
rect 26908 6020 26964 6636
rect 27020 6626 27076 6636
rect 27244 6580 27300 6638
rect 27244 6514 27300 6524
rect 27580 7084 27692 7140
rect 26908 5954 26964 5964
rect 27020 6466 27076 6478
rect 27020 6414 27022 6466
rect 27074 6414 27076 6466
rect 27020 5908 27076 6414
rect 27580 6132 27636 7084
rect 27692 7074 27748 7084
rect 27916 6690 27972 9548
rect 28140 9538 28196 9548
rect 28140 8370 28196 8382
rect 28140 8318 28142 8370
rect 28194 8318 28196 8370
rect 28028 8148 28084 8158
rect 28028 8054 28084 8092
rect 28140 7698 28196 8318
rect 28140 7646 28142 7698
rect 28194 7646 28196 7698
rect 28140 7634 28196 7646
rect 28252 8034 28308 8046
rect 28252 7982 28254 8034
rect 28306 7982 28308 8034
rect 28028 7252 28084 7262
rect 28028 7158 28084 7196
rect 28252 7140 28308 7982
rect 28364 7586 28420 11116
rect 29148 11170 29204 11182
rect 29148 11118 29150 11170
rect 29202 11118 29204 11170
rect 29148 9828 29204 11118
rect 29148 9762 29204 9772
rect 29260 11170 29316 11182
rect 29260 11118 29262 11170
rect 29314 11118 29316 11170
rect 29260 9826 29316 11118
rect 29260 9774 29262 9826
rect 29314 9774 29316 9826
rect 29260 9762 29316 9774
rect 29372 11170 29428 11182
rect 29372 11118 29374 11170
rect 29426 11118 29428 11170
rect 29372 9716 29428 11118
rect 29372 9622 29428 9660
rect 29484 9940 29540 9950
rect 28476 9604 28532 9614
rect 28476 9510 28532 9548
rect 29260 9604 29316 9614
rect 28364 7534 28366 7586
rect 28418 7534 28420 7586
rect 28364 7522 28420 7534
rect 28252 7074 28308 7084
rect 29148 7474 29204 7486
rect 29148 7422 29150 7474
rect 29202 7422 29204 7474
rect 29148 7364 29204 7422
rect 27916 6638 27918 6690
rect 27970 6638 27972 6690
rect 27916 6626 27972 6638
rect 28700 6804 28756 6814
rect 27692 6468 27748 6478
rect 27692 6466 27860 6468
rect 27692 6414 27694 6466
rect 27746 6414 27860 6466
rect 27692 6412 27860 6414
rect 27692 6402 27748 6412
rect 27692 6132 27748 6142
rect 27580 6130 27748 6132
rect 27580 6078 27694 6130
rect 27746 6078 27748 6130
rect 27580 6076 27748 6078
rect 27692 6066 27748 6076
rect 27468 5908 27524 5918
rect 27020 5852 27412 5908
rect 26796 5842 26852 5852
rect 26012 5796 26068 5806
rect 26012 5702 26068 5740
rect 26796 5684 26852 5694
rect 27020 5684 27076 5694
rect 26796 5590 26852 5628
rect 26908 5682 27076 5684
rect 26908 5630 27022 5682
rect 27074 5630 27076 5682
rect 26908 5628 27076 5630
rect 26908 5236 26964 5628
rect 27020 5618 27076 5628
rect 27132 5684 27188 5694
rect 27132 5682 27300 5684
rect 27132 5630 27134 5682
rect 27186 5630 27300 5682
rect 27132 5628 27300 5630
rect 27132 5618 27188 5628
rect 26908 5170 26964 5180
rect 27020 5124 27076 5134
rect 27020 5030 27076 5068
rect 26236 5012 26292 5022
rect 26236 4918 26292 4956
rect 26160 4732 26424 4742
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26160 4666 26424 4676
rect 27244 4676 27300 5628
rect 27356 5122 27412 5852
rect 27468 5348 27524 5852
rect 27580 5796 27636 5806
rect 27580 5702 27636 5740
rect 27580 5348 27636 5358
rect 27468 5346 27636 5348
rect 27468 5294 27582 5346
rect 27634 5294 27636 5346
rect 27468 5292 27636 5294
rect 27580 5282 27636 5292
rect 27804 5236 27860 6412
rect 28700 6018 28756 6748
rect 29148 6690 29204 7308
rect 29148 6638 29150 6690
rect 29202 6638 29204 6690
rect 28700 5966 28702 6018
rect 28754 5966 28756 6018
rect 28700 5954 28756 5966
rect 28924 6020 28980 6030
rect 29148 6020 29204 6638
rect 28924 6018 29204 6020
rect 28924 5966 28926 6018
rect 28978 5966 29204 6018
rect 28924 5964 29204 5966
rect 29260 7252 29316 9548
rect 29484 9602 29540 9884
rect 29484 9550 29486 9602
rect 29538 9550 29540 9602
rect 29484 9538 29540 9550
rect 29708 9828 29764 9838
rect 29708 8484 29764 9772
rect 29708 8418 29764 8428
rect 29484 8258 29540 8270
rect 29484 8206 29486 8258
rect 29538 8206 29540 8258
rect 29372 8148 29428 8158
rect 29372 8054 29428 8092
rect 29484 7588 29540 8206
rect 29708 8260 29764 8270
rect 29708 8166 29764 8204
rect 29820 8036 29876 11340
rect 30044 11170 30100 11182
rect 30044 11118 30046 11170
rect 30098 11118 30100 11170
rect 29932 10500 29988 10510
rect 29932 10406 29988 10444
rect 29932 10276 29988 10286
rect 29932 9828 29988 10220
rect 29932 8482 29988 9772
rect 30044 9716 30100 11118
rect 30268 10500 30324 11342
rect 30380 10612 30436 10622
rect 30380 10518 30436 10556
rect 30492 10610 30548 10622
rect 30492 10558 30494 10610
rect 30546 10558 30548 10610
rect 30268 10434 30324 10444
rect 30492 10388 30548 10558
rect 30492 10322 30548 10332
rect 30318 10220 30582 10230
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30318 10154 30582 10164
rect 30716 10052 30772 13694
rect 31164 13076 31220 13918
rect 31724 13746 31780 14252
rect 31724 13694 31726 13746
rect 31778 13694 31780 13746
rect 31724 13682 31780 13694
rect 31276 13634 31332 13646
rect 31276 13582 31278 13634
rect 31330 13582 31332 13634
rect 31276 13524 31332 13582
rect 31276 13458 31332 13468
rect 31388 13524 31444 13534
rect 31836 13524 31892 14478
rect 32060 14532 32116 14542
rect 31948 13524 32004 13534
rect 31388 13522 32004 13524
rect 31388 13470 31390 13522
rect 31442 13470 31950 13522
rect 32002 13470 32004 13522
rect 31388 13468 32004 13470
rect 31388 13458 31444 13468
rect 31276 13076 31332 13086
rect 31164 13074 31332 13076
rect 31164 13022 31278 13074
rect 31330 13022 31332 13074
rect 31164 13020 31332 13022
rect 31276 13010 31332 13020
rect 31388 12180 31444 12190
rect 31052 12178 31444 12180
rect 31052 12126 31390 12178
rect 31442 12126 31444 12178
rect 31052 12124 31444 12126
rect 30940 10724 30996 10734
rect 30828 10610 30884 10622
rect 30828 10558 30830 10610
rect 30882 10558 30884 10610
rect 30828 10500 30884 10558
rect 30940 10610 30996 10668
rect 30940 10558 30942 10610
rect 30994 10558 30996 10610
rect 30940 10546 30996 10558
rect 30828 10434 30884 10444
rect 31052 10276 31108 12124
rect 31388 12114 31444 12124
rect 31500 11956 31556 13468
rect 31948 13458 32004 13468
rect 32060 13300 32116 14476
rect 32284 13972 32340 13982
rect 32508 13972 32564 15148
rect 32620 15092 32788 15148
rect 32844 15540 32900 16828
rect 34188 16212 34244 16222
rect 33628 16210 34244 16212
rect 33628 16158 34190 16210
rect 34242 16158 34244 16210
rect 33628 16156 34244 16158
rect 33068 15540 33124 15550
rect 32844 15538 33124 15540
rect 32844 15486 33070 15538
rect 33122 15486 33124 15538
rect 32844 15484 33124 15486
rect 32620 14308 32676 15092
rect 32732 14980 32788 14990
rect 32732 14754 32788 14924
rect 32732 14702 32734 14754
rect 32786 14702 32788 14754
rect 32732 14690 32788 14702
rect 32844 14754 32900 15484
rect 33068 15474 33124 15484
rect 33628 15428 33684 16156
rect 34188 16146 34244 16156
rect 34476 15708 34740 15718
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34476 15642 34740 15652
rect 33628 15314 33684 15372
rect 33628 15262 33630 15314
rect 33682 15262 33684 15314
rect 33628 15250 33684 15262
rect 32844 14702 32846 14754
rect 32898 14702 32900 14754
rect 32844 14690 32900 14702
rect 33180 15204 33236 15214
rect 33404 15204 33460 15214
rect 33236 15202 33460 15204
rect 33236 15150 33406 15202
rect 33458 15150 33460 15202
rect 33236 15148 33460 15150
rect 33068 14532 33124 14542
rect 32732 14308 32788 14318
rect 32620 14306 32788 14308
rect 32620 14254 32734 14306
rect 32786 14254 32788 14306
rect 32620 14252 32788 14254
rect 32732 14242 32788 14252
rect 32284 13970 32564 13972
rect 32284 13918 32286 13970
rect 32338 13918 32564 13970
rect 32284 13916 32564 13918
rect 32284 13906 32340 13916
rect 31836 13244 32116 13300
rect 32396 13636 32452 13646
rect 31836 13188 31892 13244
rect 31836 12178 31892 13132
rect 31836 12126 31838 12178
rect 31890 12126 31892 12178
rect 31836 12114 31892 12126
rect 31612 11956 31668 11966
rect 31500 11954 31668 11956
rect 31500 11902 31614 11954
rect 31666 11902 31668 11954
rect 31500 11900 31668 11902
rect 31276 11508 31332 11518
rect 31164 11506 31332 11508
rect 31164 11454 31278 11506
rect 31330 11454 31332 11506
rect 31164 11452 31332 11454
rect 31164 10388 31220 11452
rect 31276 11442 31332 11452
rect 31388 10836 31444 10846
rect 31612 10836 31668 11900
rect 31948 11956 32004 11966
rect 31948 11862 32004 11900
rect 31388 10834 31668 10836
rect 31388 10782 31390 10834
rect 31442 10782 31668 10834
rect 31388 10780 31668 10782
rect 31388 10770 31444 10780
rect 31836 10724 31892 10734
rect 31724 10668 31836 10724
rect 31164 10322 31220 10332
rect 31276 10612 31332 10622
rect 30380 9828 30436 9838
rect 30380 9734 30436 9772
rect 30156 9716 30212 9726
rect 30044 9660 30156 9716
rect 29932 8430 29934 8482
rect 29986 8430 29988 8482
rect 29932 8418 29988 8430
rect 30156 9492 30212 9660
rect 30604 9714 30660 9726
rect 30604 9662 30606 9714
rect 30658 9662 30660 9714
rect 30604 9492 30660 9662
rect 30156 9436 30660 9492
rect 30156 8258 30212 9436
rect 30716 9156 30772 9996
rect 30828 10220 31108 10276
rect 30828 9938 30884 10220
rect 30828 9886 30830 9938
rect 30882 9886 30884 9938
rect 30828 9874 30884 9886
rect 30940 9940 30996 9950
rect 30940 9826 30996 9884
rect 30940 9774 30942 9826
rect 30994 9774 30996 9826
rect 30940 9762 30996 9774
rect 31276 9938 31332 10556
rect 31276 9886 31278 9938
rect 31330 9886 31332 9938
rect 31276 9380 31332 9886
rect 30716 9090 30772 9100
rect 31164 9324 31332 9380
rect 30318 8652 30582 8662
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30318 8586 30582 8596
rect 30156 8206 30158 8258
rect 30210 8206 30212 8258
rect 30156 8194 30212 8206
rect 30380 8484 30436 8494
rect 30380 8036 30436 8428
rect 30604 8372 30660 8382
rect 31164 8372 31220 9324
rect 30604 8370 31220 8372
rect 30604 8318 30606 8370
rect 30658 8318 31220 8370
rect 30604 8316 31220 8318
rect 31388 9156 31444 9166
rect 30604 8306 30660 8316
rect 30492 8260 30548 8270
rect 30492 8166 30548 8204
rect 31052 8036 31108 8316
rect 31388 8258 31444 9100
rect 31388 8206 31390 8258
rect 31442 8206 31444 8258
rect 29820 7980 30212 8036
rect 30380 7980 30772 8036
rect 31052 7980 31332 8036
rect 29484 7494 29540 7532
rect 29708 7644 29988 7700
rect 29708 7586 29764 7644
rect 29708 7534 29710 7586
rect 29762 7534 29764 7586
rect 29708 7522 29764 7534
rect 27804 5142 27860 5180
rect 27356 5070 27358 5122
rect 27410 5070 27412 5122
rect 27356 5058 27412 5070
rect 28700 5012 28756 5022
rect 27468 4900 27524 4910
rect 27468 4806 27524 4844
rect 27244 4620 27972 4676
rect 27916 4450 27972 4620
rect 27916 4398 27918 4450
rect 27970 4398 27972 4450
rect 27916 4386 27972 4398
rect 28700 4338 28756 4956
rect 28700 4286 28702 4338
rect 28754 4286 28756 4338
rect 28700 4274 28756 4286
rect 25788 4226 25956 4228
rect 25788 4174 25790 4226
rect 25842 4174 25956 4226
rect 25788 4172 25956 4174
rect 28924 4228 28980 5964
rect 29036 5682 29092 5694
rect 29036 5630 29038 5682
rect 29090 5630 29092 5682
rect 29036 5124 29092 5630
rect 29260 5346 29316 7196
rect 29820 7474 29876 7486
rect 29820 7422 29822 7474
rect 29874 7422 29876 7474
rect 29820 7028 29876 7422
rect 29596 6972 29876 7028
rect 29372 6804 29428 6814
rect 29596 6804 29652 6972
rect 29428 6748 29652 6804
rect 29708 6804 29764 6814
rect 29372 6710 29428 6748
rect 29708 6710 29764 6748
rect 29932 6692 29988 7644
rect 30156 6916 30212 7980
rect 30716 7698 30772 7980
rect 30716 7646 30718 7698
rect 30770 7646 30772 7698
rect 30716 7634 30772 7646
rect 30268 7476 30324 7486
rect 30268 7382 30324 7420
rect 31052 7476 31108 7486
rect 31052 7382 31108 7420
rect 31276 7474 31332 7980
rect 31276 7422 31278 7474
rect 31330 7422 31332 7474
rect 31276 7410 31332 7422
rect 30318 7084 30582 7094
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30318 7018 30582 7028
rect 30716 6916 30772 6926
rect 30156 6860 30324 6916
rect 29932 6244 29988 6636
rect 29932 6178 29988 6188
rect 30044 6804 30100 6814
rect 29820 6018 29876 6030
rect 29820 5966 29822 6018
rect 29874 5966 29876 6018
rect 29820 5908 29876 5966
rect 29260 5294 29262 5346
rect 29314 5294 29316 5346
rect 29260 5282 29316 5294
rect 29708 5852 29820 5908
rect 29484 5124 29540 5134
rect 29036 5122 29540 5124
rect 29036 5070 29486 5122
rect 29538 5070 29540 5122
rect 29036 5068 29540 5070
rect 29484 5058 29540 5068
rect 29708 5124 29764 5852
rect 29820 5842 29876 5852
rect 30044 5906 30100 6748
rect 30156 6690 30212 6702
rect 30156 6638 30158 6690
rect 30210 6638 30212 6690
rect 30156 6244 30212 6638
rect 30156 6178 30212 6188
rect 30044 5854 30046 5906
rect 30098 5854 30100 5906
rect 30044 5842 30100 5854
rect 30268 5908 30324 6860
rect 30380 6804 30436 6814
rect 30380 6710 30436 6748
rect 30716 6690 30772 6860
rect 30716 6638 30718 6690
rect 30770 6638 30772 6690
rect 30716 6626 30772 6638
rect 31164 6692 31220 6702
rect 31388 6692 31444 8206
rect 31724 7476 31780 10668
rect 31836 10630 31892 10668
rect 32172 10612 32228 10650
rect 32172 10546 32228 10556
rect 32172 10386 32228 10398
rect 32172 10334 32174 10386
rect 32226 10334 32228 10386
rect 31836 9156 31892 9166
rect 31836 9062 31892 9100
rect 32172 9044 32228 10334
rect 32172 8978 32228 8988
rect 32060 8146 32116 8158
rect 32060 8094 32062 8146
rect 32114 8094 32116 8146
rect 32060 7698 32116 8094
rect 32060 7646 32062 7698
rect 32114 7646 32116 7698
rect 32060 7634 32116 7646
rect 32172 7586 32228 7598
rect 32172 7534 32174 7586
rect 32226 7534 32228 7586
rect 31948 7476 32004 7486
rect 31780 7474 32004 7476
rect 31780 7422 31950 7474
rect 32002 7422 32004 7474
rect 31780 7420 32004 7422
rect 31724 7410 31780 7420
rect 31948 7410 32004 7420
rect 32172 7474 32228 7534
rect 32172 7422 32174 7474
rect 32226 7422 32228 7474
rect 32172 7410 32228 7422
rect 31724 7252 31780 7262
rect 31780 7196 32004 7252
rect 31724 7158 31780 7196
rect 31164 6690 31444 6692
rect 31164 6638 31166 6690
rect 31218 6638 31444 6690
rect 31164 6636 31444 6638
rect 31612 6916 31668 6926
rect 31164 6626 31220 6636
rect 30940 6020 30996 6030
rect 30716 5964 30940 6020
rect 30492 5908 30548 5918
rect 30268 5906 30548 5908
rect 30268 5854 30494 5906
rect 30546 5854 30548 5906
rect 30268 5852 30548 5854
rect 30492 5842 30548 5852
rect 30318 5516 30582 5526
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30318 5450 30582 5460
rect 30604 5236 30660 5246
rect 30492 5180 30604 5236
rect 29708 5030 29764 5068
rect 30380 5124 30436 5134
rect 30380 5030 30436 5068
rect 30492 5122 30548 5180
rect 30604 5170 30660 5180
rect 30492 5070 30494 5122
rect 30546 5070 30548 5122
rect 30492 5058 30548 5070
rect 30716 5122 30772 5964
rect 30940 5926 30996 5964
rect 31164 5908 31220 5918
rect 31164 5814 31220 5852
rect 31052 5794 31108 5806
rect 31052 5742 31054 5794
rect 31106 5742 31108 5794
rect 30716 5070 30718 5122
rect 30770 5070 30772 5122
rect 30716 5058 30772 5070
rect 30940 5124 30996 5134
rect 31052 5124 31108 5742
rect 30940 5122 31108 5124
rect 30940 5070 30942 5122
rect 30994 5070 31108 5122
rect 30940 5068 31108 5070
rect 31276 5122 31332 6636
rect 31612 5906 31668 6860
rect 31612 5854 31614 5906
rect 31666 5854 31668 5906
rect 31612 5842 31668 5854
rect 31836 6578 31892 6590
rect 31836 6526 31838 6578
rect 31890 6526 31892 6578
rect 31724 5796 31780 5806
rect 31724 5702 31780 5740
rect 31836 5236 31892 6526
rect 31948 5906 32004 7196
rect 31948 5854 31950 5906
rect 32002 5854 32004 5906
rect 31948 5842 32004 5854
rect 31836 5170 31892 5180
rect 32060 5682 32116 5694
rect 32060 5630 32062 5682
rect 32114 5630 32116 5682
rect 32060 5234 32116 5630
rect 32060 5182 32062 5234
rect 32114 5182 32116 5234
rect 32060 5170 32116 5182
rect 31276 5070 31278 5122
rect 31330 5070 31332 5122
rect 30940 5058 30996 5068
rect 31276 5012 31332 5070
rect 31276 4946 31332 4956
rect 31948 5012 32004 5022
rect 29596 4900 29652 4910
rect 29596 4806 29652 4844
rect 31164 4900 31220 4910
rect 31164 4450 31220 4844
rect 31164 4398 31166 4450
rect 31218 4398 31220 4450
rect 31164 4386 31220 4398
rect 31948 4338 32004 4956
rect 31948 4286 31950 4338
rect 32002 4286 32004 4338
rect 31948 4274 32004 4286
rect 29036 4228 29092 4238
rect 28924 4226 29092 4228
rect 28924 4174 29038 4226
rect 29090 4174 29092 4226
rect 28924 4172 29092 4174
rect 25788 4162 25844 4172
rect 29036 4162 29092 4172
rect 23996 4114 24052 4126
rect 23996 4062 23998 4114
rect 24050 4062 24052 4114
rect 23996 3892 24052 4062
rect 25228 4116 25284 4126
rect 23996 3836 24724 3892
rect 23660 3668 23716 3678
rect 23548 3666 23716 3668
rect 23548 3614 23662 3666
rect 23714 3614 23716 3666
rect 23548 3612 23716 3614
rect 22764 3602 22820 3612
rect 23660 3602 23716 3612
rect 24556 3668 24612 3678
rect 24556 3574 24612 3612
rect 24668 3666 24724 3836
rect 24668 3614 24670 3666
rect 24722 3614 24724 3666
rect 24668 3602 24724 3614
rect 22428 3490 22484 3500
rect 24892 3556 24948 3566
rect 24892 3462 24948 3500
rect 25228 3554 25284 4060
rect 30318 3948 30582 3958
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30318 3882 30582 3892
rect 32396 3668 32452 13580
rect 33068 13636 33124 14476
rect 33180 13746 33236 15148
rect 33404 15138 33460 15148
rect 34476 14140 34740 14150
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34476 14074 34740 14084
rect 33628 13748 33684 13758
rect 33180 13694 33182 13746
rect 33234 13694 33236 13746
rect 33180 13682 33236 13694
rect 33404 13746 33684 13748
rect 33404 13694 33630 13746
rect 33682 13694 33684 13746
rect 33404 13692 33684 13694
rect 33068 13570 33124 13580
rect 33292 13524 33348 13534
rect 33292 13430 33348 13468
rect 33404 13074 33460 13692
rect 33628 13682 33684 13692
rect 33516 13524 33572 13534
rect 33516 13430 33572 13468
rect 33404 13022 33406 13074
rect 33458 13022 33460 13074
rect 33404 13010 33460 13022
rect 34076 12962 34132 12974
rect 34076 12910 34078 12962
rect 34130 12910 34132 12962
rect 33292 11956 33348 11966
rect 33348 11900 33460 11956
rect 33292 11890 33348 11900
rect 33404 11506 33460 11900
rect 33404 11454 33406 11506
rect 33458 11454 33460 11506
rect 33404 11442 33460 11454
rect 34076 11394 34132 12910
rect 34476 12572 34740 12582
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34476 12506 34740 12516
rect 34076 11342 34078 11394
rect 34130 11342 34132 11394
rect 33068 9940 33124 9950
rect 33068 9042 33124 9884
rect 34076 9826 34132 11342
rect 34476 11004 34740 11014
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34476 10938 34740 10948
rect 34076 9774 34078 9826
rect 34130 9774 34132 9826
rect 33404 9716 33460 9726
rect 33180 9714 33460 9716
rect 33180 9662 33406 9714
rect 33458 9662 33460 9714
rect 33180 9660 33460 9662
rect 33180 9266 33236 9660
rect 33404 9650 33460 9660
rect 33180 9214 33182 9266
rect 33234 9214 33236 9266
rect 33180 9202 33236 9214
rect 34076 9156 34132 9774
rect 34476 9436 34740 9446
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34476 9370 34740 9380
rect 34076 9090 34132 9100
rect 33068 8990 33070 9042
rect 33122 8990 33124 9042
rect 33068 8978 33124 8990
rect 33292 9044 33348 9054
rect 33292 8950 33348 8988
rect 33516 8818 33572 8830
rect 33516 8766 33518 8818
rect 33570 8766 33572 8818
rect 33404 8372 33460 8382
rect 32620 7588 32676 7598
rect 33180 7588 33236 7598
rect 32620 7586 33236 7588
rect 32620 7534 32622 7586
rect 32674 7534 33182 7586
rect 33234 7534 33236 7586
rect 32620 7532 33236 7534
rect 32620 7522 32676 7532
rect 33180 7522 33236 7532
rect 33404 7588 33460 8316
rect 33404 7474 33460 7532
rect 33404 7422 33406 7474
rect 33458 7422 33460 7474
rect 33404 7410 33460 7422
rect 33068 7250 33124 7262
rect 33068 7198 33070 7250
rect 33122 7198 33124 7250
rect 33068 6916 33124 7198
rect 33516 7252 33572 8766
rect 34188 8372 34244 8382
rect 34188 8278 34244 8316
rect 34476 7868 34740 7878
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34476 7802 34740 7812
rect 33516 7186 33572 7196
rect 33068 6850 33124 6860
rect 33964 6804 34020 6814
rect 33628 6802 34020 6804
rect 33628 6750 33966 6802
rect 34018 6750 34020 6802
rect 33628 6748 34020 6750
rect 33068 6244 33124 6254
rect 32956 5908 33012 5918
rect 32956 5814 33012 5852
rect 33068 4562 33124 6188
rect 33628 6132 33684 6748
rect 33964 6738 34020 6748
rect 34476 6300 34740 6310
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34476 6234 34740 6244
rect 33404 6076 33796 6132
rect 33404 6020 33460 6076
rect 33404 5926 33460 5964
rect 33628 5908 33684 5918
rect 33516 5906 33684 5908
rect 33516 5854 33630 5906
rect 33682 5854 33684 5906
rect 33516 5852 33684 5854
rect 33180 5796 33236 5806
rect 33180 5702 33236 5740
rect 33068 4510 33070 4562
rect 33122 4510 33124 4562
rect 33068 4498 33124 4510
rect 33516 5236 33572 5852
rect 33628 5842 33684 5852
rect 33404 4340 33460 4350
rect 33516 4340 33572 5180
rect 33404 4338 33572 4340
rect 33404 4286 33406 4338
rect 33458 4286 33572 4338
rect 33404 4284 33572 4286
rect 33628 4340 33684 4350
rect 33740 4340 33796 6076
rect 34188 5236 34244 5246
rect 34188 5142 34244 5180
rect 34476 4732 34740 4742
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34476 4666 34740 4676
rect 33628 4338 33796 4340
rect 33628 4286 33630 4338
rect 33682 4286 33796 4338
rect 33628 4284 33796 4286
rect 33404 4274 33460 4284
rect 33628 4274 33684 4284
rect 32956 3668 33012 3678
rect 32396 3666 33012 3668
rect 32396 3614 32958 3666
rect 33010 3614 33012 3666
rect 32396 3612 33012 3614
rect 25228 3502 25230 3554
rect 25282 3502 25284 3554
rect 25228 3490 25284 3502
rect 31500 3556 31556 3566
rect 19628 3276 19908 3332
rect 25116 3444 25172 3454
rect 17948 2492 18340 2548
rect 17948 800 18004 2492
rect 25116 800 25172 3388
rect 26908 3444 26964 3482
rect 26908 3378 26964 3388
rect 30044 3444 30100 3482
rect 31500 3462 31556 3500
rect 32172 3556 32228 3566
rect 30044 3378 30100 3388
rect 32172 3442 32228 3500
rect 32396 3554 32452 3612
rect 32956 3602 33012 3612
rect 32396 3502 32398 3554
rect 32450 3502 32452 3554
rect 32396 3490 32452 3502
rect 32172 3390 32174 3442
rect 32226 3390 32228 3442
rect 32172 3378 32228 3390
rect 32284 3444 32340 3454
rect 26160 3164 26424 3174
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26160 3098 26424 3108
rect 32284 800 32340 3388
rect 34476 3164 34740 3174
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34476 3098 34740 3108
rect 3584 0 3696 800
rect 10752 0 10864 800
rect 17920 0 18032 800
rect 25088 0 25200 800
rect 32256 0 32368 800
<< via2 >>
rect 5370 32170 5426 32172
rect 5370 32118 5372 32170
rect 5372 32118 5424 32170
rect 5424 32118 5426 32170
rect 5370 32116 5426 32118
rect 5474 32170 5530 32172
rect 5474 32118 5476 32170
rect 5476 32118 5528 32170
rect 5528 32118 5530 32170
rect 5474 32116 5530 32118
rect 5578 32170 5634 32172
rect 5578 32118 5580 32170
rect 5580 32118 5632 32170
rect 5632 32118 5634 32170
rect 5578 32116 5634 32118
rect 13686 32170 13742 32172
rect 13686 32118 13688 32170
rect 13688 32118 13740 32170
rect 13740 32118 13742 32170
rect 13686 32116 13742 32118
rect 13790 32170 13846 32172
rect 13790 32118 13792 32170
rect 13792 32118 13844 32170
rect 13844 32118 13846 32170
rect 13790 32116 13846 32118
rect 13894 32170 13950 32172
rect 13894 32118 13896 32170
rect 13896 32118 13948 32170
rect 13948 32118 13950 32170
rect 13894 32116 13950 32118
rect 22002 32170 22058 32172
rect 22002 32118 22004 32170
rect 22004 32118 22056 32170
rect 22056 32118 22058 32170
rect 22002 32116 22058 32118
rect 22106 32170 22162 32172
rect 22106 32118 22108 32170
rect 22108 32118 22160 32170
rect 22160 32118 22162 32170
rect 22106 32116 22162 32118
rect 22210 32170 22266 32172
rect 22210 32118 22212 32170
rect 22212 32118 22264 32170
rect 22264 32118 22266 32170
rect 22210 32116 22266 32118
rect 30318 32170 30374 32172
rect 30318 32118 30320 32170
rect 30320 32118 30372 32170
rect 30372 32118 30374 32170
rect 30318 32116 30374 32118
rect 30422 32170 30478 32172
rect 30422 32118 30424 32170
rect 30424 32118 30476 32170
rect 30476 32118 30478 32170
rect 30422 32116 30478 32118
rect 30526 32170 30582 32172
rect 30526 32118 30528 32170
rect 30528 32118 30580 32170
rect 30580 32118 30582 32170
rect 30526 32116 30582 32118
rect 9528 31386 9584 31388
rect 9528 31334 9530 31386
rect 9530 31334 9582 31386
rect 9582 31334 9584 31386
rect 9528 31332 9584 31334
rect 9632 31386 9688 31388
rect 9632 31334 9634 31386
rect 9634 31334 9686 31386
rect 9686 31334 9688 31386
rect 9632 31332 9688 31334
rect 9736 31386 9792 31388
rect 9736 31334 9738 31386
rect 9738 31334 9790 31386
rect 9790 31334 9792 31386
rect 9736 31332 9792 31334
rect 17844 31386 17900 31388
rect 17844 31334 17846 31386
rect 17846 31334 17898 31386
rect 17898 31334 17900 31386
rect 17844 31332 17900 31334
rect 17948 31386 18004 31388
rect 17948 31334 17950 31386
rect 17950 31334 18002 31386
rect 18002 31334 18004 31386
rect 17948 31332 18004 31334
rect 18052 31386 18108 31388
rect 18052 31334 18054 31386
rect 18054 31334 18106 31386
rect 18106 31334 18108 31386
rect 18052 31332 18108 31334
rect 26160 31386 26216 31388
rect 26160 31334 26162 31386
rect 26162 31334 26214 31386
rect 26214 31334 26216 31386
rect 26160 31332 26216 31334
rect 26264 31386 26320 31388
rect 26264 31334 26266 31386
rect 26266 31334 26318 31386
rect 26318 31334 26320 31386
rect 26264 31332 26320 31334
rect 26368 31386 26424 31388
rect 26368 31334 26370 31386
rect 26370 31334 26422 31386
rect 26422 31334 26424 31386
rect 26368 31332 26424 31334
rect 34476 31386 34532 31388
rect 34476 31334 34478 31386
rect 34478 31334 34530 31386
rect 34530 31334 34532 31386
rect 34476 31332 34532 31334
rect 34580 31386 34636 31388
rect 34580 31334 34582 31386
rect 34582 31334 34634 31386
rect 34634 31334 34636 31386
rect 34580 31332 34636 31334
rect 34684 31386 34740 31388
rect 34684 31334 34686 31386
rect 34686 31334 34738 31386
rect 34738 31334 34740 31386
rect 34684 31332 34740 31334
rect 5370 30602 5426 30604
rect 5370 30550 5372 30602
rect 5372 30550 5424 30602
rect 5424 30550 5426 30602
rect 5370 30548 5426 30550
rect 5474 30602 5530 30604
rect 5474 30550 5476 30602
rect 5476 30550 5528 30602
rect 5528 30550 5530 30602
rect 5474 30548 5530 30550
rect 5578 30602 5634 30604
rect 5578 30550 5580 30602
rect 5580 30550 5632 30602
rect 5632 30550 5634 30602
rect 5578 30548 5634 30550
rect 13686 30602 13742 30604
rect 13686 30550 13688 30602
rect 13688 30550 13740 30602
rect 13740 30550 13742 30602
rect 13686 30548 13742 30550
rect 13790 30602 13846 30604
rect 13790 30550 13792 30602
rect 13792 30550 13844 30602
rect 13844 30550 13846 30602
rect 13790 30548 13846 30550
rect 13894 30602 13950 30604
rect 13894 30550 13896 30602
rect 13896 30550 13948 30602
rect 13948 30550 13950 30602
rect 13894 30548 13950 30550
rect 22002 30602 22058 30604
rect 22002 30550 22004 30602
rect 22004 30550 22056 30602
rect 22056 30550 22058 30602
rect 22002 30548 22058 30550
rect 22106 30602 22162 30604
rect 22106 30550 22108 30602
rect 22108 30550 22160 30602
rect 22160 30550 22162 30602
rect 22106 30548 22162 30550
rect 22210 30602 22266 30604
rect 22210 30550 22212 30602
rect 22212 30550 22264 30602
rect 22264 30550 22266 30602
rect 22210 30548 22266 30550
rect 30318 30602 30374 30604
rect 30318 30550 30320 30602
rect 30320 30550 30372 30602
rect 30372 30550 30374 30602
rect 30318 30548 30374 30550
rect 30422 30602 30478 30604
rect 30422 30550 30424 30602
rect 30424 30550 30476 30602
rect 30476 30550 30478 30602
rect 30422 30548 30478 30550
rect 30526 30602 30582 30604
rect 30526 30550 30528 30602
rect 30528 30550 30580 30602
rect 30580 30550 30582 30602
rect 30526 30548 30582 30550
rect 9528 29818 9584 29820
rect 9528 29766 9530 29818
rect 9530 29766 9582 29818
rect 9582 29766 9584 29818
rect 9528 29764 9584 29766
rect 9632 29818 9688 29820
rect 9632 29766 9634 29818
rect 9634 29766 9686 29818
rect 9686 29766 9688 29818
rect 9632 29764 9688 29766
rect 9736 29818 9792 29820
rect 9736 29766 9738 29818
rect 9738 29766 9790 29818
rect 9790 29766 9792 29818
rect 9736 29764 9792 29766
rect 17844 29818 17900 29820
rect 17844 29766 17846 29818
rect 17846 29766 17898 29818
rect 17898 29766 17900 29818
rect 17844 29764 17900 29766
rect 17948 29818 18004 29820
rect 17948 29766 17950 29818
rect 17950 29766 18002 29818
rect 18002 29766 18004 29818
rect 17948 29764 18004 29766
rect 18052 29818 18108 29820
rect 18052 29766 18054 29818
rect 18054 29766 18106 29818
rect 18106 29766 18108 29818
rect 18052 29764 18108 29766
rect 26160 29818 26216 29820
rect 26160 29766 26162 29818
rect 26162 29766 26214 29818
rect 26214 29766 26216 29818
rect 26160 29764 26216 29766
rect 26264 29818 26320 29820
rect 26264 29766 26266 29818
rect 26266 29766 26318 29818
rect 26318 29766 26320 29818
rect 26264 29764 26320 29766
rect 26368 29818 26424 29820
rect 26368 29766 26370 29818
rect 26370 29766 26422 29818
rect 26422 29766 26424 29818
rect 26368 29764 26424 29766
rect 34476 29818 34532 29820
rect 34476 29766 34478 29818
rect 34478 29766 34530 29818
rect 34530 29766 34532 29818
rect 34476 29764 34532 29766
rect 34580 29818 34636 29820
rect 34580 29766 34582 29818
rect 34582 29766 34634 29818
rect 34634 29766 34636 29818
rect 34580 29764 34636 29766
rect 34684 29818 34740 29820
rect 34684 29766 34686 29818
rect 34686 29766 34738 29818
rect 34738 29766 34740 29818
rect 34684 29764 34740 29766
rect 5370 29034 5426 29036
rect 5370 28982 5372 29034
rect 5372 28982 5424 29034
rect 5424 28982 5426 29034
rect 5370 28980 5426 28982
rect 5474 29034 5530 29036
rect 5474 28982 5476 29034
rect 5476 28982 5528 29034
rect 5528 28982 5530 29034
rect 5474 28980 5530 28982
rect 5578 29034 5634 29036
rect 5578 28982 5580 29034
rect 5580 28982 5632 29034
rect 5632 28982 5634 29034
rect 5578 28980 5634 28982
rect 13686 29034 13742 29036
rect 13686 28982 13688 29034
rect 13688 28982 13740 29034
rect 13740 28982 13742 29034
rect 13686 28980 13742 28982
rect 13790 29034 13846 29036
rect 13790 28982 13792 29034
rect 13792 28982 13844 29034
rect 13844 28982 13846 29034
rect 13790 28980 13846 28982
rect 13894 29034 13950 29036
rect 13894 28982 13896 29034
rect 13896 28982 13948 29034
rect 13948 28982 13950 29034
rect 13894 28980 13950 28982
rect 22002 29034 22058 29036
rect 22002 28982 22004 29034
rect 22004 28982 22056 29034
rect 22056 28982 22058 29034
rect 22002 28980 22058 28982
rect 22106 29034 22162 29036
rect 22106 28982 22108 29034
rect 22108 28982 22160 29034
rect 22160 28982 22162 29034
rect 22106 28980 22162 28982
rect 22210 29034 22266 29036
rect 22210 28982 22212 29034
rect 22212 28982 22264 29034
rect 22264 28982 22266 29034
rect 22210 28980 22266 28982
rect 30318 29034 30374 29036
rect 30318 28982 30320 29034
rect 30320 28982 30372 29034
rect 30372 28982 30374 29034
rect 30318 28980 30374 28982
rect 30422 29034 30478 29036
rect 30422 28982 30424 29034
rect 30424 28982 30476 29034
rect 30476 28982 30478 29034
rect 30422 28980 30478 28982
rect 30526 29034 30582 29036
rect 30526 28982 30528 29034
rect 30528 28982 30580 29034
rect 30580 28982 30582 29034
rect 30526 28980 30582 28982
rect 2492 26348 2548 26404
rect 9528 28250 9584 28252
rect 9528 28198 9530 28250
rect 9530 28198 9582 28250
rect 9582 28198 9584 28250
rect 9528 28196 9584 28198
rect 9632 28250 9688 28252
rect 9632 28198 9634 28250
rect 9634 28198 9686 28250
rect 9686 28198 9688 28250
rect 9632 28196 9688 28198
rect 9736 28250 9792 28252
rect 9736 28198 9738 28250
rect 9738 28198 9790 28250
rect 9790 28198 9792 28250
rect 9736 28196 9792 28198
rect 8428 27804 8484 27860
rect 5370 27466 5426 27468
rect 5370 27414 5372 27466
rect 5372 27414 5424 27466
rect 5424 27414 5426 27466
rect 5370 27412 5426 27414
rect 5474 27466 5530 27468
rect 5474 27414 5476 27466
rect 5476 27414 5528 27466
rect 5528 27414 5530 27466
rect 5474 27412 5530 27414
rect 5578 27466 5634 27468
rect 5578 27414 5580 27466
rect 5580 27414 5632 27466
rect 5632 27414 5634 27466
rect 5578 27412 5634 27414
rect 5180 27244 5236 27300
rect 5852 27298 5908 27300
rect 5852 27246 5854 27298
rect 5854 27246 5906 27298
rect 5906 27246 5908 27298
rect 5852 27244 5908 27246
rect 5964 27074 6020 27076
rect 5964 27022 5966 27074
rect 5966 27022 6018 27074
rect 6018 27022 6020 27074
rect 5964 27020 6020 27022
rect 4956 26908 5012 26964
rect 3276 26348 3332 26404
rect 1820 25452 1876 25508
rect 2492 22540 2548 22596
rect 3276 24892 3332 24948
rect 4060 24834 4116 24836
rect 4060 24782 4062 24834
rect 4062 24782 4114 24834
rect 4114 24782 4116 24834
rect 4060 24780 4116 24782
rect 4620 25340 4676 25396
rect 5068 25340 5124 25396
rect 5180 26908 5236 26964
rect 5068 24892 5124 24948
rect 4620 24668 4676 24724
rect 4396 24108 4452 24164
rect 5370 25898 5426 25900
rect 5370 25846 5372 25898
rect 5372 25846 5424 25898
rect 5424 25846 5426 25898
rect 5370 25844 5426 25846
rect 5474 25898 5530 25900
rect 5474 25846 5476 25898
rect 5476 25846 5528 25898
rect 5528 25846 5530 25898
rect 5474 25844 5530 25846
rect 5578 25898 5634 25900
rect 5578 25846 5580 25898
rect 5580 25846 5632 25898
rect 5632 25846 5634 25898
rect 5578 25844 5634 25846
rect 5852 25340 5908 25396
rect 5740 24780 5796 24836
rect 5628 24722 5684 24724
rect 5628 24670 5630 24722
rect 5630 24670 5682 24722
rect 5682 24670 5684 24722
rect 5628 24668 5684 24670
rect 5370 24330 5426 24332
rect 5370 24278 5372 24330
rect 5372 24278 5424 24330
rect 5424 24278 5426 24330
rect 5370 24276 5426 24278
rect 5474 24330 5530 24332
rect 5474 24278 5476 24330
rect 5476 24278 5528 24330
rect 5528 24278 5530 24330
rect 5474 24276 5530 24278
rect 5578 24330 5634 24332
rect 5578 24278 5580 24330
rect 5580 24278 5632 24330
rect 5632 24278 5634 24330
rect 5578 24276 5634 24278
rect 2716 22876 2772 22932
rect 3612 22316 3668 22372
rect 3948 21698 4004 21700
rect 3948 21646 3950 21698
rect 3950 21646 4002 21698
rect 4002 21646 4004 21698
rect 3948 21644 4004 21646
rect 4956 23212 5012 23268
rect 4844 21756 4900 21812
rect 5370 22762 5426 22764
rect 5370 22710 5372 22762
rect 5372 22710 5424 22762
rect 5424 22710 5426 22762
rect 5370 22708 5426 22710
rect 5474 22762 5530 22764
rect 5474 22710 5476 22762
rect 5476 22710 5528 22762
rect 5528 22710 5530 22762
rect 5474 22708 5530 22710
rect 5578 22762 5634 22764
rect 5578 22710 5580 22762
rect 5580 22710 5632 22762
rect 5632 22710 5634 22762
rect 5578 22708 5634 22710
rect 5628 22594 5684 22596
rect 5628 22542 5630 22594
rect 5630 22542 5682 22594
rect 5682 22542 5684 22594
rect 5628 22540 5684 22542
rect 6748 27074 6804 27076
rect 6748 27022 6750 27074
rect 6750 27022 6802 27074
rect 6802 27022 6804 27074
rect 6748 27020 6804 27022
rect 6300 26348 6356 26404
rect 6412 26908 6468 26964
rect 6076 24892 6132 24948
rect 5852 23212 5908 23268
rect 6076 22370 6132 22372
rect 6076 22318 6078 22370
rect 6078 22318 6130 22370
rect 6130 22318 6132 22370
rect 6076 22316 6132 22318
rect 5516 21810 5572 21812
rect 5516 21758 5518 21810
rect 5518 21758 5570 21810
rect 5570 21758 5572 21810
rect 5516 21756 5572 21758
rect 4620 21698 4676 21700
rect 4620 21646 4622 21698
rect 4622 21646 4674 21698
rect 4674 21646 4676 21698
rect 4620 21644 4676 21646
rect 5404 21698 5460 21700
rect 5404 21646 5406 21698
rect 5406 21646 5458 21698
rect 5458 21646 5460 21698
rect 5404 21644 5460 21646
rect 3276 20802 3332 20804
rect 3276 20750 3278 20802
rect 3278 20750 3330 20802
rect 3330 20750 3332 20802
rect 3276 20748 3332 20750
rect 2380 20578 2436 20580
rect 2380 20526 2382 20578
rect 2382 20526 2434 20578
rect 2434 20526 2436 20578
rect 2380 20524 2436 20526
rect 2940 20578 2996 20580
rect 2940 20526 2942 20578
rect 2942 20526 2994 20578
rect 2994 20526 2996 20578
rect 2940 20524 2996 20526
rect 3388 20524 3444 20580
rect 5370 21194 5426 21196
rect 5370 21142 5372 21194
rect 5372 21142 5424 21194
rect 5424 21142 5426 21194
rect 5370 21140 5426 21142
rect 5474 21194 5530 21196
rect 5474 21142 5476 21194
rect 5476 21142 5528 21194
rect 5528 21142 5530 21194
rect 5474 21140 5530 21142
rect 5578 21194 5634 21196
rect 5578 21142 5580 21194
rect 5580 21142 5632 21194
rect 5632 21142 5634 21194
rect 5578 21140 5634 21142
rect 4284 20748 4340 20804
rect 3948 20690 4004 20692
rect 3948 20638 3950 20690
rect 3950 20638 4002 20690
rect 4002 20638 4004 20690
rect 3948 20636 4004 20638
rect 3612 19964 3668 20020
rect 2492 19852 2548 19908
rect 4284 20578 4340 20580
rect 4284 20526 4286 20578
rect 4286 20526 4338 20578
rect 4338 20526 4340 20578
rect 4284 20524 4340 20526
rect 4396 20076 4452 20132
rect 4732 20748 4788 20804
rect 4620 20636 4676 20692
rect 4844 20524 4900 20580
rect 4508 19964 4564 20020
rect 6860 26962 6916 26964
rect 6860 26910 6862 26962
rect 6862 26910 6914 26962
rect 6914 26910 6916 26962
rect 6860 26908 6916 26910
rect 7308 26402 7364 26404
rect 7308 26350 7310 26402
rect 7310 26350 7362 26402
rect 7362 26350 7364 26402
rect 7308 26348 7364 26350
rect 6636 24892 6692 24948
rect 7084 25506 7140 25508
rect 7084 25454 7086 25506
rect 7086 25454 7138 25506
rect 7138 25454 7140 25506
rect 7084 25452 7140 25454
rect 6300 24108 6356 24164
rect 8204 26460 8260 26516
rect 7420 25452 7476 25508
rect 9528 26682 9584 26684
rect 9528 26630 9530 26682
rect 9530 26630 9582 26682
rect 9582 26630 9584 26682
rect 9528 26628 9584 26630
rect 9632 26682 9688 26684
rect 9632 26630 9634 26682
rect 9634 26630 9686 26682
rect 9686 26630 9688 26682
rect 9632 26628 9688 26630
rect 9736 26682 9792 26684
rect 9736 26630 9738 26682
rect 9738 26630 9790 26682
rect 9790 26630 9792 26682
rect 9736 26628 9792 26630
rect 8876 26460 8932 26516
rect 7980 25452 8036 25508
rect 10220 27858 10276 27860
rect 10220 27806 10222 27858
rect 10222 27806 10274 27858
rect 10274 27806 10276 27858
rect 10220 27804 10276 27806
rect 11004 27746 11060 27748
rect 11004 27694 11006 27746
rect 11006 27694 11058 27746
rect 11058 27694 11060 27746
rect 11004 27692 11060 27694
rect 9528 25114 9584 25116
rect 9528 25062 9530 25114
rect 9530 25062 9582 25114
rect 9582 25062 9584 25114
rect 9528 25060 9584 25062
rect 9632 25114 9688 25116
rect 9632 25062 9634 25114
rect 9634 25062 9686 25114
rect 9686 25062 9688 25114
rect 9632 25060 9688 25062
rect 9736 25114 9792 25116
rect 9736 25062 9738 25114
rect 9738 25062 9790 25114
rect 9790 25062 9792 25114
rect 9736 25060 9792 25062
rect 7756 24108 7812 24164
rect 8764 24108 8820 24164
rect 6412 22930 6468 22932
rect 6412 22878 6414 22930
rect 6414 22878 6466 22930
rect 6466 22878 6468 22930
rect 6412 22876 6468 22878
rect 6300 22540 6356 22596
rect 8988 23996 9044 24052
rect 9528 23546 9584 23548
rect 9528 23494 9530 23546
rect 9530 23494 9582 23546
rect 9582 23494 9584 23546
rect 9528 23492 9584 23494
rect 9632 23546 9688 23548
rect 9632 23494 9634 23546
rect 9634 23494 9686 23546
rect 9686 23494 9688 23546
rect 9632 23492 9688 23494
rect 9736 23546 9792 23548
rect 9736 23494 9738 23546
rect 9738 23494 9790 23546
rect 9790 23494 9792 23546
rect 9736 23492 9792 23494
rect 9996 24892 10052 24948
rect 17844 28250 17900 28252
rect 17844 28198 17846 28250
rect 17846 28198 17898 28250
rect 17898 28198 17900 28250
rect 17844 28196 17900 28198
rect 17948 28250 18004 28252
rect 17948 28198 17950 28250
rect 17950 28198 18002 28250
rect 18002 28198 18004 28250
rect 17948 28196 18004 28198
rect 18052 28250 18108 28252
rect 18052 28198 18054 28250
rect 18054 28198 18106 28250
rect 18106 28198 18108 28250
rect 18052 28196 18108 28198
rect 26160 28250 26216 28252
rect 26160 28198 26162 28250
rect 26162 28198 26214 28250
rect 26214 28198 26216 28250
rect 26160 28196 26216 28198
rect 26264 28250 26320 28252
rect 26264 28198 26266 28250
rect 26266 28198 26318 28250
rect 26318 28198 26320 28250
rect 26264 28196 26320 28198
rect 26368 28250 26424 28252
rect 26368 28198 26370 28250
rect 26370 28198 26422 28250
rect 26422 28198 26424 28250
rect 26368 28196 26424 28198
rect 34476 28250 34532 28252
rect 34476 28198 34478 28250
rect 34478 28198 34530 28250
rect 34530 28198 34532 28250
rect 34476 28196 34532 28198
rect 34580 28250 34636 28252
rect 34580 28198 34582 28250
rect 34582 28198 34634 28250
rect 34634 28198 34636 28250
rect 34580 28196 34636 28198
rect 34684 28250 34740 28252
rect 34684 28198 34686 28250
rect 34686 28198 34738 28250
rect 34738 28198 34740 28250
rect 34684 28196 34740 28198
rect 19068 27804 19124 27860
rect 12236 27692 12292 27748
rect 12460 27074 12516 27076
rect 12460 27022 12462 27074
rect 12462 27022 12514 27074
rect 12514 27022 12516 27074
rect 12460 27020 12516 27022
rect 11004 25676 11060 25732
rect 12012 25506 12068 25508
rect 12012 25454 12014 25506
rect 12014 25454 12066 25506
rect 12066 25454 12068 25506
rect 12012 25452 12068 25454
rect 10332 24556 10388 24612
rect 9996 24108 10052 24164
rect 10780 23884 10836 23940
rect 9996 23378 10052 23380
rect 9996 23326 9998 23378
rect 9998 23326 10050 23378
rect 10050 23326 10052 23378
rect 9996 23324 10052 23326
rect 9884 23266 9940 23268
rect 9884 23214 9886 23266
rect 9886 23214 9938 23266
rect 9938 23214 9940 23266
rect 9884 23212 9940 23214
rect 7084 22428 7140 22484
rect 7868 22482 7924 22484
rect 7868 22430 7870 22482
rect 7870 22430 7922 22482
rect 7922 22430 7924 22482
rect 7868 22428 7924 22430
rect 8876 23042 8932 23044
rect 8876 22990 8878 23042
rect 8878 22990 8930 23042
rect 8930 22990 8932 23042
rect 8876 22988 8932 22990
rect 8428 22204 8484 22260
rect 9528 21978 9584 21980
rect 9528 21926 9530 21978
rect 9530 21926 9582 21978
rect 9582 21926 9584 21978
rect 9528 21924 9584 21926
rect 9632 21978 9688 21980
rect 9632 21926 9634 21978
rect 9634 21926 9686 21978
rect 9686 21926 9688 21978
rect 9632 21924 9688 21926
rect 9736 21978 9792 21980
rect 9736 21926 9738 21978
rect 9738 21926 9790 21978
rect 9790 21926 9792 21978
rect 9736 21924 9792 21926
rect 10332 21532 10388 21588
rect 7644 20802 7700 20804
rect 7644 20750 7646 20802
rect 7646 20750 7698 20802
rect 7698 20750 7700 20802
rect 7644 20748 7700 20750
rect 8204 20690 8260 20692
rect 8204 20638 8206 20690
rect 8206 20638 8258 20690
rect 8258 20638 8260 20690
rect 8204 20636 8260 20638
rect 4956 20188 5012 20244
rect 5404 20076 5460 20132
rect 5180 20018 5236 20020
rect 5180 19966 5182 20018
rect 5182 19966 5234 20018
rect 5234 19966 5236 20018
rect 5180 19964 5236 19966
rect 7308 19964 7364 20020
rect 5068 19906 5124 19908
rect 5068 19854 5070 19906
rect 5070 19854 5122 19906
rect 5122 19854 5124 19906
rect 5068 19852 5124 19854
rect 5370 19626 5426 19628
rect 5370 19574 5372 19626
rect 5372 19574 5424 19626
rect 5424 19574 5426 19626
rect 5370 19572 5426 19574
rect 5474 19626 5530 19628
rect 5474 19574 5476 19626
rect 5476 19574 5528 19626
rect 5528 19574 5530 19626
rect 5474 19572 5530 19574
rect 5578 19626 5634 19628
rect 5578 19574 5580 19626
rect 5580 19574 5632 19626
rect 5632 19574 5634 19626
rect 5578 19572 5634 19574
rect 6972 18732 7028 18788
rect 6748 18508 6804 18564
rect 5370 18058 5426 18060
rect 5370 18006 5372 18058
rect 5372 18006 5424 18058
rect 5424 18006 5426 18058
rect 5370 18004 5426 18006
rect 5474 18058 5530 18060
rect 5474 18006 5476 18058
rect 5476 18006 5528 18058
rect 5528 18006 5530 18058
rect 5474 18004 5530 18006
rect 5578 18058 5634 18060
rect 5578 18006 5580 18058
rect 5580 18006 5632 18058
rect 5632 18006 5634 18058
rect 5578 18004 5634 18006
rect 1596 15148 1652 15204
rect 4620 17612 4676 17668
rect 5740 17666 5796 17668
rect 5740 17614 5742 17666
rect 5742 17614 5794 17666
rect 5794 17614 5796 17666
rect 5740 17612 5796 17614
rect 1820 15036 1876 15092
rect 2268 15036 2324 15092
rect 5964 17554 6020 17556
rect 5964 17502 5966 17554
rect 5966 17502 6018 17554
rect 6018 17502 6020 17554
rect 5964 17500 6020 17502
rect 5068 16940 5124 16996
rect 3948 16882 4004 16884
rect 3948 16830 3950 16882
rect 3950 16830 4002 16882
rect 4002 16830 4004 16882
rect 3948 16828 4004 16830
rect 5852 16828 5908 16884
rect 5370 16490 5426 16492
rect 5370 16438 5372 16490
rect 5372 16438 5424 16490
rect 5424 16438 5426 16490
rect 5370 16436 5426 16438
rect 5474 16490 5530 16492
rect 5474 16438 5476 16490
rect 5476 16438 5528 16490
rect 5528 16438 5530 16490
rect 5474 16436 5530 16438
rect 5578 16490 5634 16492
rect 5578 16438 5580 16490
rect 5580 16438 5632 16490
rect 5632 16438 5634 16490
rect 5578 16436 5634 16438
rect 3276 15036 3332 15092
rect 6524 17666 6580 17668
rect 6524 17614 6526 17666
rect 6526 17614 6578 17666
rect 6578 17614 6580 17666
rect 6524 17612 6580 17614
rect 6860 17890 6916 17892
rect 6860 17838 6862 17890
rect 6862 17838 6914 17890
rect 6914 17838 6916 17890
rect 6860 17836 6916 17838
rect 7980 19852 8036 19908
rect 7420 18674 7476 18676
rect 7420 18622 7422 18674
rect 7422 18622 7474 18674
rect 7474 18622 7476 18674
rect 7420 18620 7476 18622
rect 7196 17836 7252 17892
rect 7756 18508 7812 18564
rect 7644 17666 7700 17668
rect 7644 17614 7646 17666
rect 7646 17614 7698 17666
rect 7698 17614 7700 17666
rect 7644 17612 7700 17614
rect 7084 17500 7140 17556
rect 6748 16994 6804 16996
rect 6748 16942 6750 16994
rect 6750 16942 6802 16994
rect 6802 16942 6804 16994
rect 6748 16940 6804 16942
rect 7980 18562 8036 18564
rect 7980 18510 7982 18562
rect 7982 18510 8034 18562
rect 8034 18510 8036 18562
rect 7980 18508 8036 18510
rect 7756 17052 7812 17108
rect 7196 16940 7252 16996
rect 6300 16828 6356 16884
rect 9884 20524 9940 20580
rect 9528 20410 9584 20412
rect 9528 20358 9530 20410
rect 9530 20358 9582 20410
rect 9582 20358 9584 20410
rect 9528 20356 9584 20358
rect 9632 20410 9688 20412
rect 9632 20358 9634 20410
rect 9634 20358 9686 20410
rect 9686 20358 9688 20410
rect 9632 20356 9688 20358
rect 9736 20410 9792 20412
rect 9736 20358 9738 20410
rect 9738 20358 9790 20410
rect 9790 20358 9792 20410
rect 9736 20356 9792 20358
rect 8204 20130 8260 20132
rect 8204 20078 8206 20130
rect 8206 20078 8258 20130
rect 8258 20078 8260 20130
rect 8204 20076 8260 20078
rect 8876 19964 8932 20020
rect 9436 19964 9492 20020
rect 8988 19346 9044 19348
rect 8988 19294 8990 19346
rect 8990 19294 9042 19346
rect 9042 19294 9044 19346
rect 8988 19292 9044 19294
rect 8204 18732 8260 18788
rect 8204 18060 8260 18116
rect 8092 17276 8148 17332
rect 8316 17612 8372 17668
rect 9996 20188 10052 20244
rect 11116 24946 11172 24948
rect 11116 24894 11118 24946
rect 11118 24894 11170 24946
rect 11170 24894 11172 24946
rect 11116 24892 11172 24894
rect 11116 24556 11172 24612
rect 11004 24050 11060 24052
rect 11004 23998 11006 24050
rect 11006 23998 11058 24050
rect 11058 23998 11060 24050
rect 11004 23996 11060 23998
rect 11116 23826 11172 23828
rect 11116 23774 11118 23826
rect 11118 23774 11170 23826
rect 11170 23774 11172 23826
rect 11116 23772 11172 23774
rect 11228 23884 11284 23940
rect 12348 26290 12404 26292
rect 12348 26238 12350 26290
rect 12350 26238 12402 26290
rect 12402 26238 12404 26290
rect 12348 26236 12404 26238
rect 13686 27466 13742 27468
rect 13686 27414 13688 27466
rect 13688 27414 13740 27466
rect 13740 27414 13742 27466
rect 13686 27412 13742 27414
rect 13790 27466 13846 27468
rect 13790 27414 13792 27466
rect 13792 27414 13844 27466
rect 13844 27414 13846 27466
rect 13790 27412 13846 27414
rect 13894 27466 13950 27468
rect 13894 27414 13896 27466
rect 13896 27414 13948 27466
rect 13948 27414 13950 27466
rect 13894 27412 13950 27414
rect 16380 27132 16436 27188
rect 14364 26908 14420 26964
rect 15484 26908 15540 26964
rect 13132 26236 13188 26292
rect 12684 25564 12740 25620
rect 12348 25394 12404 25396
rect 12348 25342 12350 25394
rect 12350 25342 12402 25394
rect 12402 25342 12404 25394
rect 12348 25340 12404 25342
rect 13686 25898 13742 25900
rect 13686 25846 13688 25898
rect 13688 25846 13740 25898
rect 13740 25846 13742 25898
rect 13686 25844 13742 25846
rect 13790 25898 13846 25900
rect 13790 25846 13792 25898
rect 13792 25846 13844 25898
rect 13844 25846 13846 25898
rect 13790 25844 13846 25846
rect 13894 25898 13950 25900
rect 13894 25846 13896 25898
rect 13896 25846 13948 25898
rect 13948 25846 13950 25898
rect 13894 25844 13950 25846
rect 14140 25788 14196 25844
rect 13580 25618 13636 25620
rect 13580 25566 13582 25618
rect 13582 25566 13634 25618
rect 13634 25566 13636 25618
rect 13580 25564 13636 25566
rect 13132 25452 13188 25508
rect 13692 25506 13748 25508
rect 13692 25454 13694 25506
rect 13694 25454 13746 25506
rect 13746 25454 13748 25506
rect 13692 25452 13748 25454
rect 12908 25340 12964 25396
rect 12460 25282 12516 25284
rect 12460 25230 12462 25282
rect 12462 25230 12514 25282
rect 12514 25230 12516 25282
rect 12460 25228 12516 25230
rect 13356 25004 13412 25060
rect 14028 25340 14084 25396
rect 12124 24892 12180 24948
rect 12460 24946 12516 24948
rect 12460 24894 12462 24946
rect 12462 24894 12514 24946
rect 12514 24894 12516 24946
rect 12460 24892 12516 24894
rect 11788 24780 11844 24836
rect 11564 24108 11620 24164
rect 10892 22876 10948 22932
rect 10892 22428 10948 22484
rect 11452 23212 11508 23268
rect 11004 21756 11060 21812
rect 10668 21420 10724 21476
rect 10668 21196 10724 21252
rect 10444 20578 10500 20580
rect 10444 20526 10446 20578
rect 10446 20526 10498 20578
rect 10498 20526 10500 20578
rect 10444 20524 10500 20526
rect 10220 20076 10276 20132
rect 9996 19964 10052 20020
rect 9660 19906 9716 19908
rect 9660 19854 9662 19906
rect 9662 19854 9714 19906
rect 9714 19854 9716 19906
rect 9660 19852 9716 19854
rect 10332 19852 10388 19908
rect 9772 19180 9828 19236
rect 9100 19068 9156 19124
rect 9528 18842 9584 18844
rect 9528 18790 9530 18842
rect 9530 18790 9582 18842
rect 9582 18790 9584 18842
rect 9528 18788 9584 18790
rect 9632 18842 9688 18844
rect 9632 18790 9634 18842
rect 9634 18790 9686 18842
rect 9686 18790 9688 18842
rect 9632 18788 9688 18790
rect 9736 18842 9792 18844
rect 9736 18790 9738 18842
rect 9738 18790 9790 18842
rect 9790 18790 9792 18842
rect 9736 18788 9792 18790
rect 8428 17836 8484 17892
rect 7532 16882 7588 16884
rect 7532 16830 7534 16882
rect 7534 16830 7586 16882
rect 7586 16830 7588 16882
rect 7532 16828 7588 16830
rect 7980 16940 8036 16996
rect 8204 17106 8260 17108
rect 8204 17054 8206 17106
rect 8206 17054 8258 17106
rect 8258 17054 8260 17106
rect 8204 17052 8260 17054
rect 8428 17276 8484 17332
rect 8876 18562 8932 18564
rect 8876 18510 8878 18562
rect 8878 18510 8930 18562
rect 8930 18510 8932 18562
rect 8876 18508 8932 18510
rect 8876 18226 8932 18228
rect 8876 18174 8878 18226
rect 8878 18174 8930 18226
rect 8930 18174 8932 18226
rect 8876 18172 8932 18174
rect 8540 17612 8596 17668
rect 9100 17500 9156 17556
rect 10332 19180 10388 19236
rect 9996 18956 10052 19012
rect 9660 18562 9716 18564
rect 9660 18510 9662 18562
rect 9662 18510 9714 18562
rect 9714 18510 9716 18562
rect 9660 18508 9716 18510
rect 9884 18284 9940 18340
rect 10332 18844 10388 18900
rect 10108 18226 10164 18228
rect 10108 18174 10110 18226
rect 10110 18174 10162 18226
rect 10162 18174 10164 18226
rect 10108 18172 10164 18174
rect 9548 17890 9604 17892
rect 9548 17838 9550 17890
rect 9550 17838 9602 17890
rect 9602 17838 9604 17890
rect 9548 17836 9604 17838
rect 10892 21586 10948 21588
rect 10892 21534 10894 21586
rect 10894 21534 10946 21586
rect 10946 21534 10948 21586
rect 10892 21532 10948 21534
rect 12236 24722 12292 24724
rect 12236 24670 12238 24722
rect 12238 24670 12290 24722
rect 12290 24670 12292 24722
rect 12236 24668 12292 24670
rect 12684 24834 12740 24836
rect 12684 24782 12686 24834
rect 12686 24782 12738 24834
rect 12738 24782 12740 24834
rect 12684 24780 12740 24782
rect 13132 24780 13188 24836
rect 12460 24668 12516 24724
rect 11676 23548 11732 23604
rect 11788 23884 11844 23940
rect 11340 22764 11396 22820
rect 11340 22428 11396 22484
rect 11564 21980 11620 22036
rect 12012 23826 12068 23828
rect 12012 23774 12014 23826
rect 12014 23774 12066 23826
rect 12066 23774 12068 23826
rect 12012 23772 12068 23774
rect 12236 23772 12292 23828
rect 12124 23324 12180 23380
rect 12124 23154 12180 23156
rect 12124 23102 12126 23154
rect 12126 23102 12178 23154
rect 12178 23102 12180 23154
rect 12124 23100 12180 23102
rect 12012 21420 12068 21476
rect 10780 20524 10836 20580
rect 11452 20578 11508 20580
rect 11452 20526 11454 20578
rect 11454 20526 11506 20578
rect 11506 20526 11508 20578
rect 11452 20524 11508 20526
rect 11340 20188 11396 20244
rect 10556 19292 10612 19348
rect 11004 19740 11060 19796
rect 10556 19122 10612 19124
rect 10556 19070 10558 19122
rect 10558 19070 10610 19122
rect 10610 19070 10612 19122
rect 10556 19068 10612 19070
rect 10444 18172 10500 18228
rect 10220 17666 10276 17668
rect 10220 17614 10222 17666
rect 10222 17614 10274 17666
rect 10274 17614 10276 17666
rect 10220 17612 10276 17614
rect 9772 17388 9828 17444
rect 9528 17274 9584 17276
rect 9528 17222 9530 17274
rect 9530 17222 9582 17274
rect 9582 17222 9584 17274
rect 9528 17220 9584 17222
rect 9632 17274 9688 17276
rect 9632 17222 9634 17274
rect 9634 17222 9686 17274
rect 9686 17222 9688 17274
rect 9632 17220 9688 17222
rect 9736 17274 9792 17276
rect 9736 17222 9738 17274
rect 9738 17222 9790 17274
rect 9790 17222 9792 17274
rect 9736 17220 9792 17222
rect 9884 17106 9940 17108
rect 9884 17054 9886 17106
rect 9886 17054 9938 17106
rect 9938 17054 9940 17106
rect 9884 17052 9940 17054
rect 10556 18450 10612 18452
rect 10556 18398 10558 18450
rect 10558 18398 10610 18450
rect 10610 18398 10612 18450
rect 10556 18396 10612 18398
rect 14252 25228 14308 25284
rect 14700 25506 14756 25508
rect 14700 25454 14702 25506
rect 14702 25454 14754 25506
rect 14754 25454 14756 25506
rect 14700 25452 14756 25454
rect 14028 24892 14084 24948
rect 13244 24668 13300 24724
rect 13020 23938 13076 23940
rect 13020 23886 13022 23938
rect 13022 23886 13074 23938
rect 13074 23886 13076 23938
rect 13020 23884 13076 23886
rect 12572 23772 12628 23828
rect 12348 23548 12404 23604
rect 12572 23548 12628 23604
rect 12460 23324 12516 23380
rect 12908 23378 12964 23380
rect 12908 23326 12910 23378
rect 12910 23326 12962 23378
rect 12962 23326 12964 23378
rect 12908 23324 12964 23326
rect 12684 23266 12740 23268
rect 12684 23214 12686 23266
rect 12686 23214 12738 23266
rect 12738 23214 12740 23266
rect 12684 23212 12740 23214
rect 13020 23100 13076 23156
rect 12572 23042 12628 23044
rect 12572 22990 12574 23042
rect 12574 22990 12626 23042
rect 12626 22990 12628 23042
rect 12572 22988 12628 22990
rect 12348 21868 12404 21924
rect 12908 22370 12964 22372
rect 12908 22318 12910 22370
rect 12910 22318 12962 22370
rect 12962 22318 12964 22370
rect 12908 22316 12964 22318
rect 12348 21698 12404 21700
rect 12348 21646 12350 21698
rect 12350 21646 12402 21698
rect 12402 21646 12404 21698
rect 12348 21644 12404 21646
rect 12348 21196 12404 21252
rect 12684 21810 12740 21812
rect 12684 21758 12686 21810
rect 12686 21758 12738 21810
rect 12738 21758 12740 21810
rect 12684 21756 12740 21758
rect 13020 21420 13076 21476
rect 13686 24330 13742 24332
rect 13686 24278 13688 24330
rect 13688 24278 13740 24330
rect 13740 24278 13742 24330
rect 13686 24276 13742 24278
rect 13790 24330 13846 24332
rect 13790 24278 13792 24330
rect 13792 24278 13844 24330
rect 13844 24278 13846 24330
rect 13790 24276 13846 24278
rect 13894 24330 13950 24332
rect 13894 24278 13896 24330
rect 13896 24278 13948 24330
rect 13948 24278 13950 24330
rect 13894 24276 13950 24278
rect 13692 23884 13748 23940
rect 13692 23714 13748 23716
rect 13692 23662 13694 23714
rect 13694 23662 13746 23714
rect 13746 23662 13748 23714
rect 13692 23660 13748 23662
rect 14364 25004 14420 25060
rect 14140 24108 14196 24164
rect 13916 23826 13972 23828
rect 13916 23774 13918 23826
rect 13918 23774 13970 23826
rect 13970 23774 13972 23826
rect 13916 23772 13972 23774
rect 14140 23660 14196 23716
rect 13916 23324 13972 23380
rect 13686 22762 13742 22764
rect 13686 22710 13688 22762
rect 13688 22710 13740 22762
rect 13740 22710 13742 22762
rect 13686 22708 13742 22710
rect 13790 22762 13846 22764
rect 13790 22710 13792 22762
rect 13792 22710 13844 22762
rect 13844 22710 13846 22762
rect 13790 22708 13846 22710
rect 13894 22762 13950 22764
rect 13894 22710 13896 22762
rect 13896 22710 13948 22762
rect 13948 22710 13950 22762
rect 13894 22708 13950 22710
rect 14588 24722 14644 24724
rect 14588 24670 14590 24722
rect 14590 24670 14642 24722
rect 14642 24670 14644 24722
rect 14588 24668 14644 24670
rect 14476 24332 14532 24388
rect 14924 25394 14980 25396
rect 14924 25342 14926 25394
rect 14926 25342 14978 25394
rect 14978 25342 14980 25394
rect 14924 25340 14980 25342
rect 15484 25506 15540 25508
rect 15484 25454 15486 25506
rect 15486 25454 15538 25506
rect 15538 25454 15540 25506
rect 15484 25452 15540 25454
rect 15708 26236 15764 26292
rect 15260 24946 15316 24948
rect 15260 24894 15262 24946
rect 15262 24894 15314 24946
rect 15314 24894 15316 24946
rect 15260 24892 15316 24894
rect 14476 23660 14532 23716
rect 14588 23884 14644 23940
rect 14364 23324 14420 23380
rect 14364 23100 14420 23156
rect 13580 22204 13636 22260
rect 13244 21644 13300 21700
rect 13580 21980 13636 22036
rect 13356 21756 13412 21812
rect 12796 21026 12852 21028
rect 12796 20974 12798 21026
rect 12798 20974 12850 21026
rect 12850 20974 12852 21026
rect 12796 20972 12852 20974
rect 12124 20188 12180 20244
rect 12796 20578 12852 20580
rect 12796 20526 12798 20578
rect 12798 20526 12850 20578
rect 12850 20526 12852 20578
rect 12796 20524 12852 20526
rect 12460 20130 12516 20132
rect 12460 20078 12462 20130
rect 12462 20078 12514 20130
rect 12514 20078 12516 20130
rect 12460 20076 12516 20078
rect 10892 18956 10948 19012
rect 10780 18844 10836 18900
rect 11116 18732 11172 18788
rect 14476 21756 14532 21812
rect 13468 21698 13524 21700
rect 13468 21646 13470 21698
rect 13470 21646 13522 21698
rect 13522 21646 13524 21698
rect 13468 21644 13524 21646
rect 13686 21194 13742 21196
rect 13686 21142 13688 21194
rect 13688 21142 13740 21194
rect 13740 21142 13742 21194
rect 13686 21140 13742 21142
rect 13790 21194 13846 21196
rect 13790 21142 13792 21194
rect 13792 21142 13844 21194
rect 13844 21142 13846 21194
rect 13790 21140 13846 21142
rect 13894 21194 13950 21196
rect 13894 21142 13896 21194
rect 13896 21142 13948 21194
rect 13948 21142 13950 21194
rect 13894 21140 13950 21142
rect 13580 20748 13636 20804
rect 13132 20076 13188 20132
rect 12572 19740 12628 19796
rect 12348 19292 12404 19348
rect 14140 20802 14196 20804
rect 14140 20750 14142 20802
rect 14142 20750 14194 20802
rect 14194 20750 14196 20802
rect 14140 20748 14196 20750
rect 14364 20748 14420 20804
rect 14364 20524 14420 20580
rect 13356 19292 13412 19348
rect 13580 20076 13636 20132
rect 11900 19010 11956 19012
rect 11900 18958 11902 19010
rect 11902 18958 11954 19010
rect 11954 18958 11956 19010
rect 11900 18956 11956 18958
rect 11228 18620 11284 18676
rect 11116 18172 11172 18228
rect 11788 18450 11844 18452
rect 11788 18398 11790 18450
rect 11790 18398 11842 18450
rect 11842 18398 11844 18450
rect 11788 18396 11844 18398
rect 12348 18338 12404 18340
rect 12348 18286 12350 18338
rect 12350 18286 12402 18338
rect 12402 18286 12404 18338
rect 12348 18284 12404 18286
rect 12796 18060 12852 18116
rect 11004 17724 11060 17780
rect 10668 17554 10724 17556
rect 10668 17502 10670 17554
rect 10670 17502 10722 17554
rect 10722 17502 10724 17554
rect 10668 17500 10724 17502
rect 11116 17442 11172 17444
rect 11116 17390 11118 17442
rect 11118 17390 11170 17442
rect 11170 17390 11172 17442
rect 11116 17388 11172 17390
rect 10556 17052 10612 17108
rect 11228 17052 11284 17108
rect 10444 16940 10500 16996
rect 8316 16716 8372 16772
rect 5068 15036 5124 15092
rect 2940 14252 2996 14308
rect 3724 14252 3780 14308
rect 4620 14252 4676 14308
rect 5740 15036 5796 15092
rect 5370 14922 5426 14924
rect 5370 14870 5372 14922
rect 5372 14870 5424 14922
rect 5424 14870 5426 14922
rect 5370 14868 5426 14870
rect 5474 14922 5530 14924
rect 5474 14870 5476 14922
rect 5476 14870 5528 14922
rect 5528 14870 5530 14922
rect 5474 14868 5530 14870
rect 5578 14922 5634 14924
rect 5578 14870 5580 14922
rect 5580 14870 5632 14922
rect 5632 14870 5634 14922
rect 5578 14868 5634 14870
rect 5628 14306 5684 14308
rect 5628 14254 5630 14306
rect 5630 14254 5682 14306
rect 5682 14254 5684 14306
rect 5628 14252 5684 14254
rect 5516 13746 5572 13748
rect 5516 13694 5518 13746
rect 5518 13694 5570 13746
rect 5570 13694 5572 13746
rect 5516 13692 5572 13694
rect 5964 14028 6020 14084
rect 5964 13858 6020 13860
rect 5964 13806 5966 13858
rect 5966 13806 6018 13858
rect 6018 13806 6020 13858
rect 5964 13804 6020 13806
rect 5068 13468 5124 13524
rect 5370 13354 5426 13356
rect 5370 13302 5372 13354
rect 5372 13302 5424 13354
rect 5424 13302 5426 13354
rect 5370 13300 5426 13302
rect 5474 13354 5530 13356
rect 5474 13302 5476 13354
rect 5476 13302 5528 13354
rect 5528 13302 5530 13354
rect 5474 13300 5530 13302
rect 5578 13354 5634 13356
rect 5578 13302 5580 13354
rect 5580 13302 5632 13354
rect 5632 13302 5634 13354
rect 5578 13300 5634 13302
rect 2492 11564 2548 11620
rect 2828 12572 2884 12628
rect 2156 11394 2212 11396
rect 2156 11342 2158 11394
rect 2158 11342 2210 11394
rect 2210 11342 2212 11394
rect 2156 11340 2212 11342
rect 2604 11170 2660 11172
rect 2604 11118 2606 11170
rect 2606 11118 2658 11170
rect 2658 11118 2660 11170
rect 2604 11116 2660 11118
rect 2716 10780 2772 10836
rect 2604 9884 2660 9940
rect 2492 8540 2548 8596
rect 2156 8316 2212 8372
rect 2716 9826 2772 9828
rect 2716 9774 2718 9826
rect 2718 9774 2770 9826
rect 2770 9774 2772 9826
rect 2716 9772 2772 9774
rect 3612 12738 3668 12740
rect 3612 12686 3614 12738
rect 3614 12686 3666 12738
rect 3666 12686 3668 12738
rect 3612 12684 3668 12686
rect 3500 11954 3556 11956
rect 3500 11902 3502 11954
rect 3502 11902 3554 11954
rect 3554 11902 3556 11954
rect 3500 11900 3556 11902
rect 3052 11506 3108 11508
rect 3052 11454 3054 11506
rect 3054 11454 3106 11506
rect 3106 11454 3108 11506
rect 3052 11452 3108 11454
rect 3276 10892 3332 10948
rect 2940 10668 2996 10724
rect 3276 10722 3332 10724
rect 3276 10670 3278 10722
rect 3278 10670 3330 10722
rect 3330 10670 3332 10722
rect 3276 10668 3332 10670
rect 2940 10498 2996 10500
rect 2940 10446 2942 10498
rect 2942 10446 2994 10498
rect 2994 10446 2996 10498
rect 2940 10444 2996 10446
rect 3052 9996 3108 10052
rect 3164 9938 3220 9940
rect 3164 9886 3166 9938
rect 3166 9886 3218 9938
rect 3218 9886 3220 9938
rect 3164 9884 3220 9886
rect 3836 12124 3892 12180
rect 4172 11788 4228 11844
rect 3724 11676 3780 11732
rect 10780 16828 10836 16884
rect 12236 16882 12292 16884
rect 12236 16830 12238 16882
rect 12238 16830 12290 16882
rect 12290 16830 12292 16882
rect 12236 16828 12292 16830
rect 11676 16716 11732 16772
rect 9528 15706 9584 15708
rect 9528 15654 9530 15706
rect 9530 15654 9582 15706
rect 9582 15654 9584 15706
rect 9528 15652 9584 15654
rect 9632 15706 9688 15708
rect 9632 15654 9634 15706
rect 9634 15654 9686 15706
rect 9686 15654 9688 15706
rect 9632 15652 9688 15654
rect 9736 15706 9792 15708
rect 9736 15654 9738 15706
rect 9738 15654 9790 15706
rect 9790 15654 9792 15706
rect 9736 15652 9792 15654
rect 6300 15036 6356 15092
rect 8988 15036 9044 15092
rect 11228 15314 11284 15316
rect 11228 15262 11230 15314
rect 11230 15262 11282 15314
rect 11282 15262 11284 15314
rect 11228 15260 11284 15262
rect 9996 15036 10052 15092
rect 7308 13858 7364 13860
rect 7308 13806 7310 13858
rect 7310 13806 7362 13858
rect 7362 13806 7364 13858
rect 7308 13804 7364 13806
rect 7644 13804 7700 13860
rect 4956 12908 5012 12964
rect 4620 12460 4676 12516
rect 4508 12178 4564 12180
rect 4508 12126 4510 12178
rect 4510 12126 4562 12178
rect 4562 12126 4564 12178
rect 4508 12124 4564 12126
rect 4396 11900 4452 11956
rect 3500 11394 3556 11396
rect 3500 11342 3502 11394
rect 3502 11342 3554 11394
rect 3554 11342 3556 11394
rect 3500 11340 3556 11342
rect 3612 11116 3668 11172
rect 3612 9996 3668 10052
rect 2940 9436 2996 9492
rect 3724 9602 3780 9604
rect 3724 9550 3726 9602
rect 3726 9550 3778 9602
rect 3778 9550 3780 9602
rect 3724 9548 3780 9550
rect 3500 9436 3556 9492
rect 4060 9826 4116 9828
rect 4060 9774 4062 9826
rect 4062 9774 4114 9826
rect 4114 9774 4116 9826
rect 4060 9772 4116 9774
rect 2268 7980 2324 8036
rect 2828 8146 2884 8148
rect 2828 8094 2830 8146
rect 2830 8094 2882 8146
rect 2882 8094 2884 8146
rect 2828 8092 2884 8094
rect 3388 8092 3444 8148
rect 3948 8988 4004 9044
rect 3612 8540 3668 8596
rect 2828 7196 2884 7252
rect 2604 7084 2660 7140
rect 2828 6972 2884 7028
rect 2604 5906 2660 5908
rect 2604 5854 2606 5906
rect 2606 5854 2658 5906
rect 2658 5854 2660 5906
rect 2604 5852 2660 5854
rect 3500 7532 3556 7588
rect 3612 7420 3668 7476
rect 3500 6860 3556 6916
rect 2940 6076 2996 6132
rect 3276 6130 3332 6132
rect 3276 6078 3278 6130
rect 3278 6078 3330 6130
rect 3330 6078 3332 6130
rect 3276 6076 3332 6078
rect 3052 5906 3108 5908
rect 3052 5854 3054 5906
rect 3054 5854 3106 5906
rect 3106 5854 3108 5906
rect 3052 5852 3108 5854
rect 2492 5122 2548 5124
rect 2492 5070 2494 5122
rect 2494 5070 2546 5122
rect 2546 5070 2548 5122
rect 2492 5068 2548 5070
rect 3836 8370 3892 8372
rect 3836 8318 3838 8370
rect 3838 8318 3890 8370
rect 3890 8318 3892 8370
rect 3836 8316 3892 8318
rect 4060 8764 4116 8820
rect 5852 12962 5908 12964
rect 5852 12910 5854 12962
rect 5854 12910 5906 12962
rect 5906 12910 5908 12962
rect 5852 12908 5908 12910
rect 5068 12348 5124 12404
rect 5404 12684 5460 12740
rect 5516 12460 5572 12516
rect 5852 12236 5908 12292
rect 5292 11900 5348 11956
rect 4956 11788 5012 11844
rect 4732 11340 4788 11396
rect 4844 11116 4900 11172
rect 4396 10556 4452 10612
rect 4732 10332 4788 10388
rect 4284 9436 4340 9492
rect 4620 9266 4676 9268
rect 4620 9214 4622 9266
rect 4622 9214 4674 9266
rect 4674 9214 4676 9266
rect 4620 9212 4676 9214
rect 4284 8876 4340 8932
rect 4396 8540 4452 8596
rect 4172 8316 4228 8372
rect 4060 7868 4116 7924
rect 3836 7756 3892 7812
rect 4396 8204 4452 8260
rect 4172 7644 4228 7700
rect 4284 8092 4340 8148
rect 4508 8034 4564 8036
rect 4508 7982 4510 8034
rect 4510 7982 4562 8034
rect 4562 7982 4564 8034
rect 4508 7980 4564 7982
rect 4508 7644 4564 7700
rect 5370 11786 5426 11788
rect 5370 11734 5372 11786
rect 5372 11734 5424 11786
rect 5424 11734 5426 11786
rect 5370 11732 5426 11734
rect 5474 11786 5530 11788
rect 5474 11734 5476 11786
rect 5476 11734 5528 11786
rect 5528 11734 5530 11786
rect 5474 11732 5530 11734
rect 5578 11786 5634 11788
rect 5578 11734 5580 11786
rect 5580 11734 5632 11786
rect 5632 11734 5634 11786
rect 5578 11732 5634 11734
rect 6076 12124 6132 12180
rect 6188 12908 6244 12964
rect 5516 11394 5572 11396
rect 5516 11342 5518 11394
rect 5518 11342 5570 11394
rect 5570 11342 5572 11394
rect 5516 11340 5572 11342
rect 5068 10610 5124 10612
rect 5068 10558 5070 10610
rect 5070 10558 5122 10610
rect 5122 10558 5124 10610
rect 5068 10556 5124 10558
rect 5516 10332 5572 10388
rect 5370 10218 5426 10220
rect 5370 10166 5372 10218
rect 5372 10166 5424 10218
rect 5424 10166 5426 10218
rect 5370 10164 5426 10166
rect 5474 10218 5530 10220
rect 5474 10166 5476 10218
rect 5476 10166 5528 10218
rect 5528 10166 5530 10218
rect 5474 10164 5530 10166
rect 5578 10218 5634 10220
rect 5578 10166 5580 10218
rect 5580 10166 5632 10218
rect 5632 10166 5634 10218
rect 5578 10164 5634 10166
rect 4956 9996 5012 10052
rect 5628 9884 5684 9940
rect 5964 11228 6020 11284
rect 6076 10668 6132 10724
rect 6748 13468 6804 13524
rect 6412 12236 6468 12292
rect 6524 12348 6580 12404
rect 6524 11564 6580 11620
rect 6300 11394 6356 11396
rect 6300 11342 6302 11394
rect 6302 11342 6354 11394
rect 6354 11342 6356 11394
rect 6300 11340 6356 11342
rect 7196 12572 7252 12628
rect 7868 13356 7924 13412
rect 7532 12850 7588 12852
rect 7532 12798 7534 12850
rect 7534 12798 7586 12850
rect 7586 12798 7588 12850
rect 7532 12796 7588 12798
rect 7308 12348 7364 12404
rect 9528 14138 9584 14140
rect 8428 13468 8484 13524
rect 8540 14028 8596 14084
rect 9528 14086 9530 14138
rect 9530 14086 9582 14138
rect 9582 14086 9584 14138
rect 9528 14084 9584 14086
rect 9632 14138 9688 14140
rect 9632 14086 9634 14138
rect 9634 14086 9686 14138
rect 9686 14086 9688 14138
rect 9632 14084 9688 14086
rect 9736 14138 9792 14140
rect 9736 14086 9738 14138
rect 9738 14086 9790 14138
rect 9790 14086 9792 14138
rect 9736 14084 9792 14086
rect 7084 11900 7140 11956
rect 6860 11618 6916 11620
rect 6860 11566 6862 11618
rect 6862 11566 6914 11618
rect 6914 11566 6916 11618
rect 6860 11564 6916 11566
rect 7084 11394 7140 11396
rect 7084 11342 7086 11394
rect 7086 11342 7138 11394
rect 7138 11342 7140 11394
rect 7084 11340 7140 11342
rect 6524 10780 6580 10836
rect 6300 10556 6356 10612
rect 4956 9548 5012 9604
rect 4844 8818 4900 8820
rect 4844 8766 4846 8818
rect 4846 8766 4898 8818
rect 4898 8766 4900 8818
rect 4844 8764 4900 8766
rect 4956 8428 5012 8484
rect 4172 7084 4228 7140
rect 4732 6972 4788 7028
rect 5852 9212 5908 9268
rect 5516 9154 5572 9156
rect 5516 9102 5518 9154
rect 5518 9102 5570 9154
rect 5570 9102 5572 9154
rect 5516 9100 5572 9102
rect 5370 8650 5426 8652
rect 5370 8598 5372 8650
rect 5372 8598 5424 8650
rect 5424 8598 5426 8650
rect 5370 8596 5426 8598
rect 5474 8650 5530 8652
rect 5474 8598 5476 8650
rect 5476 8598 5528 8650
rect 5528 8598 5530 8650
rect 5474 8596 5530 8598
rect 5578 8650 5634 8652
rect 5578 8598 5580 8650
rect 5580 8598 5632 8650
rect 5632 8598 5634 8650
rect 5578 8596 5634 8598
rect 5628 8428 5684 8484
rect 5964 8540 6020 8596
rect 6188 9714 6244 9716
rect 6188 9662 6190 9714
rect 6190 9662 6242 9714
rect 6242 9662 6244 9714
rect 6188 9660 6244 9662
rect 7084 10610 7140 10612
rect 7084 10558 7086 10610
rect 7086 10558 7138 10610
rect 7138 10558 7140 10610
rect 7084 10556 7140 10558
rect 5740 7980 5796 8036
rect 4844 7308 4900 7364
rect 4844 6860 4900 6916
rect 5292 7474 5348 7476
rect 5292 7422 5294 7474
rect 5294 7422 5346 7474
rect 5346 7422 5348 7474
rect 5292 7420 5348 7422
rect 5740 7756 5796 7812
rect 5370 7082 5426 7084
rect 5068 6972 5124 7028
rect 5370 7030 5372 7082
rect 5372 7030 5424 7082
rect 5424 7030 5426 7082
rect 5370 7028 5426 7030
rect 5474 7082 5530 7084
rect 5474 7030 5476 7082
rect 5476 7030 5528 7082
rect 5528 7030 5530 7082
rect 5474 7028 5530 7030
rect 5578 7082 5634 7084
rect 5578 7030 5580 7082
rect 5580 7030 5632 7082
rect 5632 7030 5634 7082
rect 5740 7084 5796 7140
rect 5578 7028 5634 7030
rect 5068 6748 5124 6804
rect 5180 6860 5236 6916
rect 3612 6412 3668 6468
rect 4620 6466 4676 6468
rect 4620 6414 4622 6466
rect 4622 6414 4674 6466
rect 4674 6414 4676 6466
rect 4620 6412 4676 6414
rect 5628 6802 5684 6804
rect 5628 6750 5630 6802
rect 5630 6750 5682 6802
rect 5682 6750 5684 6802
rect 5628 6748 5684 6750
rect 5740 6578 5796 6580
rect 5740 6526 5742 6578
rect 5742 6526 5794 6578
rect 5794 6526 5796 6578
rect 5740 6524 5796 6526
rect 3948 6300 4004 6356
rect 5292 5964 5348 6020
rect 4396 5906 4452 5908
rect 4396 5854 4398 5906
rect 4398 5854 4450 5906
rect 4450 5854 4452 5906
rect 4396 5852 4452 5854
rect 4060 5740 4116 5796
rect 4620 5346 4676 5348
rect 4620 5294 4622 5346
rect 4622 5294 4674 5346
rect 4674 5294 4676 5346
rect 4620 5292 4676 5294
rect 4284 5122 4340 5124
rect 4284 5070 4286 5122
rect 4286 5070 4338 5122
rect 4338 5070 4340 5122
rect 4284 5068 4340 5070
rect 6076 7644 6132 7700
rect 6524 9154 6580 9156
rect 6524 9102 6526 9154
rect 6526 9102 6578 9154
rect 6578 9102 6580 9154
rect 6524 9100 6580 9102
rect 6412 9042 6468 9044
rect 6412 8990 6414 9042
rect 6414 8990 6466 9042
rect 6466 8990 6468 9042
rect 6412 8988 6468 8990
rect 6636 8428 6692 8484
rect 6524 8258 6580 8260
rect 6524 8206 6526 8258
rect 6526 8206 6578 8258
rect 6578 8206 6580 8258
rect 6524 8204 6580 8206
rect 5964 5740 6020 5796
rect 6300 7868 6356 7924
rect 5852 5628 5908 5684
rect 7084 9772 7140 9828
rect 7084 9212 7140 9268
rect 7084 8764 7140 8820
rect 6972 8652 7028 8708
rect 7420 11282 7476 11284
rect 7420 11230 7422 11282
rect 7422 11230 7474 11282
rect 7474 11230 7476 11282
rect 7420 11228 7476 11230
rect 7308 10834 7364 10836
rect 7308 10782 7310 10834
rect 7310 10782 7362 10834
rect 7362 10782 7364 10834
rect 7308 10780 7364 10782
rect 7420 10108 7476 10164
rect 8316 12572 8372 12628
rect 8204 12066 8260 12068
rect 8204 12014 8206 12066
rect 8206 12014 8258 12066
rect 8258 12014 8260 12066
rect 8204 12012 8260 12014
rect 7644 10834 7700 10836
rect 7644 10782 7646 10834
rect 7646 10782 7698 10834
rect 7698 10782 7700 10834
rect 7644 10780 7700 10782
rect 7980 11340 8036 11396
rect 7532 9996 7588 10052
rect 8204 10556 8260 10612
rect 7308 9212 7364 9268
rect 7868 9772 7924 9828
rect 7756 9042 7812 9044
rect 7756 8990 7758 9042
rect 7758 8990 7810 9042
rect 7810 8990 7812 9042
rect 7756 8988 7812 8990
rect 7644 8652 7700 8708
rect 7980 8876 8036 8932
rect 6972 8316 7028 8372
rect 7196 8146 7252 8148
rect 7196 8094 7198 8146
rect 7198 8094 7250 8146
rect 7250 8094 7252 8146
rect 7196 8092 7252 8094
rect 7420 8092 7476 8148
rect 6860 7474 6916 7476
rect 6860 7422 6862 7474
rect 6862 7422 6914 7474
rect 6914 7422 6916 7474
rect 6860 7420 6916 7422
rect 7196 7868 7252 7924
rect 7308 7756 7364 7812
rect 6636 7084 6692 7140
rect 6188 6466 6244 6468
rect 6188 6414 6190 6466
rect 6190 6414 6242 6466
rect 6242 6414 6244 6466
rect 6188 6412 6244 6414
rect 6412 6412 6468 6468
rect 6524 6188 6580 6244
rect 6188 5964 6244 6020
rect 5370 5514 5426 5516
rect 5370 5462 5372 5514
rect 5372 5462 5424 5514
rect 5424 5462 5426 5514
rect 5370 5460 5426 5462
rect 5474 5514 5530 5516
rect 5474 5462 5476 5514
rect 5476 5462 5528 5514
rect 5528 5462 5530 5514
rect 5474 5460 5530 5462
rect 5578 5514 5634 5516
rect 5578 5462 5580 5514
rect 5580 5462 5632 5514
rect 5632 5462 5634 5514
rect 5578 5460 5634 5462
rect 5180 5292 5236 5348
rect 4844 5122 4900 5124
rect 4844 5070 4846 5122
rect 4846 5070 4898 5122
rect 4898 5070 4900 5122
rect 4844 5068 4900 5070
rect 5068 5180 5124 5236
rect 4732 4562 4788 4564
rect 4732 4510 4734 4562
rect 4734 4510 4786 4562
rect 4786 4510 4788 4562
rect 4732 4508 4788 4510
rect 3612 4396 3668 4452
rect 1820 4338 1876 4340
rect 1820 4286 1822 4338
rect 1822 4286 1874 4338
rect 1874 4286 1876 4338
rect 1820 4284 1876 4286
rect 1596 4172 1652 4228
rect 3612 4172 3668 4228
rect 6188 5180 6244 5236
rect 5964 5122 6020 5124
rect 5964 5070 5966 5122
rect 5966 5070 6018 5122
rect 6018 5070 6020 5122
rect 5964 5068 6020 5070
rect 5740 4284 5796 4340
rect 5370 3946 5426 3948
rect 5370 3894 5372 3946
rect 5372 3894 5424 3946
rect 5424 3894 5426 3946
rect 5370 3892 5426 3894
rect 5474 3946 5530 3948
rect 5474 3894 5476 3946
rect 5476 3894 5528 3946
rect 5528 3894 5530 3946
rect 5474 3892 5530 3894
rect 5578 3946 5634 3948
rect 5578 3894 5580 3946
rect 5580 3894 5632 3946
rect 5632 3894 5634 3946
rect 5578 3892 5634 3894
rect 5180 3612 5236 3668
rect 6076 4956 6132 5012
rect 6412 4060 6468 4116
rect 7084 6188 7140 6244
rect 6860 4956 6916 5012
rect 6972 4450 7028 4452
rect 6972 4398 6974 4450
rect 6974 4398 7026 4450
rect 7026 4398 7028 4450
rect 6972 4396 7028 4398
rect 6748 4284 6804 4340
rect 6860 4172 6916 4228
rect 6972 4060 7028 4116
rect 6748 3612 6804 3668
rect 7868 7474 7924 7476
rect 7868 7422 7870 7474
rect 7870 7422 7922 7474
rect 7922 7422 7924 7474
rect 7868 7420 7924 7422
rect 7308 5010 7364 5012
rect 7308 4958 7310 5010
rect 7310 4958 7362 5010
rect 7362 4958 7364 5010
rect 7308 4956 7364 4958
rect 7644 5906 7700 5908
rect 7644 5854 7646 5906
rect 7646 5854 7698 5906
rect 7698 5854 7700 5906
rect 7644 5852 7700 5854
rect 7868 6466 7924 6468
rect 7868 6414 7870 6466
rect 7870 6414 7922 6466
rect 7922 6414 7924 6466
rect 7868 6412 7924 6414
rect 9772 13970 9828 13972
rect 9772 13918 9774 13970
rect 9774 13918 9826 13970
rect 9826 13918 9828 13970
rect 9772 13916 9828 13918
rect 9548 13746 9604 13748
rect 9548 13694 9550 13746
rect 9550 13694 9602 13746
rect 9602 13694 9604 13746
rect 9548 13692 9604 13694
rect 9548 13468 9604 13524
rect 12908 16828 12964 16884
rect 12348 16716 12404 16772
rect 12796 16156 12852 16212
rect 14028 20130 14084 20132
rect 14028 20078 14030 20130
rect 14030 20078 14082 20130
rect 14082 20078 14084 20130
rect 14028 20076 14084 20078
rect 14252 20018 14308 20020
rect 14252 19966 14254 20018
rect 14254 19966 14306 20018
rect 14306 19966 14308 20018
rect 14252 19964 14308 19966
rect 15036 24108 15092 24164
rect 14924 23772 14980 23828
rect 14812 23436 14868 23492
rect 15036 23154 15092 23156
rect 15036 23102 15038 23154
rect 15038 23102 15090 23154
rect 15090 23102 15092 23154
rect 15036 23100 15092 23102
rect 14812 21698 14868 21700
rect 14812 21646 14814 21698
rect 14814 21646 14866 21698
rect 14866 21646 14868 21698
rect 14812 21644 14868 21646
rect 14700 21532 14756 21588
rect 15372 23548 15428 23604
rect 15372 23212 15428 23268
rect 17164 27186 17220 27188
rect 17164 27134 17166 27186
rect 17166 27134 17218 27186
rect 17218 27134 17220 27186
rect 17164 27132 17220 27134
rect 16380 26290 16436 26292
rect 16380 26238 16382 26290
rect 16382 26238 16434 26290
rect 16434 26238 16436 26290
rect 16380 26236 16436 26238
rect 16604 25788 16660 25844
rect 16156 25394 16212 25396
rect 16156 25342 16158 25394
rect 16158 25342 16210 25394
rect 16210 25342 16212 25394
rect 16156 25340 16212 25342
rect 17724 27020 17780 27076
rect 17724 26796 17780 26852
rect 17844 26682 17900 26684
rect 17844 26630 17846 26682
rect 17846 26630 17898 26682
rect 17898 26630 17900 26682
rect 17844 26628 17900 26630
rect 17948 26682 18004 26684
rect 17948 26630 17950 26682
rect 17950 26630 18002 26682
rect 18002 26630 18004 26682
rect 17948 26628 18004 26630
rect 18052 26682 18108 26684
rect 18052 26630 18054 26682
rect 18054 26630 18106 26682
rect 18106 26630 18108 26682
rect 18052 26628 18108 26630
rect 18956 26572 19012 26628
rect 17612 26124 17668 26180
rect 16268 25282 16324 25284
rect 16268 25230 16270 25282
rect 16270 25230 16322 25282
rect 16322 25230 16324 25282
rect 16268 25228 16324 25230
rect 16380 24892 16436 24948
rect 15596 23884 15652 23940
rect 15932 23772 15988 23828
rect 15820 23436 15876 23492
rect 17164 23826 17220 23828
rect 17164 23774 17166 23826
rect 17166 23774 17218 23826
rect 17218 23774 17220 23826
rect 17164 23772 17220 23774
rect 16044 23378 16100 23380
rect 16044 23326 16046 23378
rect 16046 23326 16098 23378
rect 16098 23326 16100 23378
rect 16044 23324 16100 23326
rect 15596 23100 15652 23156
rect 15372 21474 15428 21476
rect 15372 21422 15374 21474
rect 15374 21422 15426 21474
rect 15426 21422 15428 21474
rect 15372 21420 15428 21422
rect 15484 20972 15540 21028
rect 14812 19852 14868 19908
rect 13686 19626 13742 19628
rect 13686 19574 13688 19626
rect 13688 19574 13740 19626
rect 13740 19574 13742 19626
rect 13686 19572 13742 19574
rect 13790 19626 13846 19628
rect 13790 19574 13792 19626
rect 13792 19574 13844 19626
rect 13844 19574 13846 19626
rect 13790 19572 13846 19574
rect 13894 19626 13950 19628
rect 13894 19574 13896 19626
rect 13896 19574 13948 19626
rect 13948 19574 13950 19626
rect 13894 19572 13950 19574
rect 14588 19068 14644 19124
rect 14028 18450 14084 18452
rect 14028 18398 14030 18450
rect 14030 18398 14082 18450
rect 14082 18398 14084 18450
rect 14028 18396 14084 18398
rect 13686 18058 13742 18060
rect 13686 18006 13688 18058
rect 13688 18006 13740 18058
rect 13740 18006 13742 18058
rect 13686 18004 13742 18006
rect 13790 18058 13846 18060
rect 13790 18006 13792 18058
rect 13792 18006 13844 18058
rect 13844 18006 13846 18058
rect 13790 18004 13846 18006
rect 13894 18058 13950 18060
rect 13894 18006 13896 18058
rect 13896 18006 13948 18058
rect 13948 18006 13950 18058
rect 13894 18004 13950 18006
rect 14364 17500 14420 17556
rect 14140 16828 14196 16884
rect 14028 16770 14084 16772
rect 14028 16718 14030 16770
rect 14030 16718 14082 16770
rect 14082 16718 14084 16770
rect 14028 16716 14084 16718
rect 13916 16604 13972 16660
rect 13686 16490 13742 16492
rect 13686 16438 13688 16490
rect 13688 16438 13740 16490
rect 13740 16438 13742 16490
rect 13686 16436 13742 16438
rect 13790 16490 13846 16492
rect 13790 16438 13792 16490
rect 13792 16438 13844 16490
rect 13844 16438 13846 16490
rect 13790 16436 13846 16438
rect 13894 16490 13950 16492
rect 13894 16438 13896 16490
rect 13896 16438 13948 16490
rect 13948 16438 13950 16490
rect 13894 16436 13950 16438
rect 13692 16210 13748 16212
rect 13692 16158 13694 16210
rect 13694 16158 13746 16210
rect 13746 16158 13748 16210
rect 13692 16156 13748 16158
rect 14140 15986 14196 15988
rect 14140 15934 14142 15986
rect 14142 15934 14194 15986
rect 14194 15934 14196 15986
rect 14140 15932 14196 15934
rect 14028 15372 14084 15428
rect 13468 15260 13524 15316
rect 11676 13916 11732 13972
rect 12684 14364 12740 14420
rect 10108 13858 10164 13860
rect 10108 13806 10110 13858
rect 10110 13806 10162 13858
rect 10162 13806 10164 13858
rect 10108 13804 10164 13806
rect 11116 13858 11172 13860
rect 11116 13806 11118 13858
rect 11118 13806 11170 13858
rect 11170 13806 11172 13858
rect 11116 13804 11172 13806
rect 10892 13692 10948 13748
rect 9996 13580 10052 13636
rect 9772 13020 9828 13076
rect 10780 13580 10836 13636
rect 11900 13634 11956 13636
rect 11900 13582 11902 13634
rect 11902 13582 11954 13634
rect 11954 13582 11956 13634
rect 11900 13580 11956 13582
rect 12572 13356 12628 13412
rect 12124 13074 12180 13076
rect 12124 13022 12126 13074
rect 12126 13022 12178 13074
rect 12178 13022 12180 13074
rect 12124 13020 12180 13022
rect 8652 12572 8708 12628
rect 10108 12796 10164 12852
rect 9528 12570 9584 12572
rect 9528 12518 9530 12570
rect 9530 12518 9582 12570
rect 9582 12518 9584 12570
rect 9528 12516 9584 12518
rect 9632 12570 9688 12572
rect 9632 12518 9634 12570
rect 9634 12518 9686 12570
rect 9686 12518 9688 12570
rect 9632 12516 9688 12518
rect 9736 12570 9792 12572
rect 9736 12518 9738 12570
rect 9738 12518 9790 12570
rect 9790 12518 9792 12570
rect 9736 12516 9792 12518
rect 8988 12290 9044 12292
rect 8988 12238 8990 12290
rect 8990 12238 9042 12290
rect 9042 12238 9044 12290
rect 8988 12236 9044 12238
rect 10668 12290 10724 12292
rect 10668 12238 10670 12290
rect 10670 12238 10722 12290
rect 10722 12238 10724 12290
rect 10668 12236 10724 12238
rect 8540 11618 8596 11620
rect 8540 11566 8542 11618
rect 8542 11566 8594 11618
rect 8594 11566 8596 11618
rect 8540 11564 8596 11566
rect 9212 11452 9268 11508
rect 8876 10892 8932 10948
rect 8988 11228 9044 11284
rect 8876 10668 8932 10724
rect 8764 10332 8820 10388
rect 8764 9714 8820 9716
rect 8764 9662 8766 9714
rect 8766 9662 8818 9714
rect 8818 9662 8820 9714
rect 8764 9660 8820 9662
rect 8988 9548 9044 9604
rect 8988 9100 9044 9156
rect 8092 8428 8148 8484
rect 8092 8092 8148 8148
rect 7868 6130 7924 6132
rect 7868 6078 7870 6130
rect 7870 6078 7922 6130
rect 7922 6078 7924 6130
rect 7868 6076 7924 6078
rect 8764 8146 8820 8148
rect 8764 8094 8766 8146
rect 8766 8094 8818 8146
rect 8818 8094 8820 8146
rect 8764 8092 8820 8094
rect 8988 8428 9044 8484
rect 8876 7868 8932 7924
rect 8204 6524 8260 6580
rect 8204 6076 8260 6132
rect 8316 6412 8372 6468
rect 8204 5740 8260 5796
rect 8092 5628 8148 5684
rect 7980 5404 8036 5460
rect 7644 4898 7700 4900
rect 7644 4846 7646 4898
rect 7646 4846 7698 4898
rect 7698 4846 7700 4898
rect 7644 4844 7700 4846
rect 7644 4562 7700 4564
rect 7644 4510 7646 4562
rect 7646 4510 7698 4562
rect 7698 4510 7700 4562
rect 7644 4508 7700 4510
rect 8876 7420 8932 7476
rect 8428 6018 8484 6020
rect 8428 5966 8430 6018
rect 8430 5966 8482 6018
rect 8482 5966 8484 6018
rect 8428 5964 8484 5966
rect 8540 6188 8596 6244
rect 8540 5516 8596 5572
rect 8428 5292 8484 5348
rect 8204 4956 8260 5012
rect 7868 4060 7924 4116
rect 8764 5852 8820 5908
rect 8876 5740 8932 5796
rect 9324 11116 9380 11172
rect 9996 11116 10052 11172
rect 9528 11002 9584 11004
rect 9528 10950 9530 11002
rect 9530 10950 9582 11002
rect 9582 10950 9584 11002
rect 9528 10948 9584 10950
rect 9632 11002 9688 11004
rect 9632 10950 9634 11002
rect 9634 10950 9686 11002
rect 9686 10950 9688 11002
rect 9632 10948 9688 10950
rect 9736 11002 9792 11004
rect 9736 10950 9738 11002
rect 9738 10950 9790 11002
rect 9790 10950 9792 11002
rect 9736 10948 9792 10950
rect 9436 10610 9492 10612
rect 9436 10558 9438 10610
rect 9438 10558 9490 10610
rect 9490 10558 9492 10610
rect 9436 10556 9492 10558
rect 9884 10610 9940 10612
rect 9884 10558 9886 10610
rect 9886 10558 9938 10610
rect 9938 10558 9940 10610
rect 9884 10556 9940 10558
rect 10444 11564 10500 11620
rect 11340 12738 11396 12740
rect 11340 12686 11342 12738
rect 11342 12686 11394 12738
rect 11394 12686 11396 12738
rect 11340 12684 11396 12686
rect 12012 12738 12068 12740
rect 12012 12686 12014 12738
rect 12014 12686 12066 12738
rect 12066 12686 12068 12738
rect 12012 12684 12068 12686
rect 13132 13692 13188 13748
rect 13132 12684 13188 12740
rect 10892 11452 10948 11508
rect 10444 11394 10500 11396
rect 10444 11342 10446 11394
rect 10446 11342 10498 11394
rect 10498 11342 10500 11394
rect 10444 11340 10500 11342
rect 11340 11506 11396 11508
rect 11340 11454 11342 11506
rect 11342 11454 11394 11506
rect 11394 11454 11396 11506
rect 11340 11452 11396 11454
rect 11116 11282 11172 11284
rect 11116 11230 11118 11282
rect 11118 11230 11170 11282
rect 11170 11230 11172 11282
rect 11116 11228 11172 11230
rect 10444 11116 10500 11172
rect 11340 11170 11396 11172
rect 11340 11118 11342 11170
rect 11342 11118 11394 11170
rect 11394 11118 11396 11170
rect 11340 11116 11396 11118
rect 10220 10668 10276 10724
rect 11228 10780 11284 10836
rect 10220 10498 10276 10500
rect 10220 10446 10222 10498
rect 10222 10446 10274 10498
rect 10274 10446 10276 10498
rect 10220 10444 10276 10446
rect 9212 10050 9268 10052
rect 9212 9998 9214 10050
rect 9214 9998 9266 10050
rect 9266 9998 9268 10050
rect 9212 9996 9268 9998
rect 9548 9826 9604 9828
rect 9548 9774 9550 9826
rect 9550 9774 9602 9826
rect 9602 9774 9604 9826
rect 9548 9772 9604 9774
rect 9528 9434 9584 9436
rect 9528 9382 9530 9434
rect 9530 9382 9582 9434
rect 9582 9382 9584 9434
rect 9528 9380 9584 9382
rect 9632 9434 9688 9436
rect 9632 9382 9634 9434
rect 9634 9382 9686 9434
rect 9686 9382 9688 9434
rect 9632 9380 9688 9382
rect 9736 9434 9792 9436
rect 9736 9382 9738 9434
rect 9738 9382 9790 9434
rect 9790 9382 9792 9434
rect 9736 9380 9792 9382
rect 10556 9548 10612 9604
rect 9212 9100 9268 9156
rect 9996 9042 10052 9044
rect 9996 8990 9998 9042
rect 9998 8990 10050 9042
rect 10050 8990 10052 9042
rect 9996 8988 10052 8990
rect 10220 9100 10276 9156
rect 9548 8652 9604 8708
rect 9884 8258 9940 8260
rect 9884 8206 9886 8258
rect 9886 8206 9938 8258
rect 9938 8206 9940 8258
rect 9884 8204 9940 8206
rect 9548 7980 9604 8036
rect 9884 8034 9940 8036
rect 9884 7982 9886 8034
rect 9886 7982 9938 8034
rect 9938 7982 9940 8034
rect 9884 7980 9940 7982
rect 9528 7866 9584 7868
rect 9528 7814 9530 7866
rect 9530 7814 9582 7866
rect 9582 7814 9584 7866
rect 9528 7812 9584 7814
rect 9632 7866 9688 7868
rect 9632 7814 9634 7866
rect 9634 7814 9686 7866
rect 9686 7814 9688 7866
rect 9632 7812 9688 7814
rect 9736 7866 9792 7868
rect 9736 7814 9738 7866
rect 9738 7814 9790 7866
rect 9790 7814 9792 7866
rect 9736 7812 9792 7814
rect 9772 7644 9828 7700
rect 9436 7586 9492 7588
rect 9436 7534 9438 7586
rect 9438 7534 9490 7586
rect 9490 7534 9492 7586
rect 9436 7532 9492 7534
rect 10668 8540 10724 8596
rect 10108 8316 10164 8372
rect 10108 7532 10164 7588
rect 9660 6802 9716 6804
rect 9660 6750 9662 6802
rect 9662 6750 9714 6802
rect 9714 6750 9716 6802
rect 9660 6748 9716 6750
rect 9100 6636 9156 6692
rect 9884 7420 9940 7476
rect 9772 6690 9828 6692
rect 9772 6638 9774 6690
rect 9774 6638 9826 6690
rect 9826 6638 9828 6690
rect 9772 6636 9828 6638
rect 9884 7196 9940 7252
rect 9528 6298 9584 6300
rect 9528 6246 9530 6298
rect 9530 6246 9582 6298
rect 9582 6246 9584 6298
rect 9528 6244 9584 6246
rect 9632 6298 9688 6300
rect 9632 6246 9634 6298
rect 9634 6246 9686 6298
rect 9686 6246 9688 6298
rect 9632 6244 9688 6246
rect 9736 6298 9792 6300
rect 9736 6246 9738 6298
rect 9738 6246 9790 6298
rect 9790 6246 9792 6298
rect 9736 6244 9792 6246
rect 10444 7308 10500 7364
rect 9996 6524 10052 6580
rect 9324 5852 9380 5908
rect 8652 5180 8708 5236
rect 10556 7420 10612 7476
rect 10220 6524 10276 6580
rect 11004 10332 11060 10388
rect 10780 8316 10836 8372
rect 11452 9826 11508 9828
rect 11452 9774 11454 9826
rect 11454 9774 11506 9826
rect 11506 9774 11508 9826
rect 11452 9772 11508 9774
rect 13020 11564 13076 11620
rect 12348 10332 12404 10388
rect 12012 10220 12068 10276
rect 12908 10220 12964 10276
rect 12236 10108 12292 10164
rect 11564 8988 11620 9044
rect 11228 8652 11284 8708
rect 11116 7644 11172 7700
rect 11340 8204 11396 8260
rect 11676 8652 11732 8708
rect 11452 7420 11508 7476
rect 11004 6748 11060 6804
rect 11900 8428 11956 8484
rect 10780 6524 10836 6580
rect 9324 5628 9380 5684
rect 8876 5122 8932 5124
rect 8876 5070 8878 5122
rect 8878 5070 8930 5122
rect 8930 5070 8932 5122
rect 8876 5068 8932 5070
rect 8540 4956 8596 5012
rect 10108 5404 10164 5460
rect 10668 5516 10724 5572
rect 10220 5292 10276 5348
rect 10556 5404 10612 5460
rect 9528 4730 9584 4732
rect 9528 4678 9530 4730
rect 9530 4678 9582 4730
rect 9582 4678 9584 4730
rect 9528 4676 9584 4678
rect 9632 4730 9688 4732
rect 9632 4678 9634 4730
rect 9634 4678 9686 4730
rect 9686 4678 9688 4730
rect 9632 4676 9688 4678
rect 9736 4730 9792 4732
rect 9736 4678 9738 4730
rect 9738 4678 9790 4730
rect 9790 4678 9792 4730
rect 9736 4676 9792 4678
rect 8540 4508 8596 4564
rect 8988 4562 9044 4564
rect 8988 4510 8990 4562
rect 8990 4510 9042 4562
rect 9042 4510 9044 4562
rect 8988 4508 9044 4510
rect 11116 6188 11172 6244
rect 11116 6018 11172 6020
rect 11116 5966 11118 6018
rect 11118 5966 11170 6018
rect 11170 5966 11172 6018
rect 11116 5964 11172 5966
rect 11004 5068 11060 5124
rect 12124 8258 12180 8260
rect 12124 8206 12126 8258
rect 12126 8206 12178 8258
rect 12178 8206 12180 8258
rect 12124 8204 12180 8206
rect 11900 8092 11956 8148
rect 11900 7308 11956 7364
rect 12908 9826 12964 9828
rect 12908 9774 12910 9826
rect 12910 9774 12962 9826
rect 12962 9774 12964 9826
rect 12908 9772 12964 9774
rect 12460 8652 12516 8708
rect 13020 8988 13076 9044
rect 12236 7084 12292 7140
rect 12124 6748 12180 6804
rect 11788 6636 11844 6692
rect 11564 5682 11620 5684
rect 11564 5630 11566 5682
rect 11566 5630 11618 5682
rect 11618 5630 11620 5682
rect 11564 5628 11620 5630
rect 11452 5516 11508 5572
rect 12348 6524 12404 6580
rect 12684 7308 12740 7364
rect 12348 6300 12404 6356
rect 11228 4508 11284 4564
rect 11340 5068 11396 5124
rect 8764 4338 8820 4340
rect 8764 4286 8766 4338
rect 8766 4286 8818 4338
rect 8818 4286 8820 4338
rect 8764 4284 8820 4286
rect 10668 4284 10724 4340
rect 10220 4114 10276 4116
rect 10220 4062 10222 4114
rect 10222 4062 10274 4114
rect 10274 4062 10276 4114
rect 10220 4060 10276 4062
rect 9548 3554 9604 3556
rect 9548 3502 9550 3554
rect 9550 3502 9602 3554
rect 9602 3502 9604 3554
rect 9548 3500 9604 3502
rect 11788 5234 11844 5236
rect 11788 5182 11790 5234
rect 11790 5182 11842 5234
rect 11842 5182 11844 5234
rect 11788 5180 11844 5182
rect 11788 4956 11844 5012
rect 10780 3388 10836 3444
rect 8204 3276 8260 3332
rect 9528 3162 9584 3164
rect 9528 3110 9530 3162
rect 9530 3110 9582 3162
rect 9582 3110 9584 3162
rect 9528 3108 9584 3110
rect 9632 3162 9688 3164
rect 9632 3110 9634 3162
rect 9634 3110 9686 3162
rect 9686 3110 9688 3162
rect 9632 3108 9688 3110
rect 9736 3162 9792 3164
rect 9736 3110 9738 3162
rect 9738 3110 9790 3162
rect 9790 3110 9792 3162
rect 9736 3108 9792 3110
rect 6412 2940 6468 2996
rect 12124 5068 12180 5124
rect 12124 4508 12180 4564
rect 12796 7084 12852 7140
rect 12460 6018 12516 6020
rect 12460 5966 12462 6018
rect 12462 5966 12514 6018
rect 12514 5966 12516 6018
rect 12460 5964 12516 5966
rect 14700 18338 14756 18340
rect 14700 18286 14702 18338
rect 14702 18286 14754 18338
rect 14754 18286 14756 18338
rect 14700 18284 14756 18286
rect 15372 20130 15428 20132
rect 15372 20078 15374 20130
rect 15374 20078 15426 20130
rect 15426 20078 15428 20130
rect 15372 20076 15428 20078
rect 15036 19122 15092 19124
rect 15036 19070 15038 19122
rect 15038 19070 15090 19122
rect 15090 19070 15092 19122
rect 15036 19068 15092 19070
rect 15708 21810 15764 21812
rect 15708 21758 15710 21810
rect 15710 21758 15762 21810
rect 15762 21758 15764 21810
rect 15708 21756 15764 21758
rect 16380 21810 16436 21812
rect 16380 21758 16382 21810
rect 16382 21758 16434 21810
rect 16434 21758 16436 21810
rect 16380 21756 16436 21758
rect 16716 21756 16772 21812
rect 15932 21532 15988 21588
rect 15708 20018 15764 20020
rect 15708 19966 15710 20018
rect 15710 19966 15762 20018
rect 15762 19966 15764 20018
rect 15708 19964 15764 19966
rect 15596 18396 15652 18452
rect 15260 17106 15316 17108
rect 15260 17054 15262 17106
rect 15262 17054 15314 17106
rect 15314 17054 15316 17106
rect 15260 17052 15316 17054
rect 17500 25004 17556 25060
rect 18284 26290 18340 26292
rect 18284 26238 18286 26290
rect 18286 26238 18338 26290
rect 18338 26238 18340 26290
rect 18284 26236 18340 26238
rect 18620 25506 18676 25508
rect 18620 25454 18622 25506
rect 18622 25454 18674 25506
rect 18674 25454 18676 25506
rect 18620 25452 18676 25454
rect 17836 25228 17892 25284
rect 18172 25340 18228 25396
rect 17844 25114 17900 25116
rect 17844 25062 17846 25114
rect 17846 25062 17898 25114
rect 17898 25062 17900 25114
rect 17844 25060 17900 25062
rect 17948 25114 18004 25116
rect 17948 25062 17950 25114
rect 17950 25062 18002 25114
rect 18002 25062 18004 25114
rect 17948 25060 18004 25062
rect 18052 25114 18108 25116
rect 18052 25062 18054 25114
rect 18054 25062 18106 25114
rect 18106 25062 18108 25114
rect 18052 25060 18108 25062
rect 18844 26290 18900 26292
rect 18844 26238 18846 26290
rect 18846 26238 18898 26290
rect 18898 26238 18900 26290
rect 18844 26236 18900 26238
rect 18732 25340 18788 25396
rect 18620 25228 18676 25284
rect 19628 26124 19684 26180
rect 19292 25730 19348 25732
rect 19292 25678 19294 25730
rect 19294 25678 19346 25730
rect 19346 25678 19348 25730
rect 19292 25676 19348 25678
rect 20188 27858 20244 27860
rect 20188 27806 20190 27858
rect 20190 27806 20242 27858
rect 20242 27806 20244 27858
rect 20188 27804 20244 27806
rect 22002 27466 22058 27468
rect 22002 27414 22004 27466
rect 22004 27414 22056 27466
rect 22056 27414 22058 27466
rect 22002 27412 22058 27414
rect 22106 27466 22162 27468
rect 22106 27414 22108 27466
rect 22108 27414 22160 27466
rect 22160 27414 22162 27466
rect 22106 27412 22162 27414
rect 22210 27466 22266 27468
rect 22210 27414 22212 27466
rect 22212 27414 22264 27466
rect 22264 27414 22266 27466
rect 22210 27412 22266 27414
rect 30318 27466 30374 27468
rect 30318 27414 30320 27466
rect 30320 27414 30372 27466
rect 30372 27414 30374 27466
rect 30318 27412 30374 27414
rect 30422 27466 30478 27468
rect 30422 27414 30424 27466
rect 30424 27414 30476 27466
rect 30476 27414 30478 27466
rect 30422 27412 30478 27414
rect 30526 27466 30582 27468
rect 30526 27414 30528 27466
rect 30528 27414 30580 27466
rect 30580 27414 30582 27466
rect 30526 27412 30582 27414
rect 20524 26796 20580 26852
rect 20412 26572 20468 26628
rect 22652 26572 22708 26628
rect 22540 26178 22596 26180
rect 22540 26126 22542 26178
rect 22542 26126 22594 26178
rect 22594 26126 22596 26178
rect 22540 26124 22596 26126
rect 22002 25898 22058 25900
rect 22002 25846 22004 25898
rect 22004 25846 22056 25898
rect 22056 25846 22058 25898
rect 22002 25844 22058 25846
rect 22106 25898 22162 25900
rect 22106 25846 22108 25898
rect 22108 25846 22160 25898
rect 22160 25846 22162 25898
rect 22106 25844 22162 25846
rect 22210 25898 22266 25900
rect 22210 25846 22212 25898
rect 22212 25846 22264 25898
rect 22264 25846 22266 25898
rect 22210 25844 22266 25846
rect 20076 25506 20132 25508
rect 20076 25454 20078 25506
rect 20078 25454 20130 25506
rect 20130 25454 20132 25506
rect 20076 25452 20132 25454
rect 22540 25452 22596 25508
rect 19292 25228 19348 25284
rect 17612 23212 17668 23268
rect 17388 22540 17444 22596
rect 17500 22370 17556 22372
rect 17500 22318 17502 22370
rect 17502 22318 17554 22370
rect 17554 22318 17556 22370
rect 17500 22316 17556 22318
rect 17844 23546 17900 23548
rect 17844 23494 17846 23546
rect 17846 23494 17898 23546
rect 17898 23494 17900 23546
rect 17844 23492 17900 23494
rect 17948 23546 18004 23548
rect 17948 23494 17950 23546
rect 17950 23494 18002 23546
rect 18002 23494 18004 23546
rect 17948 23492 18004 23494
rect 18052 23546 18108 23548
rect 18052 23494 18054 23546
rect 18054 23494 18106 23546
rect 18106 23494 18108 23546
rect 18052 23492 18108 23494
rect 17724 23100 17780 23156
rect 17948 23042 18004 23044
rect 17948 22990 17950 23042
rect 17950 22990 18002 23042
rect 18002 22990 18004 23042
rect 17948 22988 18004 22990
rect 17844 21978 17900 21980
rect 17844 21926 17846 21978
rect 17846 21926 17898 21978
rect 17898 21926 17900 21978
rect 17844 21924 17900 21926
rect 17948 21978 18004 21980
rect 17948 21926 17950 21978
rect 17950 21926 18002 21978
rect 18002 21926 18004 21978
rect 17948 21924 18004 21926
rect 18052 21978 18108 21980
rect 18052 21926 18054 21978
rect 18054 21926 18106 21978
rect 18106 21926 18108 21978
rect 18052 21924 18108 21926
rect 18284 21644 18340 21700
rect 18732 24892 18788 24948
rect 18620 23324 18676 23380
rect 18844 23772 18900 23828
rect 19852 25394 19908 25396
rect 19852 25342 19854 25394
rect 19854 25342 19906 25394
rect 19906 25342 19908 25394
rect 19852 25340 19908 25342
rect 20300 25282 20356 25284
rect 20300 25230 20302 25282
rect 20302 25230 20354 25282
rect 20354 25230 20356 25282
rect 20300 25228 20356 25230
rect 19516 24556 19572 24612
rect 19516 23826 19572 23828
rect 19516 23774 19518 23826
rect 19518 23774 19570 23826
rect 19570 23774 19572 23826
rect 19516 23772 19572 23774
rect 18956 23324 19012 23380
rect 19628 23324 19684 23380
rect 19068 23266 19124 23268
rect 19068 23214 19070 23266
rect 19070 23214 19122 23266
rect 19122 23214 19124 23266
rect 19068 23212 19124 23214
rect 18396 22988 18452 23044
rect 19292 22988 19348 23044
rect 19628 22876 19684 22932
rect 18956 21756 19012 21812
rect 19404 21810 19460 21812
rect 19404 21758 19406 21810
rect 19406 21758 19458 21810
rect 19458 21758 19460 21810
rect 19404 21756 19460 21758
rect 19292 21698 19348 21700
rect 19292 21646 19294 21698
rect 19294 21646 19346 21698
rect 19346 21646 19348 21698
rect 19292 21644 19348 21646
rect 19628 22258 19684 22260
rect 19628 22206 19630 22258
rect 19630 22206 19682 22258
rect 19682 22206 19684 22258
rect 19628 22204 19684 22206
rect 20300 24050 20356 24052
rect 20300 23998 20302 24050
rect 20302 23998 20354 24050
rect 20354 23998 20356 24050
rect 20300 23996 20356 23998
rect 20412 23212 20468 23268
rect 19628 21756 19684 21812
rect 19852 22316 19908 22372
rect 20076 22370 20132 22372
rect 20076 22318 20078 22370
rect 20078 22318 20130 22370
rect 20130 22318 20132 22370
rect 20076 22316 20132 22318
rect 20188 22204 20244 22260
rect 16716 20860 16772 20916
rect 16044 20802 16100 20804
rect 16044 20750 16046 20802
rect 16046 20750 16098 20802
rect 16098 20750 16100 20802
rect 16044 20748 16100 20750
rect 17164 20636 17220 20692
rect 16156 19906 16212 19908
rect 16156 19854 16158 19906
rect 16158 19854 16210 19906
rect 16210 19854 16212 19906
rect 16156 19852 16212 19854
rect 16044 18284 16100 18340
rect 16604 20076 16660 20132
rect 16380 19852 16436 19908
rect 16828 19628 16884 19684
rect 16940 18956 16996 19012
rect 16828 18508 16884 18564
rect 16492 18284 16548 18340
rect 16156 17500 16212 17556
rect 14924 16716 14980 16772
rect 15932 16994 15988 16996
rect 15932 16942 15934 16994
rect 15934 16942 15986 16994
rect 15986 16942 15988 16994
rect 15932 16940 15988 16942
rect 14924 16044 14980 16100
rect 14812 15986 14868 15988
rect 14812 15934 14814 15986
rect 14814 15934 14866 15986
rect 14866 15934 14868 15986
rect 14812 15932 14868 15934
rect 15260 16658 15316 16660
rect 15260 16606 15262 16658
rect 15262 16606 15314 16658
rect 15314 16606 15316 16658
rect 15260 16604 15316 16606
rect 15260 15932 15316 15988
rect 15148 15708 15204 15764
rect 14812 15314 14868 15316
rect 14812 15262 14814 15314
rect 14814 15262 14866 15314
rect 14866 15262 14868 15314
rect 14812 15260 14868 15262
rect 15260 15372 15316 15428
rect 15596 16716 15652 16772
rect 15484 16098 15540 16100
rect 15484 16046 15486 16098
rect 15486 16046 15538 16098
rect 15538 16046 15540 16098
rect 15484 16044 15540 16046
rect 15708 15708 15764 15764
rect 15484 15538 15540 15540
rect 15484 15486 15486 15538
rect 15486 15486 15538 15538
rect 15538 15486 15540 15538
rect 15484 15484 15540 15486
rect 16716 16994 16772 16996
rect 16716 16942 16718 16994
rect 16718 16942 16770 16994
rect 16770 16942 16772 16994
rect 16716 16940 16772 16942
rect 16156 16098 16212 16100
rect 16156 16046 16158 16098
rect 16158 16046 16210 16098
rect 16210 16046 16212 16098
rect 16156 16044 16212 16046
rect 16044 15986 16100 15988
rect 16044 15934 16046 15986
rect 16046 15934 16098 15986
rect 16098 15934 16100 15986
rect 16044 15932 16100 15934
rect 15708 15260 15764 15316
rect 13686 14922 13742 14924
rect 13686 14870 13688 14922
rect 13688 14870 13740 14922
rect 13740 14870 13742 14922
rect 13686 14868 13742 14870
rect 13790 14922 13846 14924
rect 13790 14870 13792 14922
rect 13792 14870 13844 14922
rect 13844 14870 13846 14922
rect 13790 14868 13846 14870
rect 13894 14922 13950 14924
rect 13894 14870 13896 14922
rect 13896 14870 13948 14922
rect 13948 14870 13950 14922
rect 13894 14868 13950 14870
rect 13580 14418 13636 14420
rect 13580 14366 13582 14418
rect 13582 14366 13634 14418
rect 13634 14366 13636 14418
rect 13580 14364 13636 14366
rect 14140 13970 14196 13972
rect 14140 13918 14142 13970
rect 14142 13918 14194 13970
rect 14194 13918 14196 13970
rect 14140 13916 14196 13918
rect 13686 13354 13742 13356
rect 13686 13302 13688 13354
rect 13688 13302 13740 13354
rect 13740 13302 13742 13354
rect 13686 13300 13742 13302
rect 13790 13354 13846 13356
rect 13790 13302 13792 13354
rect 13792 13302 13844 13354
rect 13844 13302 13846 13354
rect 13790 13300 13846 13302
rect 13894 13354 13950 13356
rect 13894 13302 13896 13354
rect 13896 13302 13948 13354
rect 13948 13302 13950 13354
rect 13894 13300 13950 13302
rect 13804 12738 13860 12740
rect 13804 12686 13806 12738
rect 13806 12686 13858 12738
rect 13858 12686 13860 12738
rect 13804 12684 13860 12686
rect 13686 11786 13742 11788
rect 13686 11734 13688 11786
rect 13688 11734 13740 11786
rect 13740 11734 13742 11786
rect 13686 11732 13742 11734
rect 13790 11786 13846 11788
rect 13790 11734 13792 11786
rect 13792 11734 13844 11786
rect 13844 11734 13846 11786
rect 13790 11732 13846 11734
rect 13894 11786 13950 11788
rect 13894 11734 13896 11786
rect 13896 11734 13948 11786
rect 13948 11734 13950 11786
rect 13894 11732 13950 11734
rect 14252 11506 14308 11508
rect 14252 11454 14254 11506
rect 14254 11454 14306 11506
rect 14306 11454 14308 11506
rect 14252 11452 14308 11454
rect 13468 10332 13524 10388
rect 13686 10218 13742 10220
rect 13686 10166 13688 10218
rect 13688 10166 13740 10218
rect 13740 10166 13742 10218
rect 13686 10164 13742 10166
rect 13790 10218 13846 10220
rect 13790 10166 13792 10218
rect 13792 10166 13844 10218
rect 13844 10166 13846 10218
rect 13790 10164 13846 10166
rect 13894 10218 13950 10220
rect 13894 10166 13896 10218
rect 13896 10166 13948 10218
rect 13948 10166 13950 10218
rect 13894 10164 13950 10166
rect 13692 9996 13748 10052
rect 13580 9602 13636 9604
rect 13580 9550 13582 9602
rect 13582 9550 13634 9602
rect 13634 9550 13636 9602
rect 13580 9548 13636 9550
rect 13132 7868 13188 7924
rect 14140 9548 14196 9604
rect 13804 9042 13860 9044
rect 13804 8990 13806 9042
rect 13806 8990 13858 9042
rect 13858 8990 13860 9042
rect 13804 8988 13860 8990
rect 14140 8988 14196 9044
rect 13468 8540 13524 8596
rect 13686 8650 13742 8652
rect 13686 8598 13688 8650
rect 13688 8598 13740 8650
rect 13740 8598 13742 8650
rect 13686 8596 13742 8598
rect 13790 8650 13846 8652
rect 13790 8598 13792 8650
rect 13792 8598 13844 8650
rect 13844 8598 13846 8650
rect 13790 8596 13846 8598
rect 13894 8650 13950 8652
rect 13894 8598 13896 8650
rect 13896 8598 13948 8650
rect 13948 8598 13950 8650
rect 13894 8596 13950 8598
rect 13356 8428 13412 8484
rect 13804 8428 13860 8484
rect 13468 8258 13524 8260
rect 13468 8206 13470 8258
rect 13470 8206 13522 8258
rect 13522 8206 13524 8258
rect 13468 8204 13524 8206
rect 13468 7868 13524 7924
rect 13132 6636 13188 6692
rect 12796 5852 12852 5908
rect 13686 7082 13742 7084
rect 13686 7030 13688 7082
rect 13688 7030 13740 7082
rect 13740 7030 13742 7082
rect 13686 7028 13742 7030
rect 13790 7082 13846 7084
rect 13790 7030 13792 7082
rect 13792 7030 13844 7082
rect 13844 7030 13846 7082
rect 13790 7028 13846 7030
rect 13894 7082 13950 7084
rect 13894 7030 13896 7082
rect 13896 7030 13948 7082
rect 13948 7030 13950 7082
rect 13894 7028 13950 7030
rect 13804 6300 13860 6356
rect 13580 6130 13636 6132
rect 13580 6078 13582 6130
rect 13582 6078 13634 6130
rect 13634 6078 13636 6130
rect 13580 6076 13636 6078
rect 13692 6018 13748 6020
rect 13692 5966 13694 6018
rect 13694 5966 13746 6018
rect 13746 5966 13748 6018
rect 13692 5964 13748 5966
rect 12460 5180 12516 5236
rect 12684 5122 12740 5124
rect 12684 5070 12686 5122
rect 12686 5070 12738 5122
rect 12738 5070 12740 5122
rect 12684 5068 12740 5070
rect 13686 5514 13742 5516
rect 13686 5462 13688 5514
rect 13688 5462 13740 5514
rect 13740 5462 13742 5514
rect 13686 5460 13742 5462
rect 13790 5514 13846 5516
rect 13790 5462 13792 5514
rect 13792 5462 13844 5514
rect 13844 5462 13846 5514
rect 13790 5460 13846 5462
rect 13894 5514 13950 5516
rect 13894 5462 13896 5514
rect 13896 5462 13948 5514
rect 13948 5462 13950 5514
rect 13894 5460 13950 5462
rect 13692 5292 13748 5348
rect 13132 5068 13188 5124
rect 13356 4956 13412 5012
rect 13580 4898 13636 4900
rect 13580 4846 13582 4898
rect 13582 4846 13634 4898
rect 13634 4846 13636 4898
rect 13580 4844 13636 4846
rect 13468 4508 13524 4564
rect 12572 4338 12628 4340
rect 12572 4286 12574 4338
rect 12574 4286 12626 4338
rect 12626 4286 12628 4338
rect 12572 4284 12628 4286
rect 13916 5122 13972 5124
rect 13916 5070 13918 5122
rect 13918 5070 13970 5122
rect 13970 5070 13972 5122
rect 13916 5068 13972 5070
rect 16380 15090 16436 15092
rect 16380 15038 16382 15090
rect 16382 15038 16434 15090
rect 16434 15038 16436 15090
rect 16380 15036 16436 15038
rect 16492 14924 16548 14980
rect 17052 17778 17108 17780
rect 17052 17726 17054 17778
rect 17054 17726 17106 17778
rect 17106 17726 17108 17778
rect 17052 17724 17108 17726
rect 16716 16658 16772 16660
rect 16716 16606 16718 16658
rect 16718 16606 16770 16658
rect 16770 16606 16772 16658
rect 16716 16604 16772 16606
rect 16940 16268 16996 16324
rect 16716 16044 16772 16100
rect 16940 15986 16996 15988
rect 16940 15934 16942 15986
rect 16942 15934 16994 15986
rect 16994 15934 16996 15986
rect 16940 15932 16996 15934
rect 16828 15708 16884 15764
rect 16828 15426 16884 15428
rect 16828 15374 16830 15426
rect 16830 15374 16882 15426
rect 16882 15374 16884 15426
rect 16828 15372 16884 15374
rect 16940 15036 16996 15092
rect 16716 14924 16772 14980
rect 16940 14530 16996 14532
rect 16940 14478 16942 14530
rect 16942 14478 16994 14530
rect 16994 14478 16996 14530
rect 16940 14476 16996 14478
rect 16268 13916 16324 13972
rect 15708 12796 15764 12852
rect 15820 13132 15876 13188
rect 14588 8988 14644 9044
rect 14700 10332 14756 10388
rect 14924 9996 14980 10052
rect 14924 8988 14980 9044
rect 14700 8204 14756 8260
rect 14476 7362 14532 7364
rect 14476 7310 14478 7362
rect 14478 7310 14530 7362
rect 14530 7310 14532 7362
rect 14476 7308 14532 7310
rect 14140 6188 14196 6244
rect 14924 8540 14980 8596
rect 16044 12962 16100 12964
rect 16044 12910 16046 12962
rect 16046 12910 16098 12962
rect 16098 12910 16100 12962
rect 16044 12908 16100 12910
rect 17388 20860 17444 20916
rect 17276 19964 17332 20020
rect 17612 20636 17668 20692
rect 17724 20524 17780 20580
rect 17844 20410 17900 20412
rect 17844 20358 17846 20410
rect 17846 20358 17898 20410
rect 17898 20358 17900 20410
rect 17844 20356 17900 20358
rect 17948 20410 18004 20412
rect 17948 20358 17950 20410
rect 17950 20358 18002 20410
rect 18002 20358 18004 20410
rect 17948 20356 18004 20358
rect 18052 20410 18108 20412
rect 18052 20358 18054 20410
rect 18054 20358 18106 20410
rect 18106 20358 18108 20410
rect 18052 20356 18108 20358
rect 18396 20578 18452 20580
rect 18396 20526 18398 20578
rect 18398 20526 18450 20578
rect 18450 20526 18452 20578
rect 18396 20524 18452 20526
rect 17948 20076 18004 20132
rect 18172 20018 18228 20020
rect 18172 19966 18174 20018
rect 18174 19966 18226 20018
rect 18226 19966 18228 20018
rect 18172 19964 18228 19966
rect 18284 19852 18340 19908
rect 18060 19740 18116 19796
rect 18620 20018 18676 20020
rect 18620 19966 18622 20018
rect 18622 19966 18674 20018
rect 18674 19966 18676 20018
rect 18620 19964 18676 19966
rect 18956 19740 19012 19796
rect 17276 19068 17332 19124
rect 17388 19346 17444 19348
rect 17388 19294 17390 19346
rect 17390 19294 17442 19346
rect 17442 19294 17444 19346
rect 17388 19292 17444 19294
rect 18396 19346 18452 19348
rect 18396 19294 18398 19346
rect 18398 19294 18450 19346
rect 18450 19294 18452 19346
rect 18396 19292 18452 19294
rect 17388 18956 17444 19012
rect 17500 18508 17556 18564
rect 17500 18338 17556 18340
rect 17500 18286 17502 18338
rect 17502 18286 17554 18338
rect 17554 18286 17556 18338
rect 17500 18284 17556 18286
rect 17276 17052 17332 17108
rect 17388 17500 17444 17556
rect 17844 18842 17900 18844
rect 17844 18790 17846 18842
rect 17846 18790 17898 18842
rect 17898 18790 17900 18842
rect 17844 18788 17900 18790
rect 17948 18842 18004 18844
rect 17948 18790 17950 18842
rect 17950 18790 18002 18842
rect 18002 18790 18004 18842
rect 17948 18788 18004 18790
rect 18052 18842 18108 18844
rect 18052 18790 18054 18842
rect 18054 18790 18106 18842
rect 18106 18790 18108 18842
rect 18052 18788 18108 18790
rect 17948 18172 18004 18228
rect 18172 17554 18228 17556
rect 18172 17502 18174 17554
rect 18174 17502 18226 17554
rect 18226 17502 18228 17554
rect 18172 17500 18228 17502
rect 17836 17442 17892 17444
rect 17836 17390 17838 17442
rect 17838 17390 17890 17442
rect 17890 17390 17892 17442
rect 17836 17388 17892 17390
rect 17844 17274 17900 17276
rect 17844 17222 17846 17274
rect 17846 17222 17898 17274
rect 17898 17222 17900 17274
rect 17844 17220 17900 17222
rect 17948 17274 18004 17276
rect 17948 17222 17950 17274
rect 17950 17222 18002 17274
rect 18002 17222 18004 17274
rect 17948 17220 18004 17222
rect 18052 17274 18108 17276
rect 18052 17222 18054 17274
rect 18054 17222 18106 17274
rect 18106 17222 18108 17274
rect 18052 17220 18108 17222
rect 18172 17052 18228 17108
rect 17836 16940 17892 16996
rect 17612 16716 17668 16772
rect 17612 16044 17668 16100
rect 17948 16828 18004 16884
rect 17948 16322 18004 16324
rect 17948 16270 17950 16322
rect 17950 16270 18002 16322
rect 18002 16270 18004 16322
rect 17948 16268 18004 16270
rect 18284 15874 18340 15876
rect 18284 15822 18286 15874
rect 18286 15822 18338 15874
rect 18338 15822 18340 15874
rect 18284 15820 18340 15822
rect 17844 15706 17900 15708
rect 17844 15654 17846 15706
rect 17846 15654 17898 15706
rect 17898 15654 17900 15706
rect 17844 15652 17900 15654
rect 17948 15706 18004 15708
rect 17948 15654 17950 15706
rect 17950 15654 18002 15706
rect 18002 15654 18004 15706
rect 17948 15652 18004 15654
rect 18052 15706 18108 15708
rect 18052 15654 18054 15706
rect 18054 15654 18106 15706
rect 18106 15654 18108 15706
rect 18052 15652 18108 15654
rect 17948 15148 18004 15204
rect 19628 19964 19684 20020
rect 19180 19852 19236 19908
rect 18956 18620 19012 18676
rect 18508 18396 18564 18452
rect 18508 17442 18564 17444
rect 18508 17390 18510 17442
rect 18510 17390 18562 17442
rect 18562 17390 18564 17442
rect 18508 17388 18564 17390
rect 18508 17164 18564 17220
rect 19068 17442 19124 17444
rect 19068 17390 19070 17442
rect 19070 17390 19122 17442
rect 19122 17390 19124 17442
rect 19068 17388 19124 17390
rect 18956 17052 19012 17108
rect 19628 17164 19684 17220
rect 18508 16770 18564 16772
rect 18508 16718 18510 16770
rect 18510 16718 18562 16770
rect 18562 16718 18564 16770
rect 18508 16716 18564 16718
rect 19292 16604 19348 16660
rect 18732 15986 18788 15988
rect 18732 15934 18734 15986
rect 18734 15934 18786 15986
rect 18786 15934 18788 15986
rect 18732 15932 18788 15934
rect 19068 15874 19124 15876
rect 19068 15822 19070 15874
rect 19070 15822 19122 15874
rect 19122 15822 19124 15874
rect 19068 15820 19124 15822
rect 18732 15260 18788 15316
rect 17276 14530 17332 14532
rect 17276 14478 17278 14530
rect 17278 14478 17330 14530
rect 17330 14478 17332 14530
rect 17276 14476 17332 14478
rect 17388 14252 17444 14308
rect 16604 13468 16660 13524
rect 16268 12738 16324 12740
rect 16268 12686 16270 12738
rect 16270 12686 16322 12738
rect 16322 12686 16324 12738
rect 16268 12684 16324 12686
rect 16044 8764 16100 8820
rect 15708 8428 15764 8484
rect 15036 8092 15092 8148
rect 15372 7868 15428 7924
rect 14700 5964 14756 6020
rect 14812 6188 14868 6244
rect 14252 5852 14308 5908
rect 14588 5906 14644 5908
rect 14588 5854 14590 5906
rect 14590 5854 14642 5906
rect 14642 5854 14644 5906
rect 14588 5852 14644 5854
rect 14812 5852 14868 5908
rect 13686 3946 13742 3948
rect 13686 3894 13688 3946
rect 13688 3894 13740 3946
rect 13740 3894 13742 3946
rect 13686 3892 13742 3894
rect 13790 3946 13846 3948
rect 13790 3894 13792 3946
rect 13792 3894 13844 3946
rect 13844 3894 13846 3946
rect 13790 3892 13846 3894
rect 13894 3946 13950 3948
rect 13894 3894 13896 3946
rect 13896 3894 13948 3946
rect 13948 3894 13950 3946
rect 13894 3892 13950 3894
rect 14140 3778 14196 3780
rect 14140 3726 14142 3778
rect 14142 3726 14194 3778
rect 14194 3726 14196 3778
rect 14140 3724 14196 3726
rect 14476 4844 14532 4900
rect 14924 4396 14980 4452
rect 15484 6076 15540 6132
rect 15036 4284 15092 4340
rect 15260 3778 15316 3780
rect 15260 3726 15262 3778
rect 15262 3726 15314 3778
rect 15314 3726 15316 3778
rect 15260 3724 15316 3726
rect 16828 12908 16884 12964
rect 16940 12684 16996 12740
rect 16604 8876 16660 8932
rect 16044 6188 16100 6244
rect 17388 12850 17444 12852
rect 17388 12798 17390 12850
rect 17390 12798 17442 12850
rect 17442 12798 17444 12850
rect 17388 12796 17444 12798
rect 17844 14138 17900 14140
rect 17844 14086 17846 14138
rect 17846 14086 17898 14138
rect 17898 14086 17900 14138
rect 17844 14084 17900 14086
rect 17948 14138 18004 14140
rect 17948 14086 17950 14138
rect 17950 14086 18002 14138
rect 18002 14086 18004 14138
rect 17948 14084 18004 14086
rect 18052 14138 18108 14140
rect 18052 14086 18054 14138
rect 18054 14086 18106 14138
rect 18106 14086 18108 14138
rect 18052 14084 18108 14086
rect 17724 13858 17780 13860
rect 17724 13806 17726 13858
rect 17726 13806 17778 13858
rect 17778 13806 17780 13858
rect 17724 13804 17780 13806
rect 18956 15484 19012 15540
rect 19068 15372 19124 15428
rect 19180 14364 19236 14420
rect 18844 14252 18900 14308
rect 18396 13970 18452 13972
rect 18396 13918 18398 13970
rect 18398 13918 18450 13970
rect 18450 13918 18452 13970
rect 18396 13916 18452 13918
rect 18732 13692 18788 13748
rect 17276 11618 17332 11620
rect 17276 11566 17278 11618
rect 17278 11566 17330 11618
rect 17330 11566 17332 11618
rect 17276 11564 17332 11566
rect 17612 12236 17668 12292
rect 18172 12684 18228 12740
rect 17844 12570 17900 12572
rect 17844 12518 17846 12570
rect 17846 12518 17898 12570
rect 17898 12518 17900 12570
rect 17844 12516 17900 12518
rect 17948 12570 18004 12572
rect 17948 12518 17950 12570
rect 17950 12518 18002 12570
rect 18002 12518 18004 12570
rect 17948 12516 18004 12518
rect 18052 12570 18108 12572
rect 18052 12518 18054 12570
rect 18054 12518 18106 12570
rect 18106 12518 18108 12570
rect 18052 12516 18108 12518
rect 18284 12236 18340 12292
rect 18396 12908 18452 12964
rect 18956 13468 19012 13524
rect 18508 12348 18564 12404
rect 18172 11564 18228 11620
rect 17500 11228 17556 11284
rect 17844 11002 17900 11004
rect 17844 10950 17846 11002
rect 17846 10950 17898 11002
rect 17898 10950 17900 11002
rect 17844 10948 17900 10950
rect 17948 11002 18004 11004
rect 17948 10950 17950 11002
rect 17950 10950 18002 11002
rect 18002 10950 18004 11002
rect 17948 10948 18004 10950
rect 18052 11002 18108 11004
rect 18052 10950 18054 11002
rect 18054 10950 18106 11002
rect 18106 10950 18108 11002
rect 18052 10948 18108 10950
rect 16828 9772 16884 9828
rect 17836 9826 17892 9828
rect 17836 9774 17838 9826
rect 17838 9774 17890 9826
rect 17890 9774 17892 9826
rect 17836 9772 17892 9774
rect 18508 11228 18564 11284
rect 18508 10108 18564 10164
rect 17612 9660 17668 9716
rect 17844 9434 17900 9436
rect 17844 9382 17846 9434
rect 17846 9382 17898 9434
rect 17898 9382 17900 9434
rect 17844 9380 17900 9382
rect 17948 9434 18004 9436
rect 17948 9382 17950 9434
rect 17950 9382 18002 9434
rect 18002 9382 18004 9434
rect 17948 9380 18004 9382
rect 18052 9434 18108 9436
rect 18052 9382 18054 9434
rect 18054 9382 18106 9434
rect 18106 9382 18108 9434
rect 18052 9380 18108 9382
rect 18620 9772 18676 9828
rect 18732 11228 18788 11284
rect 19068 11676 19124 11732
rect 22428 24610 22484 24612
rect 22428 24558 22430 24610
rect 22430 24558 22482 24610
rect 22482 24558 22484 24610
rect 22428 24556 22484 24558
rect 22002 24330 22058 24332
rect 22002 24278 22004 24330
rect 22004 24278 22056 24330
rect 22056 24278 22058 24330
rect 22002 24276 22058 24278
rect 22106 24330 22162 24332
rect 22106 24278 22108 24330
rect 22108 24278 22160 24330
rect 22160 24278 22162 24330
rect 22106 24276 22162 24278
rect 22210 24330 22266 24332
rect 22210 24278 22212 24330
rect 22212 24278 22264 24330
rect 22264 24278 22266 24330
rect 22210 24276 22266 24278
rect 23436 25676 23492 25732
rect 22988 24892 23044 24948
rect 23212 25228 23268 25284
rect 22764 23938 22820 23940
rect 22764 23886 22766 23938
rect 22766 23886 22818 23938
rect 22818 23886 22820 23938
rect 22764 23884 22820 23886
rect 20972 23212 21028 23268
rect 20636 22258 20692 22260
rect 20636 22206 20638 22258
rect 20638 22206 20690 22258
rect 20690 22206 20692 22258
rect 20636 22204 20692 22206
rect 20524 21698 20580 21700
rect 20524 21646 20526 21698
rect 20526 21646 20578 21698
rect 20578 21646 20580 21698
rect 20524 21644 20580 21646
rect 20412 20972 20468 21028
rect 22002 22762 22058 22764
rect 22002 22710 22004 22762
rect 22004 22710 22056 22762
rect 22056 22710 22058 22762
rect 22002 22708 22058 22710
rect 22106 22762 22162 22764
rect 22106 22710 22108 22762
rect 22108 22710 22160 22762
rect 22160 22710 22162 22762
rect 22106 22708 22162 22710
rect 22210 22762 22266 22764
rect 22210 22710 22212 22762
rect 22212 22710 22264 22762
rect 22264 22710 22266 22762
rect 22210 22708 22266 22710
rect 21420 22316 21476 22372
rect 20636 20018 20692 20020
rect 20636 19966 20638 20018
rect 20638 19966 20690 20018
rect 20690 19966 20692 20018
rect 20636 19964 20692 19966
rect 21196 20636 21252 20692
rect 22204 22258 22260 22260
rect 22204 22206 22206 22258
rect 22206 22206 22258 22258
rect 22258 22206 22260 22258
rect 22204 22204 22260 22206
rect 21980 21756 22036 21812
rect 21644 21698 21700 21700
rect 21644 21646 21646 21698
rect 21646 21646 21698 21698
rect 21698 21646 21700 21698
rect 21644 21644 21700 21646
rect 22652 21756 22708 21812
rect 21756 21420 21812 21476
rect 22002 21194 22058 21196
rect 22002 21142 22004 21194
rect 22004 21142 22056 21194
rect 22056 21142 22058 21194
rect 22002 21140 22058 21142
rect 22106 21194 22162 21196
rect 22106 21142 22108 21194
rect 22108 21142 22160 21194
rect 22160 21142 22162 21194
rect 22106 21140 22162 21142
rect 22210 21194 22266 21196
rect 22210 21142 22212 21194
rect 22212 21142 22264 21194
rect 22264 21142 22266 21194
rect 22210 21140 22266 21142
rect 22540 21026 22596 21028
rect 22540 20974 22542 21026
rect 22542 20974 22594 21026
rect 22594 20974 22596 21026
rect 22540 20972 22596 20974
rect 22988 23378 23044 23380
rect 22988 23326 22990 23378
rect 22990 23326 23042 23378
rect 23042 23326 23044 23378
rect 22988 23324 23044 23326
rect 21532 20748 21588 20804
rect 21084 20018 21140 20020
rect 21084 19966 21086 20018
rect 21086 19966 21138 20018
rect 21138 19966 21140 20018
rect 21084 19964 21140 19966
rect 20524 19292 20580 19348
rect 21308 17724 21364 17780
rect 20636 17388 20692 17444
rect 20076 16716 20132 16772
rect 21532 19906 21588 19908
rect 21532 19854 21534 19906
rect 21534 19854 21586 19906
rect 21586 19854 21588 19906
rect 21532 19852 21588 19854
rect 22876 20802 22932 20804
rect 22876 20750 22878 20802
rect 22878 20750 22930 20802
rect 22930 20750 22932 20802
rect 22876 20748 22932 20750
rect 22204 20076 22260 20132
rect 22988 20018 23044 20020
rect 22988 19966 22990 20018
rect 22990 19966 23042 20018
rect 23042 19966 23044 20018
rect 22988 19964 23044 19966
rect 21868 19906 21924 19908
rect 21868 19854 21870 19906
rect 21870 19854 21922 19906
rect 21922 19854 21924 19906
rect 21868 19852 21924 19854
rect 22002 19626 22058 19628
rect 22002 19574 22004 19626
rect 22004 19574 22056 19626
rect 22056 19574 22058 19626
rect 22002 19572 22058 19574
rect 22106 19626 22162 19628
rect 22106 19574 22108 19626
rect 22108 19574 22160 19626
rect 22160 19574 22162 19626
rect 22106 19572 22162 19574
rect 22210 19626 22266 19628
rect 22210 19574 22212 19626
rect 22212 19574 22264 19626
rect 22264 19574 22266 19626
rect 22210 19572 22266 19574
rect 21644 18620 21700 18676
rect 20972 15932 21028 15988
rect 22876 19068 22932 19124
rect 22876 18450 22932 18452
rect 22876 18398 22878 18450
rect 22878 18398 22930 18450
rect 22930 18398 22932 18450
rect 22876 18396 22932 18398
rect 24108 26124 24164 26180
rect 26160 26682 26216 26684
rect 26160 26630 26162 26682
rect 26162 26630 26214 26682
rect 26214 26630 26216 26682
rect 26160 26628 26216 26630
rect 26264 26682 26320 26684
rect 26264 26630 26266 26682
rect 26266 26630 26318 26682
rect 26318 26630 26320 26682
rect 26264 26628 26320 26630
rect 26368 26682 26424 26684
rect 26368 26630 26370 26682
rect 26370 26630 26422 26682
rect 26422 26630 26424 26682
rect 26368 26628 26424 26630
rect 34476 26682 34532 26684
rect 34476 26630 34478 26682
rect 34478 26630 34530 26682
rect 34530 26630 34532 26682
rect 34476 26628 34532 26630
rect 34580 26682 34636 26684
rect 34580 26630 34582 26682
rect 34582 26630 34634 26682
rect 34634 26630 34636 26682
rect 34580 26628 34636 26630
rect 34684 26682 34740 26684
rect 34684 26630 34686 26682
rect 34686 26630 34738 26682
rect 34738 26630 34740 26682
rect 34684 26628 34740 26630
rect 25340 25340 25396 25396
rect 25228 25228 25284 25284
rect 24332 24946 24388 24948
rect 24332 24894 24334 24946
rect 24334 24894 24386 24946
rect 24386 24894 24388 24946
rect 24332 24892 24388 24894
rect 23772 23884 23828 23940
rect 23436 23772 23492 23828
rect 24668 24668 24724 24724
rect 25564 24668 25620 24724
rect 25788 25340 25844 25396
rect 25564 23938 25620 23940
rect 25564 23886 25566 23938
rect 25566 23886 25618 23938
rect 25618 23886 25620 23938
rect 25564 23884 25620 23886
rect 24332 23772 24388 23828
rect 24780 23714 24836 23716
rect 24780 23662 24782 23714
rect 24782 23662 24834 23714
rect 24834 23662 24836 23714
rect 24780 23660 24836 23662
rect 25228 23660 25284 23716
rect 23884 23378 23940 23380
rect 23884 23326 23886 23378
rect 23886 23326 23938 23378
rect 23938 23326 23940 23378
rect 23884 23324 23940 23326
rect 24668 23378 24724 23380
rect 24668 23326 24670 23378
rect 24670 23326 24722 23378
rect 24722 23326 24724 23378
rect 24668 23324 24724 23326
rect 24444 23154 24500 23156
rect 24444 23102 24446 23154
rect 24446 23102 24498 23154
rect 24498 23102 24500 23154
rect 24444 23100 24500 23102
rect 30318 25898 30374 25900
rect 30318 25846 30320 25898
rect 30320 25846 30372 25898
rect 30372 25846 30374 25898
rect 30318 25844 30374 25846
rect 30422 25898 30478 25900
rect 30422 25846 30424 25898
rect 30424 25846 30476 25898
rect 30476 25846 30478 25898
rect 30422 25844 30478 25846
rect 30526 25898 30582 25900
rect 30526 25846 30528 25898
rect 30528 25846 30580 25898
rect 30580 25846 30582 25898
rect 30526 25844 30582 25846
rect 26160 25114 26216 25116
rect 26160 25062 26162 25114
rect 26162 25062 26214 25114
rect 26214 25062 26216 25114
rect 26160 25060 26216 25062
rect 26264 25114 26320 25116
rect 26264 25062 26266 25114
rect 26266 25062 26318 25114
rect 26318 25062 26320 25114
rect 26264 25060 26320 25062
rect 26368 25114 26424 25116
rect 26368 25062 26370 25114
rect 26370 25062 26422 25114
rect 26422 25062 26424 25114
rect 26368 25060 26424 25062
rect 26908 25394 26964 25396
rect 26908 25342 26910 25394
rect 26910 25342 26962 25394
rect 26962 25342 26964 25394
rect 26908 25340 26964 25342
rect 27356 25394 27412 25396
rect 27356 25342 27358 25394
rect 27358 25342 27410 25394
rect 27410 25342 27412 25394
rect 27356 25340 27412 25342
rect 26684 25282 26740 25284
rect 26684 25230 26686 25282
rect 26686 25230 26738 25282
rect 26738 25230 26740 25282
rect 26684 25228 26740 25230
rect 27468 24892 27524 24948
rect 25900 24780 25956 24836
rect 26012 24668 26068 24724
rect 25676 23324 25732 23380
rect 25452 23212 25508 23268
rect 25788 23996 25844 24052
rect 25788 22428 25844 22484
rect 25676 22146 25732 22148
rect 25676 22094 25678 22146
rect 25678 22094 25730 22146
rect 25730 22094 25732 22146
rect 25676 22092 25732 22094
rect 24444 21810 24500 21812
rect 24444 21758 24446 21810
rect 24446 21758 24498 21810
rect 24498 21758 24500 21810
rect 24444 21756 24500 21758
rect 25452 21810 25508 21812
rect 25452 21758 25454 21810
rect 25454 21758 25506 21810
rect 25506 21758 25508 21810
rect 25452 21756 25508 21758
rect 23548 21644 23604 21700
rect 23884 21586 23940 21588
rect 23884 21534 23886 21586
rect 23886 21534 23938 21586
rect 23938 21534 23940 21586
rect 23884 21532 23940 21534
rect 24444 20860 24500 20916
rect 24556 21420 24612 21476
rect 22540 18284 22596 18340
rect 22002 18058 22058 18060
rect 22002 18006 22004 18058
rect 22004 18006 22056 18058
rect 22056 18006 22058 18058
rect 22002 18004 22058 18006
rect 22106 18058 22162 18060
rect 22106 18006 22108 18058
rect 22108 18006 22160 18058
rect 22160 18006 22162 18058
rect 22106 18004 22162 18006
rect 22210 18058 22266 18060
rect 22210 18006 22212 18058
rect 22212 18006 22264 18058
rect 22264 18006 22266 18058
rect 22210 18004 22266 18006
rect 21756 17724 21812 17780
rect 23212 18172 23268 18228
rect 23436 20076 23492 20132
rect 21644 16156 21700 16212
rect 22540 16716 22596 16772
rect 21756 16044 21812 16100
rect 21868 16604 21924 16660
rect 22876 16604 22932 16660
rect 22002 16490 22058 16492
rect 22002 16438 22004 16490
rect 22004 16438 22056 16490
rect 22056 16438 22058 16490
rect 22002 16436 22058 16438
rect 22106 16490 22162 16492
rect 22106 16438 22108 16490
rect 22108 16438 22160 16490
rect 22160 16438 22162 16490
rect 22106 16436 22162 16438
rect 22210 16490 22266 16492
rect 22210 16438 22212 16490
rect 22212 16438 22264 16490
rect 22264 16438 22266 16490
rect 22210 16436 22266 16438
rect 22428 16098 22484 16100
rect 22428 16046 22430 16098
rect 22430 16046 22482 16098
rect 22482 16046 22484 16098
rect 22428 16044 22484 16046
rect 21532 15986 21588 15988
rect 21532 15934 21534 15986
rect 21534 15934 21586 15986
rect 21586 15934 21588 15986
rect 21532 15932 21588 15934
rect 19964 14364 20020 14420
rect 19516 13916 19572 13972
rect 19628 13804 19684 13860
rect 19852 14028 19908 14084
rect 20076 13916 20132 13972
rect 19740 13692 19796 13748
rect 19516 13468 19572 13524
rect 19740 12738 19796 12740
rect 19740 12686 19742 12738
rect 19742 12686 19794 12738
rect 19794 12686 19796 12738
rect 19740 12684 19796 12686
rect 19404 12236 19460 12292
rect 20300 13804 20356 13860
rect 20188 13746 20244 13748
rect 20188 13694 20190 13746
rect 20190 13694 20242 13746
rect 20242 13694 20244 13746
rect 20188 13692 20244 13694
rect 20300 13186 20356 13188
rect 20300 13134 20302 13186
rect 20302 13134 20354 13186
rect 20354 13134 20356 13186
rect 20300 13132 20356 13134
rect 20076 13074 20132 13076
rect 20076 13022 20078 13074
rect 20078 13022 20130 13074
rect 20130 13022 20132 13074
rect 20076 13020 20132 13022
rect 20524 14306 20580 14308
rect 20524 14254 20526 14306
rect 20526 14254 20578 14306
rect 20578 14254 20580 14306
rect 20524 14252 20580 14254
rect 20748 13020 20804 13076
rect 20524 12962 20580 12964
rect 20524 12910 20526 12962
rect 20526 12910 20578 12962
rect 20578 12910 20580 12962
rect 20524 12908 20580 12910
rect 22652 15986 22708 15988
rect 22652 15934 22654 15986
rect 22654 15934 22706 15986
rect 22706 15934 22708 15986
rect 22652 15932 22708 15934
rect 21196 14028 21252 14084
rect 19180 11452 19236 11508
rect 19628 11676 19684 11732
rect 19852 11564 19908 11620
rect 19964 12348 20020 12404
rect 20748 12572 20804 12628
rect 20636 12402 20692 12404
rect 20636 12350 20638 12402
rect 20638 12350 20690 12402
rect 20690 12350 20692 12402
rect 20636 12348 20692 12350
rect 20972 12684 21028 12740
rect 21644 14588 21700 14644
rect 21420 14252 21476 14308
rect 21308 13522 21364 13524
rect 21308 13470 21310 13522
rect 21310 13470 21362 13522
rect 21362 13470 21364 13522
rect 21308 13468 21364 13470
rect 21644 13468 21700 13524
rect 21756 13020 21812 13076
rect 22002 14922 22058 14924
rect 22002 14870 22004 14922
rect 22004 14870 22056 14922
rect 22056 14870 22058 14922
rect 22002 14868 22058 14870
rect 22106 14922 22162 14924
rect 22106 14870 22108 14922
rect 22108 14870 22160 14922
rect 22160 14870 22162 14922
rect 22106 14868 22162 14870
rect 22210 14922 22266 14924
rect 22210 14870 22212 14922
rect 22212 14870 22264 14922
rect 22264 14870 22266 14922
rect 22210 14868 22266 14870
rect 22204 13916 22260 13972
rect 21980 13522 22036 13524
rect 21980 13470 21982 13522
rect 21982 13470 22034 13522
rect 22034 13470 22036 13522
rect 21980 13468 22036 13470
rect 22002 13354 22058 13356
rect 22002 13302 22004 13354
rect 22004 13302 22056 13354
rect 22056 13302 22058 13354
rect 22002 13300 22058 13302
rect 22106 13354 22162 13356
rect 22106 13302 22108 13354
rect 22108 13302 22160 13354
rect 22160 13302 22162 13354
rect 22106 13300 22162 13302
rect 22210 13354 22266 13356
rect 22210 13302 22212 13354
rect 22212 13302 22264 13354
rect 22264 13302 22266 13354
rect 22210 13300 22266 13302
rect 22092 13186 22148 13188
rect 22092 13134 22094 13186
rect 22094 13134 22146 13186
rect 22146 13134 22148 13186
rect 22092 13132 22148 13134
rect 22652 13132 22708 13188
rect 22428 13020 22484 13076
rect 21868 12962 21924 12964
rect 21868 12910 21870 12962
rect 21870 12910 21922 12962
rect 21922 12910 21924 12962
rect 21868 12908 21924 12910
rect 22316 12962 22372 12964
rect 22316 12910 22318 12962
rect 22318 12910 22370 12962
rect 22370 12910 22372 12962
rect 22316 12908 22372 12910
rect 21644 12850 21700 12852
rect 21644 12798 21646 12850
rect 21646 12798 21698 12850
rect 21698 12798 21700 12850
rect 21644 12796 21700 12798
rect 20076 11676 20132 11732
rect 20412 11618 20468 11620
rect 20412 11566 20414 11618
rect 20414 11566 20466 11618
rect 20466 11566 20468 11618
rect 20412 11564 20468 11566
rect 21308 11676 21364 11732
rect 17724 8988 17780 9044
rect 17948 8876 18004 8932
rect 16716 7868 16772 7924
rect 16156 5906 16212 5908
rect 16156 5854 16158 5906
rect 16158 5854 16210 5906
rect 16210 5854 16212 5906
rect 16156 5852 16212 5854
rect 16828 7474 16884 7476
rect 16828 7422 16830 7474
rect 16830 7422 16882 7474
rect 16882 7422 16884 7474
rect 16828 7420 16884 7422
rect 17844 7866 17900 7868
rect 17844 7814 17846 7866
rect 17846 7814 17898 7866
rect 17898 7814 17900 7866
rect 17844 7812 17900 7814
rect 17948 7866 18004 7868
rect 17948 7814 17950 7866
rect 17950 7814 18002 7866
rect 18002 7814 18004 7866
rect 17948 7812 18004 7814
rect 18052 7866 18108 7868
rect 18052 7814 18054 7866
rect 18054 7814 18106 7866
rect 18106 7814 18108 7866
rect 18052 7812 18108 7814
rect 17164 6636 17220 6692
rect 17388 6018 17444 6020
rect 17388 5966 17390 6018
rect 17390 5966 17442 6018
rect 17442 5966 17444 6018
rect 17388 5964 17444 5966
rect 15372 3612 15428 3668
rect 16268 5628 16324 5684
rect 16268 4508 16324 4564
rect 18732 7420 18788 7476
rect 18844 10108 18900 10164
rect 19740 9996 19796 10052
rect 20972 10108 21028 10164
rect 19180 9884 19236 9940
rect 20076 9826 20132 9828
rect 20076 9774 20078 9826
rect 20078 9774 20130 9826
rect 20130 9774 20132 9826
rect 20076 9772 20132 9774
rect 20636 9826 20692 9828
rect 20636 9774 20638 9826
rect 20638 9774 20690 9826
rect 20690 9774 20692 9826
rect 20636 9772 20692 9774
rect 18956 9714 19012 9716
rect 18956 9662 18958 9714
rect 18958 9662 19010 9714
rect 19010 9662 19012 9714
rect 18956 9660 19012 9662
rect 22316 12572 22372 12628
rect 24444 20130 24500 20132
rect 24444 20078 24446 20130
rect 24446 20078 24498 20130
rect 24498 20078 24500 20130
rect 24444 20076 24500 20078
rect 25452 21362 25508 21364
rect 25452 21310 25454 21362
rect 25454 21310 25506 21362
rect 25506 21310 25508 21362
rect 25452 21308 25508 21310
rect 24668 20018 24724 20020
rect 24668 19966 24670 20018
rect 24670 19966 24722 20018
rect 24722 19966 24724 20018
rect 24668 19964 24724 19966
rect 25228 20018 25284 20020
rect 25228 19966 25230 20018
rect 25230 19966 25282 20018
rect 25282 19966 25284 20018
rect 25228 19964 25284 19966
rect 26460 23996 26516 24052
rect 26124 23772 26180 23828
rect 26160 23546 26216 23548
rect 26160 23494 26162 23546
rect 26162 23494 26214 23546
rect 26214 23494 26216 23546
rect 26160 23492 26216 23494
rect 26264 23546 26320 23548
rect 26264 23494 26266 23546
rect 26266 23494 26318 23546
rect 26318 23494 26320 23546
rect 26264 23492 26320 23494
rect 26368 23546 26424 23548
rect 26368 23494 26370 23546
rect 26370 23494 26422 23546
rect 26422 23494 26424 23546
rect 26368 23492 26424 23494
rect 26124 23100 26180 23156
rect 26124 22594 26180 22596
rect 26124 22542 26126 22594
rect 26126 22542 26178 22594
rect 26178 22542 26180 22594
rect 26124 22540 26180 22542
rect 26684 23884 26740 23940
rect 27916 23996 27972 24052
rect 28140 23938 28196 23940
rect 28140 23886 28142 23938
rect 28142 23886 28194 23938
rect 28194 23886 28196 23938
rect 28140 23884 28196 23886
rect 27132 23826 27188 23828
rect 27132 23774 27134 23826
rect 27134 23774 27186 23826
rect 27186 23774 27188 23826
rect 27132 23772 27188 23774
rect 26796 23660 26852 23716
rect 27244 23714 27300 23716
rect 27244 23662 27246 23714
rect 27246 23662 27298 23714
rect 27298 23662 27300 23714
rect 27244 23660 27300 23662
rect 27468 23714 27524 23716
rect 27468 23662 27470 23714
rect 27470 23662 27522 23714
rect 27522 23662 27524 23714
rect 27468 23660 27524 23662
rect 34476 25114 34532 25116
rect 34476 25062 34478 25114
rect 34478 25062 34530 25114
rect 34530 25062 34532 25114
rect 34476 25060 34532 25062
rect 34580 25114 34636 25116
rect 34580 25062 34582 25114
rect 34582 25062 34634 25114
rect 34634 25062 34636 25114
rect 34580 25060 34636 25062
rect 34684 25114 34740 25116
rect 34684 25062 34686 25114
rect 34686 25062 34738 25114
rect 34738 25062 34740 25114
rect 34684 25060 34740 25062
rect 28700 24892 28756 24948
rect 29372 24780 29428 24836
rect 30044 24780 30100 24836
rect 29372 23996 29428 24052
rect 29148 23826 29204 23828
rect 29148 23774 29150 23826
rect 29150 23774 29202 23826
rect 29202 23774 29204 23826
rect 29148 23772 29204 23774
rect 28364 23714 28420 23716
rect 28364 23662 28366 23714
rect 28366 23662 28418 23714
rect 28418 23662 28420 23714
rect 28364 23660 28420 23662
rect 27020 23212 27076 23268
rect 29932 23714 29988 23716
rect 29932 23662 29934 23714
rect 29934 23662 29986 23714
rect 29986 23662 29988 23714
rect 29932 23660 29988 23662
rect 30318 24330 30374 24332
rect 30318 24278 30320 24330
rect 30320 24278 30372 24330
rect 30372 24278 30374 24330
rect 30318 24276 30374 24278
rect 30422 24330 30478 24332
rect 30422 24278 30424 24330
rect 30424 24278 30476 24330
rect 30476 24278 30478 24330
rect 30422 24276 30478 24278
rect 30526 24330 30582 24332
rect 30526 24278 30528 24330
rect 30528 24278 30580 24330
rect 30580 24278 30582 24330
rect 30526 24276 30582 24278
rect 34476 23546 34532 23548
rect 34476 23494 34478 23546
rect 34478 23494 34530 23546
rect 34530 23494 34532 23546
rect 34476 23492 34532 23494
rect 34580 23546 34636 23548
rect 34580 23494 34582 23546
rect 34582 23494 34634 23546
rect 34634 23494 34636 23546
rect 34580 23492 34636 23494
rect 34684 23546 34740 23548
rect 34684 23494 34686 23546
rect 34686 23494 34738 23546
rect 34738 23494 34740 23546
rect 34684 23492 34740 23494
rect 26908 22540 26964 22596
rect 26124 22092 26180 22148
rect 26160 21978 26216 21980
rect 26160 21926 26162 21978
rect 26162 21926 26214 21978
rect 26214 21926 26216 21978
rect 26160 21924 26216 21926
rect 26264 21978 26320 21980
rect 26264 21926 26266 21978
rect 26266 21926 26318 21978
rect 26318 21926 26320 21978
rect 26264 21924 26320 21926
rect 26368 21978 26424 21980
rect 26368 21926 26370 21978
rect 26370 21926 26422 21978
rect 26422 21926 26424 21978
rect 26368 21924 26424 21926
rect 26684 21756 26740 21812
rect 26124 21532 26180 21588
rect 25900 21196 25956 21252
rect 26012 20914 26068 20916
rect 26012 20862 26014 20914
rect 26014 20862 26066 20914
rect 26066 20862 26068 20914
rect 26012 20860 26068 20862
rect 26160 20410 26216 20412
rect 26160 20358 26162 20410
rect 26162 20358 26214 20410
rect 26214 20358 26216 20410
rect 26160 20356 26216 20358
rect 26264 20410 26320 20412
rect 26264 20358 26266 20410
rect 26266 20358 26318 20410
rect 26318 20358 26320 20410
rect 26264 20356 26320 20358
rect 26368 20410 26424 20412
rect 26368 20358 26370 20410
rect 26370 20358 26422 20410
rect 26422 20358 26424 20410
rect 26368 20356 26424 20358
rect 27132 22482 27188 22484
rect 27132 22430 27134 22482
rect 27134 22430 27186 22482
rect 27186 22430 27188 22482
rect 27132 22428 27188 22430
rect 27244 22146 27300 22148
rect 27244 22094 27246 22146
rect 27246 22094 27298 22146
rect 27298 22094 27300 22146
rect 27244 22092 27300 22094
rect 27020 21756 27076 21812
rect 27244 21532 27300 21588
rect 27020 21308 27076 21364
rect 30318 22762 30374 22764
rect 30318 22710 30320 22762
rect 30320 22710 30372 22762
rect 30372 22710 30374 22762
rect 30318 22708 30374 22710
rect 30422 22762 30478 22764
rect 30422 22710 30424 22762
rect 30424 22710 30476 22762
rect 30476 22710 30478 22762
rect 30422 22708 30478 22710
rect 30526 22762 30582 22764
rect 30526 22710 30528 22762
rect 30528 22710 30580 22762
rect 30580 22710 30582 22762
rect 30526 22708 30582 22710
rect 34476 21978 34532 21980
rect 34476 21926 34478 21978
rect 34478 21926 34530 21978
rect 34530 21926 34532 21978
rect 34476 21924 34532 21926
rect 34580 21978 34636 21980
rect 34580 21926 34582 21978
rect 34582 21926 34634 21978
rect 34634 21926 34636 21978
rect 34580 21924 34636 21926
rect 34684 21978 34740 21980
rect 34684 21926 34686 21978
rect 34686 21926 34738 21978
rect 34738 21926 34740 21978
rect 34684 21924 34740 21926
rect 27468 21420 27524 21476
rect 28812 21474 28868 21476
rect 28812 21422 28814 21474
rect 28814 21422 28866 21474
rect 28866 21422 28868 21474
rect 28812 21420 28868 21422
rect 27580 21196 27636 21252
rect 30318 21194 30374 21196
rect 30318 21142 30320 21194
rect 30320 21142 30372 21194
rect 30372 21142 30374 21194
rect 30318 21140 30374 21142
rect 30422 21194 30478 21196
rect 30422 21142 30424 21194
rect 30424 21142 30476 21194
rect 30476 21142 30478 21194
rect 30422 21140 30478 21142
rect 30526 21194 30582 21196
rect 30526 21142 30528 21194
rect 30528 21142 30580 21194
rect 30580 21142 30582 21194
rect 30526 21140 30582 21142
rect 34476 20410 34532 20412
rect 34476 20358 34478 20410
rect 34478 20358 34530 20410
rect 34530 20358 34532 20410
rect 34476 20356 34532 20358
rect 34580 20410 34636 20412
rect 34580 20358 34582 20410
rect 34582 20358 34634 20410
rect 34634 20358 34636 20410
rect 34580 20356 34636 20358
rect 34684 20410 34740 20412
rect 34684 20358 34686 20410
rect 34686 20358 34738 20410
rect 34738 20358 34740 20410
rect 34684 20356 34740 20358
rect 29708 20076 29764 20132
rect 30604 20076 30660 20132
rect 27132 20018 27188 20020
rect 27132 19966 27134 20018
rect 27134 19966 27186 20018
rect 27186 19966 27188 20018
rect 27132 19964 27188 19966
rect 29148 19964 29204 20020
rect 26684 19740 26740 19796
rect 26460 19346 26516 19348
rect 26460 19294 26462 19346
rect 26462 19294 26514 19346
rect 26514 19294 26516 19346
rect 26460 19292 26516 19294
rect 27132 19292 27188 19348
rect 26160 18842 26216 18844
rect 26160 18790 26162 18842
rect 26162 18790 26214 18842
rect 26214 18790 26216 18842
rect 26160 18788 26216 18790
rect 26264 18842 26320 18844
rect 26264 18790 26266 18842
rect 26266 18790 26318 18842
rect 26318 18790 26320 18842
rect 26264 18788 26320 18790
rect 26368 18842 26424 18844
rect 26368 18790 26370 18842
rect 26370 18790 26422 18842
rect 26422 18790 26424 18842
rect 26368 18788 26424 18790
rect 23548 18450 23604 18452
rect 23548 18398 23550 18450
rect 23550 18398 23602 18450
rect 23602 18398 23604 18450
rect 23548 18396 23604 18398
rect 23548 17778 23604 17780
rect 23548 17726 23550 17778
rect 23550 17726 23602 17778
rect 23602 17726 23604 17778
rect 23548 17724 23604 17726
rect 25676 18396 25732 18452
rect 25452 18338 25508 18340
rect 25452 18286 25454 18338
rect 25454 18286 25506 18338
rect 25506 18286 25508 18338
rect 25452 18284 25508 18286
rect 23436 16604 23492 16660
rect 24556 17724 24612 17780
rect 23436 16210 23492 16212
rect 23436 16158 23438 16210
rect 23438 16158 23490 16210
rect 23490 16158 23492 16210
rect 23436 16156 23492 16158
rect 23436 14642 23492 14644
rect 23436 14590 23438 14642
rect 23438 14590 23490 14642
rect 23490 14590 23492 14642
rect 23436 14588 23492 14590
rect 24556 16604 24612 16660
rect 23660 16098 23716 16100
rect 23660 16046 23662 16098
rect 23662 16046 23714 16098
rect 23714 16046 23716 16098
rect 23660 16044 23716 16046
rect 24332 15986 24388 15988
rect 24332 15934 24334 15986
rect 24334 15934 24386 15986
rect 24386 15934 24388 15986
rect 24332 15932 24388 15934
rect 23996 15260 24052 15316
rect 26160 17274 26216 17276
rect 26160 17222 26162 17274
rect 26162 17222 26214 17274
rect 26214 17222 26216 17274
rect 26160 17220 26216 17222
rect 26264 17274 26320 17276
rect 26264 17222 26266 17274
rect 26266 17222 26318 17274
rect 26318 17222 26320 17274
rect 26264 17220 26320 17222
rect 26368 17274 26424 17276
rect 26368 17222 26370 17274
rect 26370 17222 26422 17274
rect 26422 17222 26424 17274
rect 26368 17220 26424 17222
rect 25788 16268 25844 16324
rect 26124 16716 26180 16772
rect 26236 16098 26292 16100
rect 26236 16046 26238 16098
rect 26238 16046 26290 16098
rect 26290 16046 26292 16098
rect 26236 16044 26292 16046
rect 26124 15986 26180 15988
rect 26124 15934 26126 15986
rect 26126 15934 26178 15986
rect 26178 15934 26180 15986
rect 26124 15932 26180 15934
rect 26012 15874 26068 15876
rect 26012 15822 26014 15874
rect 26014 15822 26066 15874
rect 26066 15822 26068 15874
rect 26012 15820 26068 15822
rect 26160 15706 26216 15708
rect 26160 15654 26162 15706
rect 26162 15654 26214 15706
rect 26214 15654 26216 15706
rect 26160 15652 26216 15654
rect 26264 15706 26320 15708
rect 26264 15654 26266 15706
rect 26266 15654 26318 15706
rect 26318 15654 26320 15706
rect 26264 15652 26320 15654
rect 26368 15706 26424 15708
rect 26368 15654 26370 15706
rect 26370 15654 26422 15706
rect 26422 15654 26424 15706
rect 26368 15652 26424 15654
rect 25452 14364 25508 14420
rect 22764 13020 22820 13076
rect 22988 13468 23044 13524
rect 22428 12012 22484 12068
rect 22002 11786 22058 11788
rect 22002 11734 22004 11786
rect 22004 11734 22056 11786
rect 22056 11734 22058 11786
rect 22002 11732 22058 11734
rect 22106 11786 22162 11788
rect 22106 11734 22108 11786
rect 22108 11734 22160 11786
rect 22160 11734 22162 11786
rect 22106 11732 22162 11734
rect 22210 11786 22266 11788
rect 22210 11734 22212 11786
rect 22212 11734 22264 11786
rect 22264 11734 22266 11786
rect 22210 11732 22266 11734
rect 22540 11452 22596 11508
rect 22876 12850 22932 12852
rect 22876 12798 22878 12850
rect 22878 12798 22930 12850
rect 22930 12798 22932 12850
rect 22876 12796 22932 12798
rect 22540 10834 22596 10836
rect 22540 10782 22542 10834
rect 22542 10782 22594 10834
rect 22594 10782 22596 10834
rect 22540 10780 22596 10782
rect 22092 10722 22148 10724
rect 22092 10670 22094 10722
rect 22094 10670 22146 10722
rect 22146 10670 22148 10722
rect 22092 10668 22148 10670
rect 21420 10108 21476 10164
rect 21308 10050 21364 10052
rect 21308 9998 21310 10050
rect 21310 9998 21362 10050
rect 21362 9998 21364 10050
rect 21308 9996 21364 9998
rect 21420 9938 21476 9940
rect 21420 9886 21422 9938
rect 21422 9886 21474 9938
rect 21474 9886 21476 9938
rect 21420 9884 21476 9886
rect 18956 8876 19012 8932
rect 19068 8764 19124 8820
rect 23884 13746 23940 13748
rect 23884 13694 23886 13746
rect 23886 13694 23938 13746
rect 23938 13694 23940 13746
rect 23884 13692 23940 13694
rect 26684 18172 26740 18228
rect 28028 18956 28084 19012
rect 27468 17724 27524 17780
rect 29036 17724 29092 17780
rect 28028 16940 28084 16996
rect 27580 16828 27636 16884
rect 27468 16322 27524 16324
rect 27468 16270 27470 16322
rect 27470 16270 27522 16322
rect 27522 16270 27524 16322
rect 27468 16268 27524 16270
rect 27916 15986 27972 15988
rect 27916 15934 27918 15986
rect 27918 15934 27970 15986
rect 27970 15934 27972 15986
rect 27916 15932 27972 15934
rect 27468 15874 27524 15876
rect 27468 15822 27470 15874
rect 27470 15822 27522 15874
rect 27522 15822 27524 15874
rect 27468 15820 27524 15822
rect 28924 17612 28980 17668
rect 28140 16770 28196 16772
rect 28140 16718 28142 16770
rect 28142 16718 28194 16770
rect 28194 16718 28196 16770
rect 28140 16716 28196 16718
rect 28252 15932 28308 15988
rect 28028 15820 28084 15876
rect 28140 15372 28196 15428
rect 28028 15260 28084 15316
rect 27356 15148 27412 15204
rect 27244 14530 27300 14532
rect 27244 14478 27246 14530
rect 27246 14478 27298 14530
rect 27298 14478 27300 14530
rect 27244 14476 27300 14478
rect 25676 13858 25732 13860
rect 25676 13806 25678 13858
rect 25678 13806 25730 13858
rect 25730 13806 25732 13858
rect 25676 13804 25732 13806
rect 25452 13746 25508 13748
rect 25452 13694 25454 13746
rect 25454 13694 25506 13746
rect 25506 13694 25508 13746
rect 25452 13692 25508 13694
rect 24780 13468 24836 13524
rect 24220 12066 24276 12068
rect 24220 12014 24222 12066
rect 24222 12014 24274 12066
rect 24274 12014 24276 12066
rect 24220 12012 24276 12014
rect 22002 10218 22058 10220
rect 22002 10166 22004 10218
rect 22004 10166 22056 10218
rect 22056 10166 22058 10218
rect 22002 10164 22058 10166
rect 22106 10218 22162 10220
rect 22106 10166 22108 10218
rect 22108 10166 22160 10218
rect 22160 10166 22162 10218
rect 22106 10164 22162 10166
rect 22210 10218 22266 10220
rect 22210 10166 22212 10218
rect 22212 10166 22264 10218
rect 22264 10166 22266 10218
rect 22210 10164 22266 10166
rect 23100 9996 23156 10052
rect 22092 9826 22148 9828
rect 22092 9774 22094 9826
rect 22094 9774 22146 9826
rect 22146 9774 22148 9826
rect 22092 9772 22148 9774
rect 21868 9212 21924 9268
rect 23100 9660 23156 9716
rect 22002 8650 22058 8652
rect 22002 8598 22004 8650
rect 22004 8598 22056 8650
rect 22056 8598 22058 8650
rect 22002 8596 22058 8598
rect 22106 8650 22162 8652
rect 22106 8598 22108 8650
rect 22108 8598 22160 8650
rect 22160 8598 22162 8650
rect 22106 8596 22162 8598
rect 22210 8650 22266 8652
rect 22210 8598 22212 8650
rect 22212 8598 22264 8650
rect 22264 8598 22266 8650
rect 22210 8596 22266 8598
rect 17844 6298 17900 6300
rect 17844 6246 17846 6298
rect 17846 6246 17898 6298
rect 17898 6246 17900 6298
rect 17844 6244 17900 6246
rect 17948 6298 18004 6300
rect 17948 6246 17950 6298
rect 17950 6246 18002 6298
rect 18002 6246 18004 6298
rect 17948 6244 18004 6246
rect 18052 6298 18108 6300
rect 18052 6246 18054 6298
rect 18054 6246 18106 6298
rect 18106 6246 18108 6298
rect 18052 6244 18108 6246
rect 17948 6130 18004 6132
rect 17948 6078 17950 6130
rect 17950 6078 18002 6130
rect 18002 6078 18004 6130
rect 17948 6076 18004 6078
rect 17500 5740 17556 5796
rect 16940 5068 16996 5124
rect 16828 4284 16884 4340
rect 18284 5180 18340 5236
rect 18172 5122 18228 5124
rect 18172 5070 18174 5122
rect 18174 5070 18226 5122
rect 18226 5070 18228 5122
rect 18172 5068 18228 5070
rect 17724 5010 17780 5012
rect 17724 4958 17726 5010
rect 17726 4958 17778 5010
rect 17778 4958 17780 5010
rect 17724 4956 17780 4958
rect 17276 4562 17332 4564
rect 17276 4510 17278 4562
rect 17278 4510 17330 4562
rect 17330 4510 17332 4562
rect 17276 4508 17332 4510
rect 17612 4338 17668 4340
rect 17612 4286 17614 4338
rect 17614 4286 17666 4338
rect 17666 4286 17668 4338
rect 17612 4284 17668 4286
rect 17844 4730 17900 4732
rect 17844 4678 17846 4730
rect 17846 4678 17898 4730
rect 17898 4678 17900 4730
rect 17844 4676 17900 4678
rect 17948 4730 18004 4732
rect 17948 4678 17950 4730
rect 17950 4678 18002 4730
rect 18002 4678 18004 4730
rect 17948 4676 18004 4678
rect 18052 4730 18108 4732
rect 18052 4678 18054 4730
rect 18054 4678 18106 4730
rect 18106 4678 18108 4730
rect 18052 4676 18108 4678
rect 18060 4508 18116 4564
rect 12572 3500 12628 3556
rect 14364 3554 14420 3556
rect 14364 3502 14366 3554
rect 14366 3502 14418 3554
rect 14418 3502 14420 3554
rect 14364 3500 14420 3502
rect 15484 3500 15540 3556
rect 13244 3442 13300 3444
rect 13244 3390 13246 3442
rect 13246 3390 13298 3442
rect 13298 3390 13300 3442
rect 13244 3388 13300 3390
rect 11900 3276 11956 3332
rect 17844 3162 17900 3164
rect 11788 3052 11844 3108
rect 17844 3110 17846 3162
rect 17846 3110 17898 3162
rect 17898 3110 17900 3162
rect 17844 3108 17900 3110
rect 17948 3162 18004 3164
rect 17948 3110 17950 3162
rect 17950 3110 18002 3162
rect 18002 3110 18004 3162
rect 17948 3108 18004 3110
rect 18052 3162 18108 3164
rect 18052 3110 18054 3162
rect 18054 3110 18106 3162
rect 18106 3110 18108 3162
rect 18052 3108 18108 3110
rect 18732 5068 18788 5124
rect 18620 4956 18676 5012
rect 19180 7420 19236 7476
rect 18956 6076 19012 6132
rect 19180 6802 19236 6804
rect 19180 6750 19182 6802
rect 19182 6750 19234 6802
rect 19234 6750 19236 6802
rect 19180 6748 19236 6750
rect 18844 4956 18900 5012
rect 19740 6748 19796 6804
rect 19516 6076 19572 6132
rect 21308 6076 21364 6132
rect 20076 5964 20132 6020
rect 19292 5906 19348 5908
rect 19292 5854 19294 5906
rect 19294 5854 19346 5906
rect 19346 5854 19348 5906
rect 19292 5852 19348 5854
rect 20524 6018 20580 6020
rect 20524 5966 20526 6018
rect 20526 5966 20578 6018
rect 20578 5966 20580 6018
rect 20524 5964 20580 5966
rect 20972 6018 21028 6020
rect 20972 5966 20974 6018
rect 20974 5966 21026 6018
rect 21026 5966 21028 6018
rect 20972 5964 21028 5966
rect 21756 8034 21812 8036
rect 21756 7982 21758 8034
rect 21758 7982 21810 8034
rect 21810 7982 21812 8034
rect 21756 7980 21812 7982
rect 21644 7420 21700 7476
rect 21420 5964 21476 6020
rect 21532 7196 21588 7252
rect 22204 7474 22260 7476
rect 22204 7422 22206 7474
rect 22206 7422 22258 7474
rect 22258 7422 22260 7474
rect 22204 7420 22260 7422
rect 22002 7082 22058 7084
rect 22002 7030 22004 7082
rect 22004 7030 22056 7082
rect 22056 7030 22058 7082
rect 22002 7028 22058 7030
rect 22106 7082 22162 7084
rect 22106 7030 22108 7082
rect 22108 7030 22160 7082
rect 22160 7030 22162 7082
rect 22106 7028 22162 7030
rect 22210 7082 22266 7084
rect 22210 7030 22212 7082
rect 22212 7030 22264 7082
rect 22264 7030 22266 7082
rect 22210 7028 22266 7030
rect 22092 6860 22148 6916
rect 21868 6748 21924 6804
rect 21532 5852 21588 5908
rect 21644 5964 21700 6020
rect 19180 5234 19236 5236
rect 19180 5182 19182 5234
rect 19182 5182 19234 5234
rect 19234 5182 19236 5234
rect 19180 5180 19236 5182
rect 19068 4562 19124 4564
rect 19068 4510 19070 4562
rect 19070 4510 19122 4562
rect 19122 4510 19124 4562
rect 19068 4508 19124 4510
rect 19516 4956 19572 5012
rect 19740 3554 19796 3556
rect 19740 3502 19742 3554
rect 19742 3502 19794 3554
rect 19794 3502 19796 3554
rect 19740 3500 19796 3502
rect 21644 5234 21700 5236
rect 21644 5182 21646 5234
rect 21646 5182 21698 5234
rect 21698 5182 21700 5234
rect 21644 5180 21700 5182
rect 20300 4226 20356 4228
rect 20300 4174 20302 4226
rect 20302 4174 20354 4226
rect 20354 4174 20356 4226
rect 20300 4172 20356 4174
rect 22204 6636 22260 6692
rect 22002 5514 22058 5516
rect 22002 5462 22004 5514
rect 22004 5462 22056 5514
rect 22056 5462 22058 5514
rect 22002 5460 22058 5462
rect 22106 5514 22162 5516
rect 22106 5462 22108 5514
rect 22108 5462 22160 5514
rect 22160 5462 22162 5514
rect 22106 5460 22162 5462
rect 22210 5514 22266 5516
rect 22210 5462 22212 5514
rect 22212 5462 22264 5514
rect 22264 5462 22266 5514
rect 22210 5460 22266 5462
rect 21868 4508 21924 4564
rect 21756 4284 21812 4340
rect 22540 7420 22596 7476
rect 23660 9996 23716 10052
rect 23324 7980 23380 8036
rect 22988 7474 23044 7476
rect 22988 7422 22990 7474
rect 22990 7422 23042 7474
rect 23042 7422 23044 7474
rect 22988 7420 23044 7422
rect 23324 6860 23380 6916
rect 22988 6578 23044 6580
rect 22988 6526 22990 6578
rect 22990 6526 23042 6578
rect 23042 6526 23044 6578
rect 22988 6524 23044 6526
rect 22988 6018 23044 6020
rect 22988 5966 22990 6018
rect 22990 5966 23042 6018
rect 23042 5966 23044 6018
rect 22988 5964 23044 5966
rect 22764 4956 22820 5012
rect 23548 6860 23604 6916
rect 23436 6748 23492 6804
rect 23772 8876 23828 8932
rect 24444 9714 24500 9716
rect 24444 9662 24446 9714
rect 24446 9662 24498 9714
rect 24498 9662 24500 9714
rect 24444 9660 24500 9662
rect 24668 10780 24724 10836
rect 26160 14138 26216 14140
rect 26160 14086 26162 14138
rect 26162 14086 26214 14138
rect 26214 14086 26216 14138
rect 26160 14084 26216 14086
rect 26264 14138 26320 14140
rect 26264 14086 26266 14138
rect 26266 14086 26318 14138
rect 26318 14086 26320 14138
rect 26264 14084 26320 14086
rect 26368 14138 26424 14140
rect 26368 14086 26370 14138
rect 26370 14086 26422 14138
rect 26422 14086 26424 14138
rect 26368 14084 26424 14086
rect 26796 13804 26852 13860
rect 26124 13746 26180 13748
rect 26124 13694 26126 13746
rect 26126 13694 26178 13746
rect 26178 13694 26180 13746
rect 26124 13692 26180 13694
rect 26460 13634 26516 13636
rect 26460 13582 26462 13634
rect 26462 13582 26514 13634
rect 26514 13582 26516 13634
rect 26460 13580 26516 13582
rect 26348 13356 26404 13412
rect 26160 12570 26216 12572
rect 26160 12518 26162 12570
rect 26162 12518 26214 12570
rect 26214 12518 26216 12570
rect 26160 12516 26216 12518
rect 26264 12570 26320 12572
rect 26264 12518 26266 12570
rect 26266 12518 26318 12570
rect 26318 12518 26320 12570
rect 26264 12516 26320 12518
rect 26368 12570 26424 12572
rect 26368 12518 26370 12570
rect 26370 12518 26422 12570
rect 26422 12518 26424 12570
rect 26368 12516 26424 12518
rect 25900 10668 25956 10724
rect 24668 9772 24724 9828
rect 23996 9266 24052 9268
rect 23996 9214 23998 9266
rect 23998 9214 24050 9266
rect 24050 9214 24052 9266
rect 23996 9212 24052 9214
rect 26684 12796 26740 12852
rect 26160 11002 26216 11004
rect 26160 10950 26162 11002
rect 26162 10950 26214 11002
rect 26214 10950 26216 11002
rect 26160 10948 26216 10950
rect 26264 11002 26320 11004
rect 26264 10950 26266 11002
rect 26266 10950 26318 11002
rect 26318 10950 26320 11002
rect 26264 10948 26320 10950
rect 26368 11002 26424 11004
rect 26368 10950 26370 11002
rect 26370 10950 26422 11002
rect 26422 10950 26424 11002
rect 26368 10948 26424 10950
rect 27020 13804 27076 13860
rect 27916 14700 27972 14756
rect 27468 13692 27524 13748
rect 27244 13634 27300 13636
rect 27244 13582 27246 13634
rect 27246 13582 27298 13634
rect 27298 13582 27300 13634
rect 27244 13580 27300 13582
rect 26908 13522 26964 13524
rect 26908 13470 26910 13522
rect 26910 13470 26962 13522
rect 26962 13470 26964 13522
rect 26908 13468 26964 13470
rect 27916 14476 27972 14532
rect 29372 19010 29428 19012
rect 29372 18958 29374 19010
rect 29374 18958 29426 19010
rect 29426 18958 29428 19010
rect 29372 18956 29428 18958
rect 30318 19626 30374 19628
rect 30318 19574 30320 19626
rect 30320 19574 30372 19626
rect 30372 19574 30374 19626
rect 30318 19572 30374 19574
rect 30422 19626 30478 19628
rect 30422 19574 30424 19626
rect 30424 19574 30476 19626
rect 30476 19574 30478 19626
rect 30422 19572 30478 19574
rect 30526 19626 30582 19628
rect 30526 19574 30528 19626
rect 30528 19574 30580 19626
rect 30580 19574 30582 19626
rect 30526 19572 30582 19574
rect 29372 17666 29428 17668
rect 29372 17614 29374 17666
rect 29374 17614 29426 17666
rect 29426 17614 29428 17666
rect 29372 17612 29428 17614
rect 29372 16994 29428 16996
rect 29372 16942 29374 16994
rect 29374 16942 29426 16994
rect 29426 16942 29428 16994
rect 29372 16940 29428 16942
rect 34476 18842 34532 18844
rect 34476 18790 34478 18842
rect 34478 18790 34530 18842
rect 34530 18790 34532 18842
rect 34476 18788 34532 18790
rect 34580 18842 34636 18844
rect 34580 18790 34582 18842
rect 34582 18790 34634 18842
rect 34634 18790 34636 18842
rect 34580 18788 34636 18790
rect 34684 18842 34740 18844
rect 34684 18790 34686 18842
rect 34686 18790 34738 18842
rect 34738 18790 34740 18842
rect 34684 18788 34740 18790
rect 30716 18562 30772 18564
rect 30716 18510 30718 18562
rect 30718 18510 30770 18562
rect 30770 18510 30772 18562
rect 30716 18508 30772 18510
rect 30318 18058 30374 18060
rect 30318 18006 30320 18058
rect 30320 18006 30372 18058
rect 30372 18006 30374 18058
rect 30318 18004 30374 18006
rect 30422 18058 30478 18060
rect 30422 18006 30424 18058
rect 30424 18006 30476 18058
rect 30476 18006 30478 18058
rect 30422 18004 30478 18006
rect 30526 18058 30582 18060
rect 30526 18006 30528 18058
rect 30528 18006 30580 18058
rect 30580 18006 30582 18058
rect 30526 18004 30582 18006
rect 29484 16828 29540 16884
rect 29820 16716 29876 16772
rect 29372 16098 29428 16100
rect 29372 16046 29374 16098
rect 29374 16046 29426 16098
rect 29426 16046 29428 16098
rect 29372 16044 29428 16046
rect 30380 16716 30436 16772
rect 30318 16490 30374 16492
rect 30318 16438 30320 16490
rect 30320 16438 30372 16490
rect 30372 16438 30374 16490
rect 30318 16436 30374 16438
rect 30422 16490 30478 16492
rect 30422 16438 30424 16490
rect 30424 16438 30476 16490
rect 30476 16438 30478 16490
rect 30422 16436 30478 16438
rect 30526 16490 30582 16492
rect 30526 16438 30528 16490
rect 30528 16438 30580 16490
rect 30580 16438 30582 16490
rect 30526 16436 30582 16438
rect 28924 15932 28980 15988
rect 28252 15148 28308 15204
rect 28028 13580 28084 13636
rect 27580 13356 27636 13412
rect 28812 15314 28868 15316
rect 28812 15262 28814 15314
rect 28814 15262 28866 15314
rect 28866 15262 28868 15314
rect 28812 15260 28868 15262
rect 28476 14700 28532 14756
rect 28028 12962 28084 12964
rect 28028 12910 28030 12962
rect 28030 12910 28082 12962
rect 28082 12910 28084 12962
rect 28028 12908 28084 12910
rect 28700 14476 28756 14532
rect 29148 14418 29204 14420
rect 29148 14366 29150 14418
rect 29150 14366 29202 14418
rect 29202 14366 29204 14418
rect 29148 14364 29204 14366
rect 31948 17724 32004 17780
rect 33292 17778 33348 17780
rect 33292 17726 33294 17778
rect 33294 17726 33346 17778
rect 33346 17726 33348 17778
rect 33292 17724 33348 17726
rect 34476 17274 34532 17276
rect 34476 17222 34478 17274
rect 34478 17222 34530 17274
rect 34530 17222 34532 17274
rect 34476 17220 34532 17222
rect 34580 17274 34636 17276
rect 34580 17222 34582 17274
rect 34582 17222 34634 17274
rect 34634 17222 34636 17274
rect 34580 17220 34636 17222
rect 34684 17274 34740 17276
rect 34684 17222 34686 17274
rect 34686 17222 34738 17274
rect 34738 17222 34740 17274
rect 34684 17220 34740 17222
rect 31500 16716 31556 16772
rect 31164 15708 31220 15764
rect 30380 15538 30436 15540
rect 30380 15486 30382 15538
rect 30382 15486 30434 15538
rect 30434 15486 30436 15538
rect 30380 15484 30436 15486
rect 30940 15426 30996 15428
rect 30940 15374 30942 15426
rect 30942 15374 30994 15426
rect 30994 15374 30996 15426
rect 30940 15372 30996 15374
rect 31388 15372 31444 15428
rect 30604 15202 30660 15204
rect 30604 15150 30606 15202
rect 30606 15150 30658 15202
rect 30658 15150 30660 15202
rect 30604 15148 30660 15150
rect 30492 15036 30548 15092
rect 30318 14922 30374 14924
rect 30318 14870 30320 14922
rect 30320 14870 30372 14922
rect 30372 14870 30374 14922
rect 30318 14868 30374 14870
rect 30422 14922 30478 14924
rect 30422 14870 30424 14922
rect 30424 14870 30476 14922
rect 30476 14870 30478 14922
rect 30422 14868 30478 14870
rect 30526 14922 30582 14924
rect 30526 14870 30528 14922
rect 30528 14870 30580 14922
rect 30580 14870 30582 14922
rect 30526 14868 30582 14870
rect 31500 15314 31556 15316
rect 31500 15262 31502 15314
rect 31502 15262 31554 15314
rect 31554 15262 31556 15314
rect 31500 15260 31556 15262
rect 32284 15708 32340 15764
rect 30044 14364 30100 14420
rect 32508 15148 32564 15204
rect 32172 14754 32228 14756
rect 32172 14702 32174 14754
rect 32174 14702 32226 14754
rect 32226 14702 32228 14754
rect 32172 14700 32228 14702
rect 29596 13186 29652 13188
rect 29596 13134 29598 13186
rect 29598 13134 29650 13186
rect 29650 13134 29652 13186
rect 29596 13132 29652 13134
rect 29372 12962 29428 12964
rect 29372 12910 29374 12962
rect 29374 12910 29426 12962
rect 29426 12910 29428 12962
rect 29372 12908 29428 12910
rect 30318 13354 30374 13356
rect 30318 13302 30320 13354
rect 30320 13302 30372 13354
rect 30372 13302 30374 13354
rect 30318 13300 30374 13302
rect 30422 13354 30478 13356
rect 30422 13302 30424 13354
rect 30424 13302 30476 13354
rect 30476 13302 30478 13354
rect 30422 13300 30478 13302
rect 30526 13354 30582 13356
rect 30526 13302 30528 13354
rect 30528 13302 30580 13354
rect 30580 13302 30582 13354
rect 30526 13300 30582 13302
rect 30318 11786 30374 11788
rect 30318 11734 30320 11786
rect 30320 11734 30372 11786
rect 30372 11734 30374 11786
rect 30318 11732 30374 11734
rect 30422 11786 30478 11788
rect 30422 11734 30424 11786
rect 30424 11734 30476 11786
rect 30476 11734 30478 11786
rect 30422 11732 30478 11734
rect 30526 11786 30582 11788
rect 30526 11734 30528 11786
rect 30528 11734 30580 11786
rect 30580 11734 30582 11786
rect 30526 11732 30582 11734
rect 26908 9996 26964 10052
rect 27132 9996 27188 10052
rect 27804 9884 27860 9940
rect 26796 9660 26852 9716
rect 26160 9434 26216 9436
rect 26160 9382 26162 9434
rect 26162 9382 26214 9434
rect 26214 9382 26216 9434
rect 26160 9380 26216 9382
rect 26264 9434 26320 9436
rect 26264 9382 26266 9434
rect 26266 9382 26318 9434
rect 26318 9382 26320 9434
rect 26264 9380 26320 9382
rect 26368 9434 26424 9436
rect 26368 9382 26370 9434
rect 26370 9382 26422 9434
rect 26422 9382 26424 9434
rect 26368 9380 26424 9382
rect 27244 9826 27300 9828
rect 27244 9774 27246 9826
rect 27246 9774 27298 9826
rect 27298 9774 27300 9826
rect 27244 9772 27300 9774
rect 27916 9548 27972 9604
rect 25340 8930 25396 8932
rect 25340 8878 25342 8930
rect 25342 8878 25394 8930
rect 25394 8878 25396 8930
rect 25340 8876 25396 8878
rect 23772 7196 23828 7252
rect 25900 8204 25956 8260
rect 26908 8258 26964 8260
rect 26908 8206 26910 8258
rect 26910 8206 26962 8258
rect 26962 8206 26964 8258
rect 26908 8204 26964 8206
rect 26160 7866 26216 7868
rect 26160 7814 26162 7866
rect 26162 7814 26214 7866
rect 26214 7814 26216 7866
rect 26160 7812 26216 7814
rect 26264 7866 26320 7868
rect 26264 7814 26266 7866
rect 26266 7814 26318 7866
rect 26318 7814 26320 7866
rect 26264 7812 26320 7814
rect 26368 7866 26424 7868
rect 26368 7814 26370 7866
rect 26370 7814 26422 7866
rect 26422 7814 26424 7866
rect 26368 7812 26424 7814
rect 24108 7196 24164 7252
rect 23660 6636 23716 6692
rect 24780 6578 24836 6580
rect 24780 6526 24782 6578
rect 24782 6526 24834 6578
rect 24834 6526 24836 6578
rect 24780 6524 24836 6526
rect 24220 5964 24276 6020
rect 24108 5852 24164 5908
rect 22002 3946 22058 3948
rect 22002 3894 22004 3946
rect 22004 3894 22056 3946
rect 22056 3894 22058 3946
rect 22002 3892 22058 3894
rect 22106 3946 22162 3948
rect 22106 3894 22108 3946
rect 22108 3894 22160 3946
rect 22160 3894 22162 3946
rect 22106 3892 22162 3894
rect 22210 3946 22266 3948
rect 22210 3894 22212 3946
rect 22212 3894 22264 3946
rect 22264 3894 22266 3946
rect 22210 3892 22266 3894
rect 20748 3554 20804 3556
rect 20748 3502 20750 3554
rect 20750 3502 20802 3554
rect 20802 3502 20804 3554
rect 20748 3500 20804 3502
rect 22764 4562 22820 4564
rect 22764 4510 22766 4562
rect 22766 4510 22818 4562
rect 22818 4510 22820 4562
rect 22764 4508 22820 4510
rect 23100 4338 23156 4340
rect 23100 4286 23102 4338
rect 23102 4286 23154 4338
rect 23154 4286 23156 4338
rect 23100 4284 23156 4286
rect 23772 5180 23828 5236
rect 23436 4956 23492 5012
rect 23324 4060 23380 4116
rect 22764 3612 22820 3668
rect 25340 6524 25396 6580
rect 26236 7474 26292 7476
rect 26236 7422 26238 7474
rect 26238 7422 26290 7474
rect 26290 7422 26292 7474
rect 26236 7420 26292 7422
rect 26012 6860 26068 6916
rect 26684 6748 26740 6804
rect 26460 6690 26516 6692
rect 26460 6638 26462 6690
rect 26462 6638 26514 6690
rect 26514 6638 26516 6690
rect 26460 6636 26516 6638
rect 26160 6298 26216 6300
rect 26160 6246 26162 6298
rect 26162 6246 26214 6298
rect 26214 6246 26216 6298
rect 26160 6244 26216 6246
rect 26264 6298 26320 6300
rect 26264 6246 26266 6298
rect 26266 6246 26318 6298
rect 26318 6246 26320 6298
rect 26264 6244 26320 6246
rect 26368 6298 26424 6300
rect 26368 6246 26370 6298
rect 26370 6246 26422 6298
rect 26422 6246 26424 6298
rect 26368 6244 26424 6246
rect 25452 6018 25508 6020
rect 25452 5966 25454 6018
rect 25454 5966 25506 6018
rect 25506 5966 25508 6018
rect 25452 5964 25508 5966
rect 25228 5906 25284 5908
rect 25228 5854 25230 5906
rect 25230 5854 25282 5906
rect 25282 5854 25284 5906
rect 25228 5852 25284 5854
rect 24332 5794 24388 5796
rect 24332 5742 24334 5794
rect 24334 5742 24386 5794
rect 24386 5742 24388 5794
rect 24332 5740 24388 5742
rect 25564 5740 25620 5796
rect 23660 4226 23716 4228
rect 23660 4174 23662 4226
rect 23662 4174 23714 4226
rect 23714 4174 23716 4226
rect 23660 4172 23716 4174
rect 27692 7308 27748 7364
rect 27244 6524 27300 6580
rect 27692 7084 27748 7140
rect 26908 5964 26964 6020
rect 26796 5852 26852 5908
rect 28028 8146 28084 8148
rect 28028 8094 28030 8146
rect 28030 8094 28082 8146
rect 28082 8094 28084 8146
rect 28028 8092 28084 8094
rect 28028 7250 28084 7252
rect 28028 7198 28030 7250
rect 28030 7198 28082 7250
rect 28082 7198 28084 7250
rect 28028 7196 28084 7198
rect 29148 9772 29204 9828
rect 29372 9714 29428 9716
rect 29372 9662 29374 9714
rect 29374 9662 29426 9714
rect 29426 9662 29428 9714
rect 29372 9660 29428 9662
rect 29484 9884 29540 9940
rect 28476 9602 28532 9604
rect 28476 9550 28478 9602
rect 28478 9550 28530 9602
rect 28530 9550 28532 9602
rect 28476 9548 28532 9550
rect 29260 9548 29316 9604
rect 28252 7084 28308 7140
rect 29148 7308 29204 7364
rect 28700 6748 28756 6804
rect 26012 5794 26068 5796
rect 26012 5742 26014 5794
rect 26014 5742 26066 5794
rect 26066 5742 26068 5794
rect 26012 5740 26068 5742
rect 26796 5682 26852 5684
rect 26796 5630 26798 5682
rect 26798 5630 26850 5682
rect 26850 5630 26852 5682
rect 26796 5628 26852 5630
rect 26908 5180 26964 5236
rect 27020 5122 27076 5124
rect 27020 5070 27022 5122
rect 27022 5070 27074 5122
rect 27074 5070 27076 5122
rect 27020 5068 27076 5070
rect 26236 5010 26292 5012
rect 26236 4958 26238 5010
rect 26238 4958 26290 5010
rect 26290 4958 26292 5010
rect 26236 4956 26292 4958
rect 26160 4730 26216 4732
rect 26160 4678 26162 4730
rect 26162 4678 26214 4730
rect 26214 4678 26216 4730
rect 26160 4676 26216 4678
rect 26264 4730 26320 4732
rect 26264 4678 26266 4730
rect 26266 4678 26318 4730
rect 26318 4678 26320 4730
rect 26264 4676 26320 4678
rect 26368 4730 26424 4732
rect 26368 4678 26370 4730
rect 26370 4678 26422 4730
rect 26422 4678 26424 4730
rect 26368 4676 26424 4678
rect 27468 5906 27524 5908
rect 27468 5854 27470 5906
rect 27470 5854 27522 5906
rect 27522 5854 27524 5906
rect 27468 5852 27524 5854
rect 27580 5794 27636 5796
rect 27580 5742 27582 5794
rect 27582 5742 27634 5794
rect 27634 5742 27636 5794
rect 27580 5740 27636 5742
rect 29708 9826 29764 9828
rect 29708 9774 29710 9826
rect 29710 9774 29762 9826
rect 29762 9774 29764 9826
rect 29708 9772 29764 9774
rect 29708 8428 29764 8484
rect 29372 8146 29428 8148
rect 29372 8094 29374 8146
rect 29374 8094 29426 8146
rect 29426 8094 29428 8146
rect 29372 8092 29428 8094
rect 29708 8258 29764 8260
rect 29708 8206 29710 8258
rect 29710 8206 29762 8258
rect 29762 8206 29764 8258
rect 29708 8204 29764 8206
rect 29932 10498 29988 10500
rect 29932 10446 29934 10498
rect 29934 10446 29986 10498
rect 29986 10446 29988 10498
rect 29932 10444 29988 10446
rect 29932 10220 29988 10276
rect 29932 9772 29988 9828
rect 30380 10610 30436 10612
rect 30380 10558 30382 10610
rect 30382 10558 30434 10610
rect 30434 10558 30436 10610
rect 30380 10556 30436 10558
rect 30268 10444 30324 10500
rect 30492 10332 30548 10388
rect 30318 10218 30374 10220
rect 30318 10166 30320 10218
rect 30320 10166 30372 10218
rect 30372 10166 30374 10218
rect 30318 10164 30374 10166
rect 30422 10218 30478 10220
rect 30422 10166 30424 10218
rect 30424 10166 30476 10218
rect 30476 10166 30478 10218
rect 30422 10164 30478 10166
rect 30526 10218 30582 10220
rect 30526 10166 30528 10218
rect 30528 10166 30580 10218
rect 30580 10166 30582 10218
rect 30526 10164 30582 10166
rect 31276 13468 31332 13524
rect 32060 14476 32116 14532
rect 30940 10668 30996 10724
rect 30828 10444 30884 10500
rect 32732 14924 32788 14980
rect 34476 15706 34532 15708
rect 34476 15654 34478 15706
rect 34478 15654 34530 15706
rect 34530 15654 34532 15706
rect 34476 15652 34532 15654
rect 34580 15706 34636 15708
rect 34580 15654 34582 15706
rect 34582 15654 34634 15706
rect 34634 15654 34636 15706
rect 34580 15652 34636 15654
rect 34684 15706 34740 15708
rect 34684 15654 34686 15706
rect 34686 15654 34738 15706
rect 34738 15654 34740 15706
rect 34684 15652 34740 15654
rect 33628 15372 33684 15428
rect 33180 15148 33236 15204
rect 33068 14530 33124 14532
rect 33068 14478 33070 14530
rect 33070 14478 33122 14530
rect 33122 14478 33124 14530
rect 33068 14476 33124 14478
rect 32396 13580 32452 13636
rect 31836 13132 31892 13188
rect 31948 11954 32004 11956
rect 31948 11902 31950 11954
rect 31950 11902 32002 11954
rect 32002 11902 32004 11954
rect 31948 11900 32004 11902
rect 31836 10722 31892 10724
rect 31836 10670 31838 10722
rect 31838 10670 31890 10722
rect 31890 10670 31892 10722
rect 31836 10668 31892 10670
rect 31164 10332 31220 10388
rect 31276 10556 31332 10612
rect 30716 9996 30772 10052
rect 30380 9826 30436 9828
rect 30380 9774 30382 9826
rect 30382 9774 30434 9826
rect 30434 9774 30436 9826
rect 30380 9772 30436 9774
rect 30156 9660 30212 9716
rect 30940 9884 30996 9940
rect 30716 9100 30772 9156
rect 30318 8650 30374 8652
rect 30318 8598 30320 8650
rect 30320 8598 30372 8650
rect 30372 8598 30374 8650
rect 30318 8596 30374 8598
rect 30422 8650 30478 8652
rect 30422 8598 30424 8650
rect 30424 8598 30476 8650
rect 30476 8598 30478 8650
rect 30422 8596 30478 8598
rect 30526 8650 30582 8652
rect 30526 8598 30528 8650
rect 30528 8598 30580 8650
rect 30580 8598 30582 8650
rect 30526 8596 30582 8598
rect 30380 8428 30436 8484
rect 31388 9100 31444 9156
rect 30492 8258 30548 8260
rect 30492 8206 30494 8258
rect 30494 8206 30546 8258
rect 30546 8206 30548 8258
rect 30492 8204 30548 8206
rect 29484 7586 29540 7588
rect 29484 7534 29486 7586
rect 29486 7534 29538 7586
rect 29538 7534 29540 7586
rect 29484 7532 29540 7534
rect 29260 7196 29316 7252
rect 27804 5234 27860 5236
rect 27804 5182 27806 5234
rect 27806 5182 27858 5234
rect 27858 5182 27860 5234
rect 27804 5180 27860 5182
rect 28700 4956 28756 5012
rect 27468 4898 27524 4900
rect 27468 4846 27470 4898
rect 27470 4846 27522 4898
rect 27522 4846 27524 4898
rect 27468 4844 27524 4846
rect 29372 6802 29428 6804
rect 29372 6750 29374 6802
rect 29374 6750 29426 6802
rect 29426 6750 29428 6802
rect 29372 6748 29428 6750
rect 29708 6802 29764 6804
rect 29708 6750 29710 6802
rect 29710 6750 29762 6802
rect 29762 6750 29764 6802
rect 29708 6748 29764 6750
rect 30268 7474 30324 7476
rect 30268 7422 30270 7474
rect 30270 7422 30322 7474
rect 30322 7422 30324 7474
rect 30268 7420 30324 7422
rect 31052 7474 31108 7476
rect 31052 7422 31054 7474
rect 31054 7422 31106 7474
rect 31106 7422 31108 7474
rect 31052 7420 31108 7422
rect 30318 7082 30374 7084
rect 30318 7030 30320 7082
rect 30320 7030 30372 7082
rect 30372 7030 30374 7082
rect 30318 7028 30374 7030
rect 30422 7082 30478 7084
rect 30422 7030 30424 7082
rect 30424 7030 30476 7082
rect 30476 7030 30478 7082
rect 30422 7028 30478 7030
rect 30526 7082 30582 7084
rect 30526 7030 30528 7082
rect 30528 7030 30580 7082
rect 30580 7030 30582 7082
rect 30526 7028 30582 7030
rect 29932 6636 29988 6692
rect 29932 6188 29988 6244
rect 30044 6748 30100 6804
rect 29820 5852 29876 5908
rect 30156 6188 30212 6244
rect 30716 6860 30772 6916
rect 30380 6802 30436 6804
rect 30380 6750 30382 6802
rect 30382 6750 30434 6802
rect 30434 6750 30436 6802
rect 30380 6748 30436 6750
rect 32172 10610 32228 10612
rect 32172 10558 32174 10610
rect 32174 10558 32226 10610
rect 32226 10558 32228 10610
rect 32172 10556 32228 10558
rect 31836 9154 31892 9156
rect 31836 9102 31838 9154
rect 31838 9102 31890 9154
rect 31890 9102 31892 9154
rect 31836 9100 31892 9102
rect 32172 8988 32228 9044
rect 31724 7420 31780 7476
rect 31724 7250 31780 7252
rect 31724 7198 31726 7250
rect 31726 7198 31778 7250
rect 31778 7198 31780 7250
rect 31724 7196 31780 7198
rect 31612 6860 31668 6916
rect 30940 6018 30996 6020
rect 30940 5966 30942 6018
rect 30942 5966 30994 6018
rect 30994 5966 30996 6018
rect 30940 5964 30996 5966
rect 30318 5514 30374 5516
rect 30318 5462 30320 5514
rect 30320 5462 30372 5514
rect 30372 5462 30374 5514
rect 30318 5460 30374 5462
rect 30422 5514 30478 5516
rect 30422 5462 30424 5514
rect 30424 5462 30476 5514
rect 30476 5462 30478 5514
rect 30422 5460 30478 5462
rect 30526 5514 30582 5516
rect 30526 5462 30528 5514
rect 30528 5462 30580 5514
rect 30580 5462 30582 5514
rect 30526 5460 30582 5462
rect 30604 5180 30660 5236
rect 29708 5122 29764 5124
rect 29708 5070 29710 5122
rect 29710 5070 29762 5122
rect 29762 5070 29764 5122
rect 29708 5068 29764 5070
rect 30380 5122 30436 5124
rect 30380 5070 30382 5122
rect 30382 5070 30434 5122
rect 30434 5070 30436 5122
rect 30380 5068 30436 5070
rect 31164 5906 31220 5908
rect 31164 5854 31166 5906
rect 31166 5854 31218 5906
rect 31218 5854 31220 5906
rect 31164 5852 31220 5854
rect 31724 5794 31780 5796
rect 31724 5742 31726 5794
rect 31726 5742 31778 5794
rect 31778 5742 31780 5794
rect 31724 5740 31780 5742
rect 31836 5180 31892 5236
rect 31276 4956 31332 5012
rect 31948 4956 32004 5012
rect 29596 4898 29652 4900
rect 29596 4846 29598 4898
rect 29598 4846 29650 4898
rect 29650 4846 29652 4898
rect 29596 4844 29652 4846
rect 31164 4844 31220 4900
rect 25228 4060 25284 4116
rect 24556 3666 24612 3668
rect 24556 3614 24558 3666
rect 24558 3614 24610 3666
rect 24610 3614 24612 3666
rect 24556 3612 24612 3614
rect 22428 3500 22484 3556
rect 24892 3554 24948 3556
rect 24892 3502 24894 3554
rect 24894 3502 24946 3554
rect 24946 3502 24948 3554
rect 24892 3500 24948 3502
rect 30318 3946 30374 3948
rect 30318 3894 30320 3946
rect 30320 3894 30372 3946
rect 30372 3894 30374 3946
rect 30318 3892 30374 3894
rect 30422 3946 30478 3948
rect 30422 3894 30424 3946
rect 30424 3894 30476 3946
rect 30476 3894 30478 3946
rect 30422 3892 30478 3894
rect 30526 3946 30582 3948
rect 30526 3894 30528 3946
rect 30528 3894 30580 3946
rect 30580 3894 30582 3946
rect 30526 3892 30582 3894
rect 34476 14138 34532 14140
rect 34476 14086 34478 14138
rect 34478 14086 34530 14138
rect 34530 14086 34532 14138
rect 34476 14084 34532 14086
rect 34580 14138 34636 14140
rect 34580 14086 34582 14138
rect 34582 14086 34634 14138
rect 34634 14086 34636 14138
rect 34580 14084 34636 14086
rect 34684 14138 34740 14140
rect 34684 14086 34686 14138
rect 34686 14086 34738 14138
rect 34738 14086 34740 14138
rect 34684 14084 34740 14086
rect 33068 13580 33124 13636
rect 33292 13522 33348 13524
rect 33292 13470 33294 13522
rect 33294 13470 33346 13522
rect 33346 13470 33348 13522
rect 33292 13468 33348 13470
rect 33516 13522 33572 13524
rect 33516 13470 33518 13522
rect 33518 13470 33570 13522
rect 33570 13470 33572 13522
rect 33516 13468 33572 13470
rect 33292 11900 33348 11956
rect 34476 12570 34532 12572
rect 34476 12518 34478 12570
rect 34478 12518 34530 12570
rect 34530 12518 34532 12570
rect 34476 12516 34532 12518
rect 34580 12570 34636 12572
rect 34580 12518 34582 12570
rect 34582 12518 34634 12570
rect 34634 12518 34636 12570
rect 34580 12516 34636 12518
rect 34684 12570 34740 12572
rect 34684 12518 34686 12570
rect 34686 12518 34738 12570
rect 34738 12518 34740 12570
rect 34684 12516 34740 12518
rect 33068 9884 33124 9940
rect 34476 11002 34532 11004
rect 34476 10950 34478 11002
rect 34478 10950 34530 11002
rect 34530 10950 34532 11002
rect 34476 10948 34532 10950
rect 34580 11002 34636 11004
rect 34580 10950 34582 11002
rect 34582 10950 34634 11002
rect 34634 10950 34636 11002
rect 34580 10948 34636 10950
rect 34684 11002 34740 11004
rect 34684 10950 34686 11002
rect 34686 10950 34738 11002
rect 34738 10950 34740 11002
rect 34684 10948 34740 10950
rect 34476 9434 34532 9436
rect 34476 9382 34478 9434
rect 34478 9382 34530 9434
rect 34530 9382 34532 9434
rect 34476 9380 34532 9382
rect 34580 9434 34636 9436
rect 34580 9382 34582 9434
rect 34582 9382 34634 9434
rect 34634 9382 34636 9434
rect 34580 9380 34636 9382
rect 34684 9434 34740 9436
rect 34684 9382 34686 9434
rect 34686 9382 34738 9434
rect 34738 9382 34740 9434
rect 34684 9380 34740 9382
rect 34076 9100 34132 9156
rect 33292 9042 33348 9044
rect 33292 8990 33294 9042
rect 33294 8990 33346 9042
rect 33346 8990 33348 9042
rect 33292 8988 33348 8990
rect 33404 8316 33460 8372
rect 33404 7532 33460 7588
rect 34188 8370 34244 8372
rect 34188 8318 34190 8370
rect 34190 8318 34242 8370
rect 34242 8318 34244 8370
rect 34188 8316 34244 8318
rect 34476 7866 34532 7868
rect 34476 7814 34478 7866
rect 34478 7814 34530 7866
rect 34530 7814 34532 7866
rect 34476 7812 34532 7814
rect 34580 7866 34636 7868
rect 34580 7814 34582 7866
rect 34582 7814 34634 7866
rect 34634 7814 34636 7866
rect 34580 7812 34636 7814
rect 34684 7866 34740 7868
rect 34684 7814 34686 7866
rect 34686 7814 34738 7866
rect 34738 7814 34740 7866
rect 34684 7812 34740 7814
rect 33516 7196 33572 7252
rect 33068 6860 33124 6916
rect 33068 6188 33124 6244
rect 32956 5906 33012 5908
rect 32956 5854 32958 5906
rect 32958 5854 33010 5906
rect 33010 5854 33012 5906
rect 32956 5852 33012 5854
rect 34476 6298 34532 6300
rect 34476 6246 34478 6298
rect 34478 6246 34530 6298
rect 34530 6246 34532 6298
rect 34476 6244 34532 6246
rect 34580 6298 34636 6300
rect 34580 6246 34582 6298
rect 34582 6246 34634 6298
rect 34634 6246 34636 6298
rect 34580 6244 34636 6246
rect 34684 6298 34740 6300
rect 34684 6246 34686 6298
rect 34686 6246 34738 6298
rect 34738 6246 34740 6298
rect 34684 6244 34740 6246
rect 33404 6018 33460 6020
rect 33404 5966 33406 6018
rect 33406 5966 33458 6018
rect 33458 5966 33460 6018
rect 33404 5964 33460 5966
rect 33180 5794 33236 5796
rect 33180 5742 33182 5794
rect 33182 5742 33234 5794
rect 33234 5742 33236 5794
rect 33180 5740 33236 5742
rect 33516 5180 33572 5236
rect 34188 5234 34244 5236
rect 34188 5182 34190 5234
rect 34190 5182 34242 5234
rect 34242 5182 34244 5234
rect 34188 5180 34244 5182
rect 34476 4730 34532 4732
rect 34476 4678 34478 4730
rect 34478 4678 34530 4730
rect 34530 4678 34532 4730
rect 34476 4676 34532 4678
rect 34580 4730 34636 4732
rect 34580 4678 34582 4730
rect 34582 4678 34634 4730
rect 34634 4678 34636 4730
rect 34580 4676 34636 4678
rect 34684 4730 34740 4732
rect 34684 4678 34686 4730
rect 34686 4678 34738 4730
rect 34738 4678 34740 4730
rect 34684 4676 34740 4678
rect 31500 3554 31556 3556
rect 31500 3502 31502 3554
rect 31502 3502 31554 3554
rect 31554 3502 31556 3554
rect 31500 3500 31556 3502
rect 25116 3388 25172 3444
rect 26908 3442 26964 3444
rect 26908 3390 26910 3442
rect 26910 3390 26962 3442
rect 26962 3390 26964 3442
rect 26908 3388 26964 3390
rect 32172 3500 32228 3556
rect 30044 3442 30100 3444
rect 30044 3390 30046 3442
rect 30046 3390 30098 3442
rect 30098 3390 30100 3442
rect 30044 3388 30100 3390
rect 32284 3388 32340 3444
rect 26160 3162 26216 3164
rect 26160 3110 26162 3162
rect 26162 3110 26214 3162
rect 26214 3110 26216 3162
rect 26160 3108 26216 3110
rect 26264 3162 26320 3164
rect 26264 3110 26266 3162
rect 26266 3110 26318 3162
rect 26318 3110 26320 3162
rect 26264 3108 26320 3110
rect 26368 3162 26424 3164
rect 26368 3110 26370 3162
rect 26370 3110 26422 3162
rect 26422 3110 26424 3162
rect 26368 3108 26424 3110
rect 34476 3162 34532 3164
rect 34476 3110 34478 3162
rect 34478 3110 34530 3162
rect 34530 3110 34532 3162
rect 34476 3108 34532 3110
rect 34580 3162 34636 3164
rect 34580 3110 34582 3162
rect 34582 3110 34634 3162
rect 34634 3110 34636 3162
rect 34580 3108 34636 3110
rect 34684 3162 34740 3164
rect 34684 3110 34686 3162
rect 34686 3110 34738 3162
rect 34738 3110 34740 3162
rect 34684 3108 34740 3110
<< metal3 >>
rect 5360 32116 5370 32172
rect 5426 32116 5474 32172
rect 5530 32116 5578 32172
rect 5634 32116 5644 32172
rect 13676 32116 13686 32172
rect 13742 32116 13790 32172
rect 13846 32116 13894 32172
rect 13950 32116 13960 32172
rect 21992 32116 22002 32172
rect 22058 32116 22106 32172
rect 22162 32116 22210 32172
rect 22266 32116 22276 32172
rect 30308 32116 30318 32172
rect 30374 32116 30422 32172
rect 30478 32116 30526 32172
rect 30582 32116 30592 32172
rect 9518 31332 9528 31388
rect 9584 31332 9632 31388
rect 9688 31332 9736 31388
rect 9792 31332 9802 31388
rect 17834 31332 17844 31388
rect 17900 31332 17948 31388
rect 18004 31332 18052 31388
rect 18108 31332 18118 31388
rect 26150 31332 26160 31388
rect 26216 31332 26264 31388
rect 26320 31332 26368 31388
rect 26424 31332 26434 31388
rect 34466 31332 34476 31388
rect 34532 31332 34580 31388
rect 34636 31332 34684 31388
rect 34740 31332 34750 31388
rect 5360 30548 5370 30604
rect 5426 30548 5474 30604
rect 5530 30548 5578 30604
rect 5634 30548 5644 30604
rect 13676 30548 13686 30604
rect 13742 30548 13790 30604
rect 13846 30548 13894 30604
rect 13950 30548 13960 30604
rect 21992 30548 22002 30604
rect 22058 30548 22106 30604
rect 22162 30548 22210 30604
rect 22266 30548 22276 30604
rect 30308 30548 30318 30604
rect 30374 30548 30422 30604
rect 30478 30548 30526 30604
rect 30582 30548 30592 30604
rect 9518 29764 9528 29820
rect 9584 29764 9632 29820
rect 9688 29764 9736 29820
rect 9792 29764 9802 29820
rect 17834 29764 17844 29820
rect 17900 29764 17948 29820
rect 18004 29764 18052 29820
rect 18108 29764 18118 29820
rect 26150 29764 26160 29820
rect 26216 29764 26264 29820
rect 26320 29764 26368 29820
rect 26424 29764 26434 29820
rect 34466 29764 34476 29820
rect 34532 29764 34580 29820
rect 34636 29764 34684 29820
rect 34740 29764 34750 29820
rect 5360 28980 5370 29036
rect 5426 28980 5474 29036
rect 5530 28980 5578 29036
rect 5634 28980 5644 29036
rect 13676 28980 13686 29036
rect 13742 28980 13790 29036
rect 13846 28980 13894 29036
rect 13950 28980 13960 29036
rect 21992 28980 22002 29036
rect 22058 28980 22106 29036
rect 22162 28980 22210 29036
rect 22266 28980 22276 29036
rect 30308 28980 30318 29036
rect 30374 28980 30422 29036
rect 30478 28980 30526 29036
rect 30582 28980 30592 29036
rect 9518 28196 9528 28252
rect 9584 28196 9632 28252
rect 9688 28196 9736 28252
rect 9792 28196 9802 28252
rect 17834 28196 17844 28252
rect 17900 28196 17948 28252
rect 18004 28196 18052 28252
rect 18108 28196 18118 28252
rect 26150 28196 26160 28252
rect 26216 28196 26264 28252
rect 26320 28196 26368 28252
rect 26424 28196 26434 28252
rect 34466 28196 34476 28252
rect 34532 28196 34580 28252
rect 34636 28196 34684 28252
rect 34740 28196 34750 28252
rect 8418 27804 8428 27860
rect 8484 27804 10220 27860
rect 10276 27804 10286 27860
rect 19058 27804 19068 27860
rect 19124 27804 20188 27860
rect 20244 27804 20254 27860
rect 10994 27692 11004 27748
rect 11060 27692 12236 27748
rect 12292 27692 12302 27748
rect 5360 27412 5370 27468
rect 5426 27412 5474 27468
rect 5530 27412 5578 27468
rect 5634 27412 5644 27468
rect 13676 27412 13686 27468
rect 13742 27412 13790 27468
rect 13846 27412 13894 27468
rect 13950 27412 13960 27468
rect 21992 27412 22002 27468
rect 22058 27412 22106 27468
rect 22162 27412 22210 27468
rect 22266 27412 22276 27468
rect 30308 27412 30318 27468
rect 30374 27412 30422 27468
rect 30478 27412 30526 27468
rect 30582 27412 30592 27468
rect 5170 27244 5180 27300
rect 5236 27244 5852 27300
rect 5908 27244 5918 27300
rect 5180 27076 5236 27244
rect 16370 27132 16380 27188
rect 16436 27132 17164 27188
rect 17220 27132 17230 27188
rect 4956 27020 5236 27076
rect 5954 27020 5964 27076
rect 6020 27020 6748 27076
rect 6804 27020 6814 27076
rect 12450 27020 12460 27076
rect 12516 27020 17724 27076
rect 17780 27020 17790 27076
rect 4956 26964 5012 27020
rect 4946 26908 4956 26964
rect 5012 26908 5022 26964
rect 5170 26908 5180 26964
rect 5236 26908 6412 26964
rect 6468 26908 6860 26964
rect 6916 26908 6926 26964
rect 14354 26908 14364 26964
rect 14420 26908 15484 26964
rect 15540 26908 15550 26964
rect 17714 26796 17724 26852
rect 17780 26796 20524 26852
rect 20580 26796 20590 26852
rect 9518 26628 9528 26684
rect 9584 26628 9632 26684
rect 9688 26628 9736 26684
rect 9792 26628 9802 26684
rect 17834 26628 17844 26684
rect 17900 26628 17948 26684
rect 18004 26628 18052 26684
rect 18108 26628 18118 26684
rect 26150 26628 26160 26684
rect 26216 26628 26264 26684
rect 26320 26628 26368 26684
rect 26424 26628 26434 26684
rect 34466 26628 34476 26684
rect 34532 26628 34580 26684
rect 34636 26628 34684 26684
rect 34740 26628 34750 26684
rect 18946 26572 18956 26628
rect 19012 26572 20412 26628
rect 20468 26572 22652 26628
rect 22708 26572 22718 26628
rect 8194 26460 8204 26516
rect 8260 26460 8876 26516
rect 8932 26460 8942 26516
rect 2482 26348 2492 26404
rect 2548 26348 3276 26404
rect 3332 26348 3342 26404
rect 6290 26348 6300 26404
rect 6356 26348 7308 26404
rect 7364 26348 7374 26404
rect 12338 26236 12348 26292
rect 12404 26236 13132 26292
rect 13188 26236 13198 26292
rect 15698 26236 15708 26292
rect 15764 26236 16380 26292
rect 16436 26236 16446 26292
rect 18274 26236 18284 26292
rect 18340 26236 18844 26292
rect 18900 26236 18910 26292
rect 17602 26124 17612 26180
rect 17668 26124 19628 26180
rect 19684 26124 19694 26180
rect 22530 26124 22540 26180
rect 22596 26124 24108 26180
rect 24164 26124 24174 26180
rect 5360 25844 5370 25900
rect 5426 25844 5474 25900
rect 5530 25844 5578 25900
rect 5634 25844 5644 25900
rect 13676 25844 13686 25900
rect 13742 25844 13790 25900
rect 13846 25844 13894 25900
rect 13950 25844 13960 25900
rect 21992 25844 22002 25900
rect 22058 25844 22106 25900
rect 22162 25844 22210 25900
rect 22266 25844 22276 25900
rect 30308 25844 30318 25900
rect 30374 25844 30422 25900
rect 30478 25844 30526 25900
rect 30582 25844 30592 25900
rect 14130 25788 14140 25844
rect 14196 25788 16604 25844
rect 16660 25788 16670 25844
rect 10994 25676 11004 25732
rect 11060 25676 14756 25732
rect 19282 25676 19292 25732
rect 19348 25676 23436 25732
rect 23492 25676 23502 25732
rect 12674 25564 12684 25620
rect 12740 25564 13580 25620
rect 13636 25564 13646 25620
rect 14700 25508 14756 25676
rect 1810 25452 1820 25508
rect 1876 25452 7084 25508
rect 7140 25452 7420 25508
rect 7476 25452 7980 25508
rect 8036 25452 8046 25508
rect 12002 25452 12012 25508
rect 12068 25452 12348 25508
rect 12404 25452 12414 25508
rect 13122 25452 13132 25508
rect 13188 25452 13692 25508
rect 13748 25452 13758 25508
rect 14690 25452 14700 25508
rect 14756 25452 15484 25508
rect 15540 25452 15550 25508
rect 18610 25452 18620 25508
rect 18676 25452 20076 25508
rect 20132 25452 22540 25508
rect 22596 25452 22606 25508
rect 4610 25340 4620 25396
rect 4676 25340 5068 25396
rect 5124 25340 5852 25396
rect 5908 25340 5918 25396
rect 12338 25340 12348 25396
rect 12404 25340 12460 25396
rect 12516 25340 12526 25396
rect 12898 25340 12908 25396
rect 12964 25340 14028 25396
rect 14084 25340 14094 25396
rect 14914 25340 14924 25396
rect 14980 25340 15148 25396
rect 16146 25340 16156 25396
rect 16212 25340 18172 25396
rect 18228 25340 18732 25396
rect 18788 25340 19852 25396
rect 19908 25340 19918 25396
rect 23212 25340 25340 25396
rect 25396 25340 25406 25396
rect 25778 25340 25788 25396
rect 25844 25340 26908 25396
rect 26964 25340 27356 25396
rect 27412 25340 27422 25396
rect 15092 25284 15148 25340
rect 23212 25284 23268 25340
rect 12450 25228 12460 25284
rect 12516 25228 14252 25284
rect 14308 25228 14318 25284
rect 15092 25228 16268 25284
rect 16324 25228 16334 25284
rect 17826 25228 17836 25284
rect 17892 25228 18620 25284
rect 18676 25228 18686 25284
rect 19282 25228 19292 25284
rect 19348 25228 20300 25284
rect 20356 25228 23212 25284
rect 23268 25228 23278 25284
rect 25218 25228 25228 25284
rect 25284 25228 26684 25284
rect 26740 25228 26750 25284
rect 9518 25060 9528 25116
rect 9584 25060 9632 25116
rect 9688 25060 9736 25116
rect 9792 25060 9802 25116
rect 17834 25060 17844 25116
rect 17900 25060 17948 25116
rect 18004 25060 18052 25116
rect 18108 25060 18118 25116
rect 26150 25060 26160 25116
rect 26216 25060 26264 25116
rect 26320 25060 26368 25116
rect 26424 25060 26434 25116
rect 34466 25060 34476 25116
rect 34532 25060 34580 25116
rect 34636 25060 34684 25116
rect 34740 25060 34750 25116
rect 13346 25004 13356 25060
rect 13412 25004 14364 25060
rect 14420 25004 17500 25060
rect 17556 25004 17566 25060
rect 17500 24948 17556 25004
rect 3266 24892 3276 24948
rect 3332 24836 3388 24948
rect 5058 24892 5068 24948
rect 5124 24892 6076 24948
rect 6132 24892 6636 24948
rect 6692 24892 6702 24948
rect 9986 24892 9996 24948
rect 10052 24892 11116 24948
rect 11172 24892 11182 24948
rect 12114 24892 12124 24948
rect 12180 24892 12460 24948
rect 12516 24892 12526 24948
rect 14018 24892 14028 24948
rect 14084 24892 15260 24948
rect 15316 24892 16380 24948
rect 16436 24892 16446 24948
rect 17500 24892 18732 24948
rect 18788 24892 18798 24948
rect 22978 24892 22988 24948
rect 23044 24892 24332 24948
rect 24388 24892 24398 24948
rect 27458 24892 27468 24948
rect 27524 24892 28700 24948
rect 28756 24892 28766 24948
rect 3332 24780 4060 24836
rect 4116 24780 5740 24836
rect 5796 24780 5806 24836
rect 11778 24780 11788 24836
rect 11844 24780 12684 24836
rect 12740 24780 13132 24836
rect 13188 24780 13198 24836
rect 25890 24780 25900 24836
rect 25956 24780 29372 24836
rect 29428 24780 30044 24836
rect 30100 24780 30110 24836
rect 4610 24668 4620 24724
rect 4676 24668 5628 24724
rect 5684 24668 5694 24724
rect 12198 24668 12236 24724
rect 12292 24668 12302 24724
rect 12450 24668 12460 24724
rect 12516 24668 13244 24724
rect 13300 24668 13310 24724
rect 14550 24668 14588 24724
rect 14644 24668 14654 24724
rect 24658 24668 24668 24724
rect 24724 24668 25564 24724
rect 25620 24668 26012 24724
rect 26068 24668 26078 24724
rect 10322 24556 10332 24612
rect 10388 24556 11116 24612
rect 11172 24556 11182 24612
rect 19506 24556 19516 24612
rect 19572 24556 22428 24612
rect 22484 24556 22494 24612
rect 14466 24332 14476 24388
rect 14532 24332 14542 24388
rect 5360 24276 5370 24332
rect 5426 24276 5474 24332
rect 5530 24276 5578 24332
rect 5634 24276 5644 24332
rect 13676 24276 13686 24332
rect 13742 24276 13790 24332
rect 13846 24276 13894 24332
rect 13950 24276 13960 24332
rect 14476 24164 14532 24332
rect 21992 24276 22002 24332
rect 22058 24276 22106 24332
rect 22162 24276 22210 24332
rect 22266 24276 22276 24332
rect 30308 24276 30318 24332
rect 30374 24276 30422 24332
rect 30478 24276 30526 24332
rect 30582 24276 30592 24332
rect 4386 24108 4396 24164
rect 4452 24108 6300 24164
rect 6356 24108 6366 24164
rect 7746 24108 7756 24164
rect 7812 24108 8764 24164
rect 8820 24108 8830 24164
rect 9986 24108 9996 24164
rect 10052 24108 11564 24164
rect 11620 24108 14140 24164
rect 14196 24108 14206 24164
rect 14476 24108 15036 24164
rect 15092 24108 15102 24164
rect 8978 23996 8988 24052
rect 9044 23996 11004 24052
rect 11060 23996 11070 24052
rect 11890 23996 11900 24052
rect 11956 23996 13468 24052
rect 13524 23996 13534 24052
rect 14588 23996 20300 24052
rect 20356 23996 20366 24052
rect 25778 23996 25788 24052
rect 25844 23996 26460 24052
rect 26516 23996 27916 24052
rect 27972 23996 29372 24052
rect 29428 23996 29438 24052
rect 14588 23940 14644 23996
rect 10770 23884 10780 23940
rect 10836 23884 11228 23940
rect 11284 23884 11294 23940
rect 11778 23884 11788 23940
rect 11844 23884 12852 23940
rect 13010 23884 13020 23940
rect 13076 23884 13692 23940
rect 13748 23884 14588 23940
rect 14644 23884 14654 23940
rect 14924 23884 15596 23940
rect 15652 23884 15662 23940
rect 22754 23884 22764 23940
rect 22820 23884 23772 23940
rect 23828 23884 23838 23940
rect 25554 23884 25564 23940
rect 25620 23884 26684 23940
rect 26740 23884 28140 23940
rect 28196 23884 28206 23940
rect 11106 23772 11116 23828
rect 11172 23772 12012 23828
rect 12068 23772 12078 23828
rect 12226 23772 12236 23828
rect 12292 23772 12330 23828
rect 12534 23772 12572 23828
rect 12628 23772 12638 23828
rect 9518 23492 9528 23548
rect 9584 23492 9632 23548
rect 9688 23492 9736 23548
rect 9792 23492 9802 23548
rect 11116 23492 11172 23772
rect 12796 23716 12852 23884
rect 14924 23828 14980 23884
rect 13906 23772 13916 23828
rect 13972 23772 14924 23828
rect 14980 23772 14990 23828
rect 15922 23772 15932 23828
rect 15988 23772 17164 23828
rect 17220 23772 17230 23828
rect 18834 23772 18844 23828
rect 18900 23772 19516 23828
rect 19572 23772 19582 23828
rect 23426 23772 23436 23828
rect 23492 23772 24332 23828
rect 24388 23772 26124 23828
rect 26180 23772 26190 23828
rect 27122 23772 27132 23828
rect 27188 23772 29148 23828
rect 29204 23772 29214 23828
rect 12796 23660 13692 23716
rect 13748 23660 13758 23716
rect 14130 23660 14140 23716
rect 14196 23660 14476 23716
rect 14532 23660 14542 23716
rect 24770 23660 24780 23716
rect 24836 23660 25228 23716
rect 25284 23660 26796 23716
rect 26852 23660 27244 23716
rect 27300 23660 27310 23716
rect 27458 23660 27468 23716
rect 27524 23660 28364 23716
rect 28420 23660 29932 23716
rect 29988 23660 29998 23716
rect 11666 23548 11676 23604
rect 11732 23548 11900 23604
rect 11956 23548 11966 23604
rect 12338 23548 12348 23604
rect 12404 23548 12442 23604
rect 12562 23548 12572 23604
rect 12628 23548 12666 23604
rect 13458 23548 13468 23604
rect 13524 23548 15372 23604
rect 15428 23548 15438 23604
rect 17834 23492 17844 23548
rect 17900 23492 17948 23548
rect 18004 23492 18052 23548
rect 18108 23492 18118 23548
rect 26150 23492 26160 23548
rect 26216 23492 26264 23548
rect 26320 23492 26368 23548
rect 26424 23492 26434 23548
rect 34466 23492 34476 23548
rect 34532 23492 34580 23548
rect 34636 23492 34684 23548
rect 34740 23492 34750 23548
rect 11116 23436 11228 23492
rect 11284 23436 11294 23492
rect 12460 23436 14812 23492
rect 14868 23436 15820 23492
rect 15876 23436 15886 23492
rect 12460 23380 12516 23436
rect 9986 23324 9996 23380
rect 10052 23324 12124 23380
rect 12180 23324 12460 23380
rect 12516 23324 12526 23380
rect 12898 23324 12908 23380
rect 12964 23324 13916 23380
rect 13972 23324 14364 23380
rect 14420 23324 14430 23380
rect 16034 23324 16044 23380
rect 16100 23324 18620 23380
rect 18676 23324 18686 23380
rect 18946 23324 18956 23380
rect 19012 23324 19628 23380
rect 19684 23324 19694 23380
rect 22978 23324 22988 23380
rect 23044 23324 23884 23380
rect 23940 23324 23950 23380
rect 24658 23324 24668 23380
rect 24724 23324 25676 23380
rect 25732 23324 25742 23380
rect 4946 23212 4956 23268
rect 5012 23212 5852 23268
rect 5908 23212 5918 23268
rect 9874 23212 9884 23268
rect 9940 23212 11452 23268
rect 11508 23212 12684 23268
rect 12740 23212 12750 23268
rect 15362 23212 15372 23268
rect 15428 23212 17612 23268
rect 17668 23212 19068 23268
rect 19124 23212 19134 23268
rect 20402 23212 20412 23268
rect 20468 23212 20972 23268
rect 21028 23212 25452 23268
rect 25508 23212 27020 23268
rect 27076 23212 27086 23268
rect 12114 23100 12124 23156
rect 12180 23100 13020 23156
rect 13076 23100 13086 23156
rect 14354 23100 14364 23156
rect 14420 23100 15036 23156
rect 15092 23100 15102 23156
rect 15586 23100 15596 23156
rect 15652 23100 17724 23156
rect 17780 23100 19348 23156
rect 24434 23100 24444 23156
rect 24500 23100 26124 23156
rect 26180 23100 26190 23156
rect 19292 23044 19348 23100
rect 8866 22988 8876 23044
rect 8932 22988 12572 23044
rect 12628 22988 12638 23044
rect 17938 22988 17948 23044
rect 18004 22988 18396 23044
rect 18452 22988 18462 23044
rect 19282 22988 19292 23044
rect 19348 22988 19358 23044
rect 2706 22876 2716 22932
rect 2772 22876 6412 22932
rect 6468 22876 6478 22932
rect 10882 22876 10892 22932
rect 10948 22876 19628 22932
rect 19684 22876 19694 22932
rect 11218 22764 11228 22820
rect 11284 22764 11340 22820
rect 11396 22764 11406 22820
rect 5360 22708 5370 22764
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5634 22708 5644 22764
rect 13676 22708 13686 22764
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13950 22708 13960 22764
rect 21992 22708 22002 22764
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22266 22708 22276 22764
rect 30308 22708 30318 22764
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30582 22708 30592 22764
rect 2482 22540 2492 22596
rect 2548 22540 5628 22596
rect 5684 22540 5694 22596
rect 6290 22540 6300 22596
rect 6356 22540 17388 22596
rect 17444 22540 17454 22596
rect 26114 22540 26124 22596
rect 26180 22540 26908 22596
rect 26964 22540 26974 22596
rect 7074 22428 7084 22484
rect 7140 22428 7868 22484
rect 7924 22428 7934 22484
rect 10882 22428 10892 22484
rect 10948 22428 11340 22484
rect 11396 22428 11406 22484
rect 25778 22428 25788 22484
rect 25844 22428 27132 22484
rect 27188 22428 27198 22484
rect 3602 22316 3612 22372
rect 3668 22316 6076 22372
rect 6132 22316 6142 22372
rect 12898 22316 12908 22372
rect 12964 22316 17500 22372
rect 17556 22316 19852 22372
rect 19908 22316 19918 22372
rect 20066 22316 20076 22372
rect 20132 22316 21420 22372
rect 21476 22316 21486 22372
rect 8418 22204 8428 22260
rect 8484 22204 13580 22260
rect 13636 22204 13646 22260
rect 19618 22204 19628 22260
rect 19684 22204 20188 22260
rect 20244 22204 20254 22260
rect 20626 22204 20636 22260
rect 20692 22204 22204 22260
rect 22260 22204 22270 22260
rect 25666 22092 25676 22148
rect 25732 22092 26124 22148
rect 26180 22092 27244 22148
rect 27300 22092 27310 22148
rect 11554 21980 11564 22036
rect 11620 21980 13580 22036
rect 13636 21980 13646 22036
rect 9518 21924 9528 21980
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9792 21924 9802 21980
rect 17834 21924 17844 21980
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 18108 21924 18118 21980
rect 26150 21924 26160 21980
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26424 21924 26434 21980
rect 34466 21924 34476 21980
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34740 21924 34750 21980
rect 12338 21868 12348 21924
rect 12404 21868 12414 21924
rect 12348 21812 12404 21868
rect 4834 21756 4844 21812
rect 4900 21756 5516 21812
rect 5572 21756 5582 21812
rect 10994 21756 11004 21812
rect 11060 21756 12404 21812
rect 12674 21756 12684 21812
rect 12740 21756 13356 21812
rect 13412 21756 13422 21812
rect 14466 21756 14476 21812
rect 14532 21756 15708 21812
rect 15764 21756 16380 21812
rect 16436 21756 16446 21812
rect 16706 21756 16716 21812
rect 16772 21756 18956 21812
rect 19012 21756 19022 21812
rect 19394 21756 19404 21812
rect 19460 21756 19628 21812
rect 19684 21756 20580 21812
rect 21970 21756 21980 21812
rect 22036 21756 22652 21812
rect 22708 21756 24444 21812
rect 24500 21756 24510 21812
rect 25442 21756 25452 21812
rect 25508 21756 26684 21812
rect 26740 21756 27020 21812
rect 27076 21756 27086 21812
rect 20524 21700 20580 21756
rect 3938 21644 3948 21700
rect 4004 21644 4620 21700
rect 4676 21644 5404 21700
rect 5460 21644 5470 21700
rect 12338 21644 12348 21700
rect 12404 21644 13244 21700
rect 13300 21644 13310 21700
rect 13458 21644 13468 21700
rect 13524 21644 14812 21700
rect 14868 21644 14878 21700
rect 18274 21644 18284 21700
rect 18340 21644 19292 21700
rect 19348 21644 19358 21700
rect 20514 21644 20524 21700
rect 20580 21644 21644 21700
rect 21700 21644 23548 21700
rect 23604 21644 23614 21700
rect 10322 21532 10332 21588
rect 10388 21532 10892 21588
rect 10948 21532 10958 21588
rect 14690 21532 14700 21588
rect 14756 21532 15932 21588
rect 15988 21532 15998 21588
rect 23874 21532 23884 21588
rect 23940 21532 26124 21588
rect 26180 21532 27244 21588
rect 27300 21532 27310 21588
rect 10658 21420 10668 21476
rect 10724 21420 12012 21476
rect 12068 21420 12078 21476
rect 13010 21420 13020 21476
rect 13076 21420 15372 21476
rect 15428 21420 15438 21476
rect 21746 21420 21756 21476
rect 21812 21420 24556 21476
rect 24612 21420 24622 21476
rect 27458 21420 27468 21476
rect 27524 21420 28812 21476
rect 28868 21420 28878 21476
rect 25442 21308 25452 21364
rect 25508 21308 27020 21364
rect 27076 21308 27086 21364
rect 10658 21196 10668 21252
rect 10724 21196 12348 21252
rect 12404 21196 12414 21252
rect 25890 21196 25900 21252
rect 25956 21196 27580 21252
rect 27636 21196 27646 21252
rect 5360 21140 5370 21196
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5634 21140 5644 21196
rect 13676 21140 13686 21196
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13950 21140 13960 21196
rect 21992 21140 22002 21196
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22266 21140 22276 21196
rect 30308 21140 30318 21196
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30582 21140 30592 21196
rect 12786 20972 12796 21028
rect 12852 20972 15484 21028
rect 15540 20972 15550 21028
rect 20402 20972 20412 21028
rect 20468 20972 22540 21028
rect 22596 20972 22606 21028
rect 16706 20860 16716 20916
rect 16772 20860 17388 20916
rect 17444 20860 17454 20916
rect 24434 20860 24444 20916
rect 24500 20860 26012 20916
rect 26068 20860 26078 20916
rect 3266 20748 3276 20804
rect 3332 20748 4284 20804
rect 4340 20748 4732 20804
rect 4788 20748 7644 20804
rect 7700 20748 7710 20804
rect 13570 20748 13580 20804
rect 13636 20748 14140 20804
rect 14196 20748 14206 20804
rect 14354 20748 14364 20804
rect 14420 20748 16044 20804
rect 16100 20748 16110 20804
rect 21522 20748 21532 20804
rect 21588 20748 22876 20804
rect 22932 20748 22942 20804
rect 3938 20636 3948 20692
rect 4004 20636 4620 20692
rect 4676 20636 8204 20692
rect 8260 20636 8270 20692
rect 17154 20636 17164 20692
rect 17220 20636 17612 20692
rect 17668 20636 21196 20692
rect 21252 20636 21262 20692
rect 2370 20524 2380 20580
rect 2436 20524 2940 20580
rect 2996 20524 3388 20580
rect 3444 20524 4284 20580
rect 4340 20524 4844 20580
rect 4900 20524 4910 20580
rect 9874 20524 9884 20580
rect 9940 20524 10444 20580
rect 10500 20524 10780 20580
rect 10836 20524 10846 20580
rect 11442 20524 11452 20580
rect 11508 20524 12796 20580
rect 12852 20524 14364 20580
rect 14420 20524 14430 20580
rect 17714 20524 17724 20580
rect 17780 20524 18396 20580
rect 18452 20524 18462 20580
rect 9518 20356 9528 20412
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9792 20356 9802 20412
rect 17834 20356 17844 20412
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 18108 20356 18118 20412
rect 26150 20356 26160 20412
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26424 20356 26434 20412
rect 34466 20356 34476 20412
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34740 20356 34750 20412
rect 4946 20188 4956 20244
rect 5012 20188 9996 20244
rect 10052 20188 10062 20244
rect 11330 20188 11340 20244
rect 11396 20188 12124 20244
rect 12180 20188 12190 20244
rect 4386 20076 4396 20132
rect 4452 20076 5404 20132
rect 5460 20076 5470 20132
rect 8194 20076 8204 20132
rect 8260 20076 10220 20132
rect 10276 20076 12460 20132
rect 12516 20076 12526 20132
rect 13122 20076 13132 20132
rect 13188 20076 13580 20132
rect 13636 20076 14028 20132
rect 14084 20076 14094 20132
rect 15092 20076 15372 20132
rect 15428 20076 16604 20132
rect 16660 20076 17948 20132
rect 18004 20076 18014 20132
rect 22194 20076 22204 20132
rect 22260 20076 23436 20132
rect 23492 20076 24444 20132
rect 24500 20076 24510 20132
rect 29698 20076 29708 20132
rect 29764 20076 30604 20132
rect 30660 20076 30670 20132
rect 15092 20020 15148 20076
rect 3602 19964 3612 20020
rect 3668 19964 4508 20020
rect 4564 19964 5180 20020
rect 5236 19964 5246 20020
rect 7298 19964 7308 20020
rect 7364 19964 8876 20020
rect 8932 19964 9436 20020
rect 9492 19964 9502 20020
rect 9986 19964 9996 20020
rect 10052 19964 14252 20020
rect 14308 19964 15148 20020
rect 15698 19964 15708 20020
rect 15764 19964 17276 20020
rect 17332 19964 17342 20020
rect 18162 19964 18172 20020
rect 18228 19964 18620 20020
rect 18676 19964 18686 20020
rect 19618 19964 19628 20020
rect 19684 19964 20636 20020
rect 20692 19964 20702 20020
rect 21074 19964 21084 20020
rect 21140 19964 22988 20020
rect 23044 19964 23054 20020
rect 24658 19964 24668 20020
rect 24724 19964 25228 20020
rect 25284 19964 25294 20020
rect 27122 19964 27132 20020
rect 27188 19964 29148 20020
rect 29204 19964 29214 20020
rect 2482 19852 2492 19908
rect 2548 19852 5068 19908
rect 5124 19852 5134 19908
rect 7970 19852 7980 19908
rect 8036 19852 9660 19908
rect 9716 19852 9726 19908
rect 10322 19852 10332 19908
rect 10388 19852 14588 19908
rect 14644 19852 14654 19908
rect 14802 19852 14812 19908
rect 14868 19852 16156 19908
rect 16212 19852 16222 19908
rect 16370 19852 16380 19908
rect 16436 19852 18284 19908
rect 18340 19852 19180 19908
rect 19236 19852 19246 19908
rect 21522 19852 21532 19908
rect 21588 19852 21868 19908
rect 21924 19852 21934 19908
rect 10994 19740 11004 19796
rect 11060 19740 12572 19796
rect 12628 19740 12638 19796
rect 18050 19740 18060 19796
rect 18116 19740 18956 19796
rect 19012 19740 19022 19796
rect 19180 19740 26684 19796
rect 26740 19740 26750 19796
rect 19180 19684 19236 19740
rect 16818 19628 16828 19684
rect 16884 19628 19236 19684
rect 5360 19572 5370 19628
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5634 19572 5644 19628
rect 13676 19572 13686 19628
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13950 19572 13960 19628
rect 21992 19572 22002 19628
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22266 19572 22276 19628
rect 30308 19572 30318 19628
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30582 19572 30592 19628
rect 8978 19292 8988 19348
rect 9044 19292 10556 19348
rect 10612 19292 10622 19348
rect 12338 19292 12348 19348
rect 12404 19292 13356 19348
rect 13412 19292 13422 19348
rect 17378 19292 17388 19348
rect 17444 19292 18396 19348
rect 18452 19292 20524 19348
rect 20580 19292 20590 19348
rect 26450 19292 26460 19348
rect 26516 19292 27132 19348
rect 27188 19292 27198 19348
rect 9762 19180 9772 19236
rect 9828 19180 10332 19236
rect 10388 19180 10398 19236
rect 9090 19068 9100 19124
rect 9156 19068 10556 19124
rect 10612 19068 10622 19124
rect 14578 19068 14588 19124
rect 14644 19068 15036 19124
rect 15092 19068 17276 19124
rect 17332 19068 22876 19124
rect 22932 19068 22942 19124
rect 8204 18956 9996 19012
rect 10052 18956 10062 19012
rect 10882 18956 10892 19012
rect 10948 18956 11900 19012
rect 11956 18956 11966 19012
rect 16930 18956 16940 19012
rect 16996 18956 17388 19012
rect 17444 18956 17454 19012
rect 28018 18956 28028 19012
rect 28084 18956 29372 19012
rect 29428 18956 29438 19012
rect 8204 18788 8260 18956
rect 10322 18844 10332 18900
rect 10388 18844 10780 18900
rect 10836 18844 10846 18900
rect 9518 18788 9528 18844
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9792 18788 9802 18844
rect 17834 18788 17844 18844
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 18108 18788 18118 18844
rect 26150 18788 26160 18844
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26424 18788 26434 18844
rect 34466 18788 34476 18844
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34740 18788 34750 18844
rect 6962 18732 6972 18788
rect 7028 18732 8204 18788
rect 8260 18732 8270 18788
rect 11078 18732 11116 18788
rect 11172 18732 11182 18788
rect 7410 18620 7420 18676
rect 7476 18620 11228 18676
rect 11284 18620 11294 18676
rect 18946 18620 18956 18676
rect 19012 18620 21644 18676
rect 21700 18620 21710 18676
rect 6738 18508 6748 18564
rect 6804 18508 7756 18564
rect 7812 18508 7822 18564
rect 7970 18508 7980 18564
rect 8036 18508 8876 18564
rect 8932 18508 8942 18564
rect 9100 18508 9660 18564
rect 9716 18508 9726 18564
rect 16818 18508 16828 18564
rect 16884 18508 17500 18564
rect 17556 18508 17566 18564
rect 30706 18508 30716 18564
rect 30772 18508 30782 18564
rect 7756 18452 7812 18508
rect 9100 18452 9156 18508
rect 30716 18452 30772 18508
rect 7756 18396 9156 18452
rect 10546 18396 10556 18452
rect 10612 18396 11788 18452
rect 11844 18396 11854 18452
rect 14018 18396 14028 18452
rect 14084 18396 15596 18452
rect 15652 18396 18508 18452
rect 18564 18396 18574 18452
rect 22866 18396 22876 18452
rect 22932 18396 23548 18452
rect 23604 18396 23614 18452
rect 25666 18396 25676 18452
rect 25732 18396 30772 18452
rect 9874 18284 9884 18340
rect 9940 18284 12348 18340
rect 12404 18284 12414 18340
rect 14690 18284 14700 18340
rect 14756 18284 16044 18340
rect 16100 18284 16110 18340
rect 16482 18284 16492 18340
rect 16548 18284 17500 18340
rect 17556 18284 17566 18340
rect 22530 18284 22540 18340
rect 22596 18284 25452 18340
rect 25508 18284 25518 18340
rect 25452 18228 25508 18284
rect 8866 18172 8876 18228
rect 8932 18172 10108 18228
rect 10164 18172 10174 18228
rect 10434 18172 10444 18228
rect 10500 18172 11116 18228
rect 11172 18172 11182 18228
rect 17938 18172 17948 18228
rect 18004 18172 23212 18228
rect 23268 18172 23278 18228
rect 25452 18172 26684 18228
rect 26740 18172 26750 18228
rect 8194 18060 8204 18116
rect 8260 18060 12796 18116
rect 12852 18060 12862 18116
rect 5360 18004 5370 18060
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5634 18004 5644 18060
rect 13676 18004 13686 18060
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13950 18004 13960 18060
rect 21992 18004 22002 18060
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22266 18004 22276 18060
rect 30308 18004 30318 18060
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30582 18004 30592 18060
rect 6850 17836 6860 17892
rect 6916 17836 7196 17892
rect 7252 17836 7262 17892
rect 8418 17836 8428 17892
rect 8484 17836 9548 17892
rect 9604 17836 9614 17892
rect 10994 17724 11004 17780
rect 11060 17724 11116 17780
rect 11172 17724 11182 17780
rect 17014 17724 17052 17780
rect 17108 17724 17118 17780
rect 21298 17724 21308 17780
rect 21364 17724 21756 17780
rect 21812 17724 23548 17780
rect 23604 17724 24556 17780
rect 24612 17724 24622 17780
rect 27458 17724 27468 17780
rect 27524 17724 29036 17780
rect 29092 17724 29102 17780
rect 31938 17724 31948 17780
rect 32004 17724 33292 17780
rect 33348 17724 33358 17780
rect 4610 17612 4620 17668
rect 4676 17612 5740 17668
rect 5796 17612 6524 17668
rect 6580 17612 6590 17668
rect 7084 17612 7644 17668
rect 7700 17612 8316 17668
rect 8372 17612 8382 17668
rect 8530 17612 8540 17668
rect 8596 17612 10220 17668
rect 10276 17612 10286 17668
rect 28914 17612 28924 17668
rect 28980 17612 29372 17668
rect 29428 17612 29438 17668
rect 7084 17556 7140 17612
rect 5954 17500 5964 17556
rect 6020 17500 7084 17556
rect 7140 17500 7150 17556
rect 9090 17500 9100 17556
rect 9156 17500 10668 17556
rect 10724 17500 10734 17556
rect 14354 17500 14364 17556
rect 14420 17500 16156 17556
rect 16212 17500 17388 17556
rect 17444 17500 18172 17556
rect 18228 17500 18238 17556
rect 9762 17388 9772 17444
rect 9828 17388 11116 17444
rect 11172 17388 11182 17444
rect 17826 17388 17836 17444
rect 17892 17388 18508 17444
rect 18564 17388 18574 17444
rect 19058 17388 19068 17444
rect 19124 17388 20636 17444
rect 20692 17388 20702 17444
rect 8082 17276 8092 17332
rect 8148 17276 8428 17332
rect 8484 17276 8494 17332
rect 9518 17220 9528 17276
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9792 17220 9802 17276
rect 17834 17220 17844 17276
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 18108 17220 18118 17276
rect 26150 17220 26160 17276
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26424 17220 26434 17276
rect 34466 17220 34476 17276
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34740 17220 34750 17276
rect 18498 17164 18508 17220
rect 18564 17164 19628 17220
rect 19684 17164 19694 17220
rect 7746 17052 7756 17108
rect 7812 17052 8204 17108
rect 8260 17052 8270 17108
rect 9874 17052 9884 17108
rect 9940 17052 10556 17108
rect 10612 17052 11228 17108
rect 11284 17052 11294 17108
rect 15250 17052 15260 17108
rect 15316 17052 17276 17108
rect 17332 17052 17342 17108
rect 18162 17052 18172 17108
rect 18228 17052 18956 17108
rect 19012 17052 19022 17108
rect 5058 16940 5068 16996
rect 5124 16940 6748 16996
rect 6804 16940 7196 16996
rect 7252 16940 7262 16996
rect 7970 16940 7980 16996
rect 8036 16940 10444 16996
rect 10500 16940 10510 16996
rect 15922 16940 15932 16996
rect 15988 16940 16716 16996
rect 16772 16940 17836 16996
rect 17892 16940 17902 16996
rect 28018 16940 28028 16996
rect 28084 16940 29372 16996
rect 29428 16940 29438 16996
rect 15932 16884 15988 16940
rect 3938 16828 3948 16884
rect 4004 16828 5852 16884
rect 5908 16828 5918 16884
rect 6290 16828 6300 16884
rect 6356 16828 7532 16884
rect 7588 16828 7598 16884
rect 10770 16828 10780 16884
rect 10836 16828 12236 16884
rect 12292 16828 12302 16884
rect 12898 16828 12908 16884
rect 12964 16828 14140 16884
rect 14196 16828 15988 16884
rect 17042 16828 17052 16884
rect 17108 16828 17948 16884
rect 18004 16828 18014 16884
rect 27570 16828 27580 16884
rect 27636 16828 29484 16884
rect 29540 16828 29550 16884
rect 8306 16716 8316 16772
rect 8372 16716 11676 16772
rect 11732 16716 11742 16772
rect 12338 16716 12348 16772
rect 12404 16716 14028 16772
rect 14084 16716 14094 16772
rect 14914 16716 14924 16772
rect 14980 16716 15596 16772
rect 15652 16716 15662 16772
rect 17602 16716 17612 16772
rect 17668 16716 18508 16772
rect 18564 16716 18574 16772
rect 20066 16716 20076 16772
rect 20132 16716 22540 16772
rect 22596 16716 22606 16772
rect 26114 16716 26124 16772
rect 26180 16716 28140 16772
rect 28196 16716 28206 16772
rect 29810 16716 29820 16772
rect 29876 16716 30380 16772
rect 30436 16716 31500 16772
rect 31556 16716 31566 16772
rect 13906 16604 13916 16660
rect 13972 16604 15260 16660
rect 15316 16604 15326 16660
rect 16706 16604 16716 16660
rect 16772 16604 19292 16660
rect 19348 16604 19358 16660
rect 21858 16604 21868 16660
rect 21924 16604 22876 16660
rect 22932 16604 23436 16660
rect 23492 16604 24556 16660
rect 24612 16604 24622 16660
rect 5360 16436 5370 16492
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5634 16436 5644 16492
rect 13676 16436 13686 16492
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13950 16436 13960 16492
rect 21992 16436 22002 16492
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22266 16436 22276 16492
rect 30308 16436 30318 16492
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30582 16436 30592 16492
rect 16930 16268 16940 16324
rect 16996 16268 17948 16324
rect 18004 16268 18014 16324
rect 25778 16268 25788 16324
rect 25844 16268 27468 16324
rect 27524 16268 27534 16324
rect 12786 16156 12796 16212
rect 12852 16156 13692 16212
rect 13748 16156 13758 16212
rect 21634 16156 21644 16212
rect 21700 16156 23436 16212
rect 23492 16156 23502 16212
rect 14914 16044 14924 16100
rect 14980 16044 15484 16100
rect 15540 16044 15550 16100
rect 16146 16044 16156 16100
rect 16212 16044 16716 16100
rect 16772 16044 17612 16100
rect 17668 16044 17678 16100
rect 21746 16044 21756 16100
rect 21812 16044 22428 16100
rect 22484 16044 23660 16100
rect 23716 16044 23726 16100
rect 26226 16044 26236 16100
rect 26292 16044 29372 16100
rect 29428 16044 29438 16100
rect 14130 15932 14140 15988
rect 14196 15932 14812 15988
rect 14868 15932 14878 15988
rect 15250 15932 15260 15988
rect 15316 15932 16044 15988
rect 16100 15932 16110 15988
rect 16930 15932 16940 15988
rect 16996 15932 18732 15988
rect 18788 15932 18798 15988
rect 20962 15932 20972 15988
rect 21028 15932 21532 15988
rect 21588 15932 21598 15988
rect 22642 15932 22652 15988
rect 22708 15932 24332 15988
rect 24388 15932 24398 15988
rect 26114 15932 26124 15988
rect 26180 15932 27916 15988
rect 27972 15932 27982 15988
rect 28242 15932 28252 15988
rect 28308 15932 28924 15988
rect 28980 15932 28990 15988
rect 18274 15820 18284 15876
rect 18340 15820 19068 15876
rect 19124 15820 19134 15876
rect 26002 15820 26012 15876
rect 26068 15820 27468 15876
rect 27524 15820 28028 15876
rect 28084 15820 28094 15876
rect 15138 15708 15148 15764
rect 15204 15708 15708 15764
rect 15764 15708 16828 15764
rect 16884 15708 16894 15764
rect 31154 15708 31164 15764
rect 31220 15708 32284 15764
rect 32340 15708 32350 15764
rect 9518 15652 9528 15708
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9792 15652 9802 15708
rect 17834 15652 17844 15708
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 18108 15652 18118 15708
rect 26150 15652 26160 15708
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26424 15652 26434 15708
rect 34466 15652 34476 15708
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34740 15652 34750 15708
rect 15474 15484 15484 15540
rect 15540 15484 18956 15540
rect 19012 15484 19022 15540
rect 30370 15484 30380 15540
rect 30436 15484 31444 15540
rect 31388 15428 31444 15484
rect 14018 15372 14028 15428
rect 14084 15372 15260 15428
rect 15316 15372 16436 15428
rect 16818 15372 16828 15428
rect 16884 15372 19068 15428
rect 19124 15372 19134 15428
rect 28130 15372 28140 15428
rect 28196 15372 30940 15428
rect 30996 15372 31006 15428
rect 31378 15372 31388 15428
rect 31444 15372 33628 15428
rect 33684 15372 33694 15428
rect 16380 15316 16436 15372
rect 11218 15260 11228 15316
rect 11284 15260 13468 15316
rect 13524 15260 13534 15316
rect 14802 15260 14812 15316
rect 14868 15260 15708 15316
rect 15764 15260 15774 15316
rect 16380 15260 18732 15316
rect 18788 15260 18798 15316
rect 23986 15260 23996 15316
rect 24052 15260 28028 15316
rect 28084 15260 28094 15316
rect 28802 15260 28812 15316
rect 28868 15260 31500 15316
rect 31556 15260 31566 15316
rect 1586 15148 1596 15204
rect 1652 15148 17948 15204
rect 18004 15148 18014 15204
rect 27346 15148 27356 15204
rect 27412 15148 28252 15204
rect 28308 15148 28318 15204
rect 30594 15148 30604 15204
rect 30660 15148 32508 15204
rect 32564 15148 33180 15204
rect 33236 15148 33246 15204
rect 1810 15036 1820 15092
rect 1876 15036 2268 15092
rect 2324 15036 3276 15092
rect 3332 15036 5068 15092
rect 5124 15036 5740 15092
rect 5796 15036 6300 15092
rect 6356 15036 6366 15092
rect 8978 15036 8988 15092
rect 9044 15036 9996 15092
rect 10052 15036 10062 15092
rect 16370 15036 16380 15092
rect 16436 15036 16940 15092
rect 16996 15036 17006 15092
rect 30482 15036 30492 15092
rect 30548 15036 32788 15092
rect 32732 14980 32788 15036
rect 16482 14924 16492 14980
rect 16548 14924 16716 14980
rect 16772 14924 16782 14980
rect 32722 14924 32732 14980
rect 32788 14924 32798 14980
rect 5360 14868 5370 14924
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5634 14868 5644 14924
rect 13676 14868 13686 14924
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13950 14868 13960 14924
rect 21992 14868 22002 14924
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22266 14868 22276 14924
rect 30308 14868 30318 14924
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30582 14868 30592 14924
rect 27906 14700 27916 14756
rect 27972 14700 28476 14756
rect 28532 14700 32172 14756
rect 32228 14700 32238 14756
rect 21634 14588 21644 14644
rect 21700 14588 23436 14644
rect 23492 14588 23502 14644
rect 16930 14476 16940 14532
rect 16996 14476 17276 14532
rect 17332 14476 17342 14532
rect 27234 14476 27244 14532
rect 27300 14476 27916 14532
rect 27972 14476 28700 14532
rect 28756 14476 28766 14532
rect 32050 14476 32060 14532
rect 32116 14476 33068 14532
rect 33124 14476 33134 14532
rect 12674 14364 12684 14420
rect 12740 14364 13580 14420
rect 13636 14364 19180 14420
rect 19236 14364 19964 14420
rect 20020 14364 20030 14420
rect 25442 14364 25452 14420
rect 25508 14364 29148 14420
rect 29204 14364 30044 14420
rect 30100 14364 30110 14420
rect 2930 14252 2940 14308
rect 2996 14252 3724 14308
rect 3780 14252 3790 14308
rect 4610 14252 4620 14308
rect 4676 14252 5628 14308
rect 5684 14252 5694 14308
rect 17378 14252 17388 14308
rect 17444 14252 18844 14308
rect 18900 14252 18910 14308
rect 20514 14252 20524 14308
rect 20580 14252 21420 14308
rect 21476 14252 21486 14308
rect 9518 14084 9528 14140
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9792 14084 9802 14140
rect 17834 14084 17844 14140
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 18108 14084 18118 14140
rect 26150 14084 26160 14140
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26424 14084 26434 14140
rect 34466 14084 34476 14140
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34740 14084 34750 14140
rect 5954 14028 5964 14084
rect 6020 14028 8540 14084
rect 8596 14028 8606 14084
rect 19842 14028 19852 14084
rect 19908 14028 21196 14084
rect 21252 14028 21262 14084
rect 8540 13972 8596 14028
rect 8540 13916 9772 13972
rect 9828 13916 9838 13972
rect 11666 13916 11676 13972
rect 11732 13916 14140 13972
rect 14196 13916 16268 13972
rect 16324 13916 16334 13972
rect 18386 13916 18396 13972
rect 18452 13916 19516 13972
rect 19572 13916 19582 13972
rect 20066 13916 20076 13972
rect 20132 13916 22204 13972
rect 22260 13916 22270 13972
rect 5954 13804 5964 13860
rect 6020 13804 7308 13860
rect 7364 13804 7374 13860
rect 7634 13804 7644 13860
rect 7700 13804 9940 13860
rect 10098 13804 10108 13860
rect 10164 13804 11116 13860
rect 11172 13804 11182 13860
rect 17714 13804 17724 13860
rect 17780 13804 19628 13860
rect 19684 13804 20300 13860
rect 20356 13804 20366 13860
rect 25666 13804 25676 13860
rect 25732 13804 26796 13860
rect 26852 13804 27020 13860
rect 27076 13804 27086 13860
rect 9884 13748 9940 13804
rect 5506 13692 5516 13748
rect 5572 13692 9548 13748
rect 9604 13692 9614 13748
rect 9884 13692 10892 13748
rect 10948 13692 13132 13748
rect 13188 13692 13198 13748
rect 18722 13692 18732 13748
rect 18788 13692 19740 13748
rect 19796 13692 20188 13748
rect 20244 13692 20254 13748
rect 23874 13692 23884 13748
rect 23940 13692 25452 13748
rect 25508 13692 25518 13748
rect 26114 13692 26124 13748
rect 26180 13692 27468 13748
rect 27524 13692 27534 13748
rect 9986 13580 9996 13636
rect 10052 13580 10780 13636
rect 10836 13580 11900 13636
rect 11956 13580 11966 13636
rect 26450 13580 26460 13636
rect 26516 13580 27244 13636
rect 27300 13580 27310 13636
rect 28018 13580 28028 13636
rect 28084 13580 32396 13636
rect 32452 13580 32462 13636
rect 33058 13580 33068 13636
rect 33124 13580 33572 13636
rect 33516 13524 33572 13580
rect 5058 13468 5068 13524
rect 5124 13468 6748 13524
rect 6804 13468 8428 13524
rect 8484 13468 8494 13524
rect 9538 13468 9548 13524
rect 9604 13468 12852 13524
rect 16594 13468 16604 13524
rect 16660 13468 18956 13524
rect 19012 13468 19022 13524
rect 19506 13468 19516 13524
rect 19572 13468 21308 13524
rect 21364 13468 21374 13524
rect 21634 13468 21644 13524
rect 21700 13468 21980 13524
rect 22036 13468 22988 13524
rect 23044 13468 23054 13524
rect 24770 13468 24780 13524
rect 24836 13468 26908 13524
rect 26964 13468 26974 13524
rect 31266 13468 31276 13524
rect 31332 13468 33292 13524
rect 33348 13468 33358 13524
rect 33506 13468 33516 13524
rect 33572 13468 33582 13524
rect 7868 13412 7924 13468
rect 8428 13412 8484 13468
rect 7858 13356 7868 13412
rect 7924 13356 7934 13412
rect 8428 13356 12572 13412
rect 12628 13356 12638 13412
rect 5360 13300 5370 13356
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5634 13300 5644 13356
rect 12796 13188 12852 13468
rect 26338 13356 26348 13412
rect 26404 13356 27580 13412
rect 27636 13356 27646 13412
rect 13676 13300 13686 13356
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13950 13300 13960 13356
rect 21992 13300 22002 13356
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22266 13300 22276 13356
rect 30308 13300 30318 13356
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30582 13300 30592 13356
rect 12796 13132 15820 13188
rect 15876 13132 15886 13188
rect 20290 13132 20300 13188
rect 20356 13132 22092 13188
rect 22148 13132 22652 13188
rect 22708 13132 22718 13188
rect 29586 13132 29596 13188
rect 29652 13132 31836 13188
rect 31892 13132 31902 13188
rect 9762 13020 9772 13076
rect 9828 13020 12124 13076
rect 12180 13020 12190 13076
rect 20066 13020 20076 13076
rect 20132 13020 20748 13076
rect 20804 13020 20814 13076
rect 21746 13020 21756 13076
rect 21812 13020 22428 13076
rect 22484 13020 22494 13076
rect 22754 13020 22764 13076
rect 22820 13020 22830 13076
rect 22764 12964 22820 13020
rect 4946 12908 4956 12964
rect 5012 12908 5852 12964
rect 5908 12908 6188 12964
rect 6244 12908 6254 12964
rect 16034 12908 16044 12964
rect 16100 12908 16828 12964
rect 16884 12908 18396 12964
rect 18452 12908 18462 12964
rect 20514 12908 20524 12964
rect 20580 12908 21868 12964
rect 21924 12908 21934 12964
rect 22306 12908 22316 12964
rect 22372 12908 22820 12964
rect 26852 12908 28028 12964
rect 28084 12908 29372 12964
rect 29428 12908 29438 12964
rect 7522 12796 7532 12852
rect 7588 12796 10108 12852
rect 10164 12796 10174 12852
rect 15698 12796 15708 12852
rect 15764 12796 17388 12852
rect 17444 12796 17454 12852
rect 20972 12740 21028 12908
rect 26852 12852 26908 12908
rect 21634 12796 21644 12852
rect 21700 12796 22876 12852
rect 22932 12796 22942 12852
rect 26674 12796 26684 12852
rect 26740 12796 26908 12852
rect 3602 12684 3612 12740
rect 3668 12684 5404 12740
rect 5460 12684 5470 12740
rect 11330 12684 11340 12740
rect 11396 12684 12012 12740
rect 12068 12684 12078 12740
rect 13122 12684 13132 12740
rect 13188 12684 13804 12740
rect 13860 12684 13870 12740
rect 16258 12684 16268 12740
rect 16324 12684 16940 12740
rect 16996 12684 17006 12740
rect 18162 12684 18172 12740
rect 18228 12684 19740 12740
rect 19796 12684 19806 12740
rect 20962 12684 20972 12740
rect 21028 12684 21038 12740
rect 2818 12572 2828 12628
rect 2884 12572 7196 12628
rect 7252 12572 8316 12628
rect 8372 12572 8652 12628
rect 8708 12572 8718 12628
rect 20738 12572 20748 12628
rect 20804 12572 22316 12628
rect 22372 12572 22382 12628
rect 9518 12516 9528 12572
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9792 12516 9802 12572
rect 17834 12516 17844 12572
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 18108 12516 18118 12572
rect 26150 12516 26160 12572
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26424 12516 26434 12572
rect 34466 12516 34476 12572
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34740 12516 34750 12572
rect 4610 12460 4620 12516
rect 4676 12460 5516 12516
rect 5572 12460 5582 12516
rect 5058 12348 5068 12404
rect 5124 12348 6524 12404
rect 6580 12348 7308 12404
rect 7364 12348 7374 12404
rect 18498 12348 18508 12404
rect 18564 12348 19964 12404
rect 20020 12348 20636 12404
rect 20692 12348 20702 12404
rect 5842 12236 5852 12292
rect 5908 12236 6412 12292
rect 6468 12236 8988 12292
rect 9044 12236 10668 12292
rect 10724 12236 10734 12292
rect 17602 12236 17612 12292
rect 17668 12236 18284 12292
rect 18340 12236 19404 12292
rect 19460 12236 19470 12292
rect 3826 12124 3836 12180
rect 3892 12124 4508 12180
rect 4564 12124 6076 12180
rect 6132 12124 6142 12180
rect 4956 12012 8204 12068
rect 8260 12012 8270 12068
rect 22418 12012 22428 12068
rect 22484 12012 24220 12068
rect 24276 12012 24286 12068
rect 3490 11900 3500 11956
rect 3556 11900 4396 11956
rect 4452 11900 4462 11956
rect 4956 11844 5012 12012
rect 5282 11900 5292 11956
rect 5348 11900 7084 11956
rect 7140 11900 7150 11956
rect 31938 11900 31948 11956
rect 32004 11900 33292 11956
rect 33348 11900 33358 11956
rect 4162 11788 4172 11844
rect 4228 11788 4956 11844
rect 5012 11788 5022 11844
rect 5360 11732 5370 11788
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5634 11732 5644 11788
rect 13676 11732 13686 11788
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13950 11732 13960 11788
rect 21992 11732 22002 11788
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22266 11732 22276 11788
rect 30308 11732 30318 11788
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30582 11732 30592 11788
rect 3714 11676 3724 11732
rect 3780 11676 4732 11732
rect 4788 11676 4798 11732
rect 19058 11676 19068 11732
rect 19124 11676 19134 11732
rect 19618 11676 19628 11732
rect 19684 11676 20076 11732
rect 20132 11676 21308 11732
rect 21364 11676 21374 11732
rect 19068 11620 19124 11676
rect 2482 11564 2492 11620
rect 2548 11564 6524 11620
rect 6580 11564 6590 11620
rect 6850 11564 6860 11620
rect 6916 11564 8540 11620
rect 8596 11564 8606 11620
rect 10434 11564 10444 11620
rect 10500 11564 13020 11620
rect 13076 11564 13086 11620
rect 17266 11564 17276 11620
rect 17332 11564 18172 11620
rect 18228 11564 18238 11620
rect 18956 11564 19124 11620
rect 19842 11564 19852 11620
rect 19908 11564 20412 11620
rect 20468 11564 20478 11620
rect 3042 11452 3052 11508
rect 3108 11452 5572 11508
rect 9202 11452 9212 11508
rect 9268 11452 10892 11508
rect 10948 11452 10958 11508
rect 11330 11452 11340 11508
rect 11396 11452 14252 11508
rect 14308 11452 14318 11508
rect 5516 11396 5572 11452
rect 2146 11340 2156 11396
rect 2212 11340 3500 11396
rect 3556 11340 4732 11396
rect 4788 11340 4798 11396
rect 5506 11340 5516 11396
rect 5572 11340 5582 11396
rect 6290 11340 6300 11396
rect 6356 11340 7084 11396
rect 7140 11340 7150 11396
rect 7970 11340 7980 11396
rect 8036 11340 10444 11396
rect 10500 11340 10510 11396
rect 18956 11284 19012 11564
rect 19170 11452 19180 11508
rect 19236 11452 22540 11508
rect 22596 11452 22606 11508
rect 5954 11228 5964 11284
rect 6020 11228 7420 11284
rect 7476 11228 7486 11284
rect 8978 11228 8988 11284
rect 9044 11228 11116 11284
rect 11172 11228 11182 11284
rect 17490 11228 17500 11284
rect 17556 11228 18508 11284
rect 18564 11228 18574 11284
rect 18722 11228 18732 11284
rect 18788 11228 19012 11284
rect 2594 11116 2604 11172
rect 2660 11116 3612 11172
rect 3668 11116 3678 11172
rect 4834 11116 4844 11172
rect 4900 11116 9324 11172
rect 9380 11116 9996 11172
rect 10052 11116 10062 11172
rect 10434 11116 10444 11172
rect 10500 11116 11340 11172
rect 11396 11116 11406 11172
rect 9518 10948 9528 11004
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9792 10948 9802 11004
rect 17834 10948 17844 11004
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 18108 10948 18118 11004
rect 26150 10948 26160 11004
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26424 10948 26434 11004
rect 34466 10948 34476 11004
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34740 10948 34750 11004
rect 3238 10892 3276 10948
rect 3332 10892 3342 10948
rect 8838 10892 8876 10948
rect 8932 10892 8942 10948
rect 2706 10780 2716 10836
rect 2772 10780 2782 10836
rect 6514 10780 6524 10836
rect 6580 10780 7308 10836
rect 7364 10780 7374 10836
rect 7634 10780 7644 10836
rect 7700 10780 11228 10836
rect 11284 10780 11294 10836
rect 22530 10780 22540 10836
rect 22596 10780 24668 10836
rect 24724 10780 24734 10836
rect 2716 10612 2772 10780
rect 2930 10668 2940 10724
rect 2996 10668 3276 10724
rect 3332 10668 6076 10724
rect 6132 10668 8876 10724
rect 8932 10668 10220 10724
rect 10276 10668 10286 10724
rect 22082 10668 22092 10724
rect 22148 10668 25900 10724
rect 25956 10668 25966 10724
rect 30930 10668 30940 10724
rect 30996 10668 31836 10724
rect 31892 10668 31902 10724
rect 2716 10556 2996 10612
rect 4386 10556 4396 10612
rect 4452 10556 5068 10612
rect 5124 10556 6300 10612
rect 6356 10556 6366 10612
rect 7074 10556 7084 10612
rect 7140 10556 7150 10612
rect 8194 10556 8204 10612
rect 8260 10556 9436 10612
rect 9492 10556 9502 10612
rect 9846 10556 9884 10612
rect 9940 10556 9950 10612
rect 30370 10556 30380 10612
rect 30436 10556 31276 10612
rect 31332 10556 32172 10612
rect 32228 10556 32238 10612
rect 2940 10500 2996 10556
rect 7084 10500 7140 10556
rect 2930 10444 2940 10500
rect 2996 10444 3006 10500
rect 4722 10444 4732 10500
rect 4788 10444 6804 10500
rect 7084 10444 10220 10500
rect 10276 10444 10286 10500
rect 29922 10444 29932 10500
rect 29988 10444 30268 10500
rect 30324 10444 30828 10500
rect 30884 10444 30894 10500
rect 4722 10332 4732 10388
rect 4788 10332 5516 10388
rect 5572 10332 5582 10388
rect 6748 10276 6804 10444
rect 8754 10332 8764 10388
rect 8820 10332 10108 10388
rect 10164 10332 11004 10388
rect 11060 10332 11070 10388
rect 12338 10332 12348 10388
rect 12404 10332 13468 10388
rect 13524 10332 14700 10388
rect 14756 10332 14766 10388
rect 29932 10332 30492 10388
rect 30548 10332 31164 10388
rect 31220 10332 31230 10388
rect 29932 10276 29988 10332
rect 6748 10220 12012 10276
rect 12068 10220 12908 10276
rect 12964 10220 12974 10276
rect 29922 10220 29932 10276
rect 29988 10220 29998 10276
rect 5360 10164 5370 10220
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5634 10164 5644 10220
rect 7382 10108 7420 10164
rect 7476 10108 12236 10164
rect 12292 10108 12302 10164
rect 12908 10052 12964 10220
rect 13676 10164 13686 10220
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13950 10164 13960 10220
rect 21992 10164 22002 10220
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22266 10164 22276 10220
rect 30308 10164 30318 10220
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30582 10164 30592 10220
rect 18498 10108 18508 10164
rect 18564 10108 18844 10164
rect 18900 10108 20972 10164
rect 21028 10108 21420 10164
rect 21476 10108 21588 10164
rect 21532 10052 21588 10108
rect 3042 9996 3052 10052
rect 3108 9996 3612 10052
rect 3668 9996 3678 10052
rect 4918 9996 4956 10052
rect 5012 9996 5022 10052
rect 7522 9996 7532 10052
rect 7588 9996 9212 10052
rect 9268 9996 9278 10052
rect 12908 9996 13692 10052
rect 13748 9996 14924 10052
rect 14980 9996 14990 10052
rect 19730 9996 19740 10052
rect 19796 9996 21308 10052
rect 21364 9996 21374 10052
rect 21532 9996 23100 10052
rect 23156 9996 23166 10052
rect 23650 9996 23660 10052
rect 23716 9996 26908 10052
rect 26964 9996 26974 10052
rect 27122 9996 27132 10052
rect 27188 9996 30716 10052
rect 30772 9996 30782 10052
rect 2594 9884 2604 9940
rect 2660 9884 3164 9940
rect 3220 9884 5628 9940
rect 5684 9884 5694 9940
rect 19170 9884 19180 9940
rect 19236 9884 21420 9940
rect 21476 9884 21486 9940
rect 27794 9884 27804 9940
rect 27860 9884 29484 9940
rect 29540 9884 29550 9940
rect 29708 9884 30940 9940
rect 30996 9884 33068 9940
rect 33124 9884 33134 9940
rect 29708 9828 29764 9884
rect 2706 9772 2716 9828
rect 2772 9772 3276 9828
rect 3332 9772 4060 9828
rect 4116 9772 4126 9828
rect 7074 9772 7084 9828
rect 7140 9772 7868 9828
rect 7924 9772 9548 9828
rect 9604 9772 10556 9828
rect 10612 9772 11452 9828
rect 11508 9772 11518 9828
rect 12898 9772 12908 9828
rect 12964 9772 16828 9828
rect 16884 9772 17836 9828
rect 17892 9772 17902 9828
rect 18610 9772 18620 9828
rect 18676 9772 20076 9828
rect 20132 9772 20636 9828
rect 20692 9772 22092 9828
rect 22148 9772 22158 9828
rect 24658 9772 24668 9828
rect 24724 9772 27244 9828
rect 27300 9772 27310 9828
rect 29138 9772 29148 9828
rect 29204 9772 29708 9828
rect 29764 9772 29774 9828
rect 29922 9772 29932 9828
rect 29988 9772 30380 9828
rect 30436 9772 30446 9828
rect 6178 9660 6188 9716
rect 6244 9660 8764 9716
rect 8820 9660 8830 9716
rect 17602 9660 17612 9716
rect 17668 9660 18956 9716
rect 19012 9660 19022 9716
rect 23090 9660 23100 9716
rect 23156 9660 24444 9716
rect 24500 9660 24510 9716
rect 26786 9660 26796 9716
rect 26852 9604 26908 9716
rect 29362 9660 29372 9716
rect 29428 9660 30156 9716
rect 30212 9660 30222 9716
rect 3714 9548 3724 9604
rect 3780 9548 4956 9604
rect 5012 9548 8988 9604
rect 9044 9548 10556 9604
rect 10612 9548 10622 9604
rect 13570 9548 13580 9604
rect 13636 9548 14140 9604
rect 14196 9548 14206 9604
rect 26852 9548 27916 9604
rect 27972 9548 27982 9604
rect 28466 9548 28476 9604
rect 28532 9548 29260 9604
rect 29316 9548 29326 9604
rect 2930 9436 2940 9492
rect 2996 9436 3500 9492
rect 3556 9436 4284 9492
rect 4340 9436 4350 9492
rect 9518 9380 9528 9436
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9792 9380 9802 9436
rect 17834 9380 17844 9436
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 18108 9380 18118 9436
rect 26150 9380 26160 9436
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 26424 9380 26434 9436
rect 34466 9380 34476 9436
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34740 9380 34750 9436
rect 4610 9212 4620 9268
rect 4676 9212 5852 9268
rect 5908 9212 5918 9268
rect 7074 9212 7084 9268
rect 7140 9212 7308 9268
rect 7364 9212 7374 9268
rect 21858 9212 21868 9268
rect 21924 9212 23996 9268
rect 24052 9212 24062 9268
rect 5506 9100 5516 9156
rect 5572 9100 6524 9156
rect 6580 9100 6590 9156
rect 8978 9100 8988 9156
rect 9044 9100 9212 9156
rect 9268 9100 10220 9156
rect 10276 9100 10286 9156
rect 30706 9100 30716 9156
rect 30772 9100 31388 9156
rect 31444 9100 31836 9156
rect 31892 9100 34076 9156
rect 34132 9100 34142 9156
rect 3938 8988 3948 9044
rect 4004 8988 6412 9044
rect 6468 8988 7756 9044
rect 7812 8988 7822 9044
rect 9958 8988 9996 9044
rect 10052 8988 10062 9044
rect 11554 8988 11564 9044
rect 11620 8988 13020 9044
rect 13076 8988 13086 9044
rect 13794 8988 13804 9044
rect 13860 8988 14140 9044
rect 14196 8988 14588 9044
rect 14644 8988 14654 9044
rect 14914 8988 14924 9044
rect 14980 8988 17724 9044
rect 17780 8988 17790 9044
rect 32162 8988 32172 9044
rect 32228 8988 33292 9044
rect 33348 8988 33358 9044
rect 13020 8932 13076 8988
rect 4274 8876 4284 8932
rect 4340 8876 7980 8932
rect 8036 8876 8046 8932
rect 13020 8876 15148 8932
rect 16594 8876 16604 8932
rect 16660 8876 17948 8932
rect 18004 8876 18956 8932
rect 19012 8876 19022 8932
rect 23762 8876 23772 8932
rect 23828 8876 25340 8932
rect 25396 8876 25406 8932
rect 15092 8820 15148 8876
rect 4050 8764 4060 8820
rect 4116 8764 4172 8820
rect 4228 8764 4238 8820
rect 4834 8764 4844 8820
rect 4900 8764 7084 8820
rect 7140 8764 7150 8820
rect 12460 8764 14980 8820
rect 15092 8764 16044 8820
rect 16100 8764 19068 8820
rect 19124 8764 19134 8820
rect 12460 8708 12516 8764
rect 14924 8708 14980 8764
rect 6850 8652 6860 8708
rect 6916 8652 6972 8708
rect 7028 8652 7644 8708
rect 7700 8652 8876 8708
rect 8932 8652 9548 8708
rect 9604 8652 9614 8708
rect 11218 8652 11228 8708
rect 11284 8652 11676 8708
rect 11732 8652 11742 8708
rect 12450 8652 12460 8708
rect 12516 8652 12526 8708
rect 14924 8652 15148 8708
rect 5360 8596 5370 8652
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5634 8596 5644 8652
rect 13676 8596 13686 8652
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13950 8596 13960 8652
rect 2482 8540 2492 8596
rect 2548 8540 3612 8596
rect 3668 8540 4396 8596
rect 4452 8540 4462 8596
rect 5954 8540 5964 8596
rect 6020 8540 7196 8596
rect 7252 8540 7262 8596
rect 10658 8540 10668 8596
rect 10724 8540 13468 8596
rect 13524 8540 13534 8596
rect 14914 8540 14924 8596
rect 14980 8540 14990 8596
rect 14924 8484 14980 8540
rect 4946 8428 4956 8484
rect 5012 8428 5628 8484
rect 5684 8428 5694 8484
rect 6598 8428 6636 8484
rect 6692 8428 6702 8484
rect 8082 8428 8092 8484
rect 8148 8428 8988 8484
rect 9044 8428 9054 8484
rect 11890 8428 11900 8484
rect 11956 8428 13356 8484
rect 13412 8428 13422 8484
rect 13794 8428 13804 8484
rect 13860 8428 14980 8484
rect 15092 8484 15148 8652
rect 21992 8596 22002 8652
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22266 8596 22276 8652
rect 30308 8596 30318 8652
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30582 8596 30592 8652
rect 15092 8428 15708 8484
rect 15764 8428 15774 8484
rect 29698 8428 29708 8484
rect 29764 8428 30380 8484
rect 30436 8428 30446 8484
rect 2146 8316 2156 8372
rect 2212 8316 3836 8372
rect 3892 8316 3902 8372
rect 4162 8316 4172 8372
rect 4228 8316 6972 8372
rect 7028 8316 10108 8372
rect 10164 8316 10780 8372
rect 10836 8316 10846 8372
rect 33394 8316 33404 8372
rect 33460 8316 34188 8372
rect 34244 8316 34254 8372
rect 4386 8204 4396 8260
rect 4452 8204 4956 8260
rect 5012 8204 6524 8260
rect 6580 8204 6590 8260
rect 6748 8204 9044 8260
rect 9874 8204 9884 8260
rect 9940 8204 11340 8260
rect 11396 8204 11406 8260
rect 12114 8204 12124 8260
rect 12180 8204 13468 8260
rect 13524 8204 14700 8260
rect 14756 8204 15092 8260
rect 25890 8204 25900 8260
rect 25956 8204 26908 8260
rect 26964 8204 26974 8260
rect 29698 8204 29708 8260
rect 29764 8204 30492 8260
rect 30548 8204 30558 8260
rect 6748 8148 6804 8204
rect 8988 8148 9044 8204
rect 15036 8148 15092 8204
rect 2818 8092 2828 8148
rect 2884 8092 3388 8148
rect 3444 8092 4284 8148
rect 4340 8092 6804 8148
rect 7186 8092 7196 8148
rect 7252 8092 7420 8148
rect 7476 8092 7486 8148
rect 8082 8092 8092 8148
rect 8148 8092 8764 8148
rect 8820 8092 8830 8148
rect 8988 8092 11900 8148
rect 11956 8092 11966 8148
rect 15026 8092 15036 8148
rect 15092 8092 15102 8148
rect 28018 8092 28028 8148
rect 28084 8092 29372 8148
rect 29428 8092 29438 8148
rect 2258 7980 2268 8036
rect 2324 7980 4508 8036
rect 4564 7980 4574 8036
rect 5730 7980 5740 8036
rect 5796 7980 9548 8036
rect 9604 7980 9614 8036
rect 9846 7980 9884 8036
rect 9940 7980 9950 8036
rect 21746 7980 21756 8036
rect 21812 7980 23324 8036
rect 23380 7980 23390 8036
rect 6300 7924 6356 7980
rect 4050 7868 4060 7924
rect 4116 7868 5068 7924
rect 5124 7868 5134 7924
rect 6290 7868 6300 7924
rect 6356 7868 6366 7924
rect 7158 7868 7196 7924
rect 7252 7868 8876 7924
rect 8932 7868 8942 7924
rect 13094 7868 13132 7924
rect 13188 7868 13198 7924
rect 13458 7868 13468 7924
rect 13524 7868 15372 7924
rect 15428 7868 16716 7924
rect 16772 7868 16782 7924
rect 9518 7812 9528 7868
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9792 7812 9802 7868
rect 17834 7812 17844 7868
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 18108 7812 18118 7868
rect 26150 7812 26160 7868
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26424 7812 26434 7868
rect 34466 7812 34476 7868
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34740 7812 34750 7868
rect 3826 7756 3836 7812
rect 3892 7756 5740 7812
rect 5796 7756 7308 7812
rect 7364 7756 7374 7812
rect 3938 7644 3948 7700
rect 4004 7644 4172 7700
rect 4228 7644 4238 7700
rect 4498 7644 4508 7700
rect 4564 7644 6076 7700
rect 6132 7644 6142 7700
rect 9762 7644 9772 7700
rect 9828 7644 11116 7700
rect 11172 7644 11182 7700
rect 3490 7532 3500 7588
rect 3556 7532 9436 7588
rect 9492 7532 10108 7588
rect 10164 7532 10174 7588
rect 29474 7532 29484 7588
rect 29540 7532 33404 7588
rect 33460 7532 33470 7588
rect 3602 7420 3612 7476
rect 3668 7420 5292 7476
rect 5348 7420 5358 7476
rect 6850 7420 6860 7476
rect 6916 7420 7868 7476
rect 7924 7420 7934 7476
rect 8866 7420 8876 7476
rect 8932 7420 9884 7476
rect 9940 7420 10556 7476
rect 10612 7420 10622 7476
rect 11414 7420 11452 7476
rect 11508 7420 11518 7476
rect 16818 7420 16828 7476
rect 16884 7420 18732 7476
rect 18788 7420 19180 7476
rect 19236 7420 19246 7476
rect 21634 7420 21644 7476
rect 21700 7420 22204 7476
rect 22260 7420 22540 7476
rect 22596 7420 22606 7476
rect 22978 7420 22988 7476
rect 23044 7420 26236 7476
rect 26292 7420 26302 7476
rect 30258 7420 30268 7476
rect 30324 7420 31052 7476
rect 31108 7420 31724 7476
rect 31780 7420 31790 7476
rect 4834 7308 4844 7364
rect 4900 7308 10444 7364
rect 10500 7308 10510 7364
rect 11890 7308 11900 7364
rect 11956 7308 12684 7364
rect 12740 7308 14476 7364
rect 14532 7308 14542 7364
rect 27682 7308 27692 7364
rect 27748 7308 29148 7364
rect 29204 7308 29214 7364
rect 2818 7196 2828 7252
rect 2884 7196 4172 7252
rect 4228 7196 9884 7252
rect 9940 7196 9950 7252
rect 21522 7196 21532 7252
rect 21588 7196 23772 7252
rect 23828 7196 23838 7252
rect 24098 7196 24108 7252
rect 24164 7196 28028 7252
rect 28084 7196 28094 7252
rect 29250 7196 29260 7252
rect 29316 7196 31724 7252
rect 31780 7196 33516 7252
rect 33572 7196 33582 7252
rect 2594 7084 2604 7140
rect 2660 7084 4172 7140
rect 4228 7084 4238 7140
rect 5730 7084 5740 7140
rect 5796 7084 5834 7140
rect 6626 7084 6636 7140
rect 6692 7084 7644 7140
rect 7700 7084 7710 7140
rect 12226 7084 12236 7140
rect 12292 7084 12796 7140
rect 12852 7084 12862 7140
rect 26852 7084 27692 7140
rect 27748 7084 28252 7140
rect 28308 7084 28318 7140
rect 5360 7028 5370 7084
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5634 7028 5644 7084
rect 2818 6972 2828 7028
rect 2884 6972 4732 7028
rect 4788 6972 4798 7028
rect 5030 6972 5068 7028
rect 5124 6972 5134 7028
rect 6636 6916 6692 7084
rect 13676 7028 13686 7084
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13950 7028 13960 7084
rect 21992 7028 22002 7084
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22266 7028 22276 7084
rect 26852 6916 26908 7084
rect 30308 7028 30318 7084
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30582 7028 30592 7084
rect 3490 6860 3500 6916
rect 3556 6860 4844 6916
rect 4900 6860 4910 6916
rect 5170 6860 5180 6916
rect 5236 6860 6692 6916
rect 22082 6860 22092 6916
rect 22148 6860 23324 6916
rect 23380 6860 23548 6916
rect 23604 6860 23614 6916
rect 26002 6860 26012 6916
rect 26068 6860 26908 6916
rect 30706 6860 30716 6916
rect 30772 6860 31612 6916
rect 31668 6860 33068 6916
rect 33124 6860 33134 6916
rect 5058 6748 5068 6804
rect 5124 6748 5628 6804
rect 5684 6748 5694 6804
rect 9650 6748 9660 6804
rect 9716 6748 9996 6804
rect 10052 6748 10062 6804
rect 10994 6748 11004 6804
rect 11060 6748 12124 6804
rect 12180 6748 12190 6804
rect 19170 6748 19180 6804
rect 19236 6748 19740 6804
rect 19796 6748 19806 6804
rect 21858 6748 21868 6804
rect 21924 6748 23436 6804
rect 23492 6748 23502 6804
rect 26674 6748 26684 6804
rect 26740 6748 28700 6804
rect 28756 6748 29372 6804
rect 29428 6748 29438 6804
rect 29698 6748 29708 6804
rect 29764 6748 30044 6804
rect 30100 6748 30380 6804
rect 30436 6748 30446 6804
rect 9090 6636 9100 6692
rect 9156 6636 9772 6692
rect 9828 6636 11788 6692
rect 11844 6636 11854 6692
rect 13122 6636 13132 6692
rect 13188 6636 17164 6692
rect 17220 6636 17230 6692
rect 22194 6636 22204 6692
rect 22260 6636 23660 6692
rect 23716 6636 23726 6692
rect 26450 6636 26460 6692
rect 26516 6636 29932 6692
rect 29988 6636 29998 6692
rect 5730 6524 5740 6580
rect 5796 6524 8204 6580
rect 8260 6524 8270 6580
rect 9986 6524 9996 6580
rect 10052 6524 10220 6580
rect 10276 6524 10780 6580
rect 10836 6524 12348 6580
rect 12404 6524 12414 6580
rect 22978 6524 22988 6580
rect 23044 6524 24780 6580
rect 24836 6524 24846 6580
rect 25330 6524 25340 6580
rect 25396 6524 27244 6580
rect 27300 6524 27310 6580
rect 3602 6412 3612 6468
rect 3668 6412 4620 6468
rect 4676 6412 6188 6468
rect 6244 6412 6254 6468
rect 6402 6412 6412 6468
rect 6468 6412 7420 6468
rect 7476 6412 7486 6468
rect 7858 6412 7868 6468
rect 7924 6412 8316 6468
rect 8372 6412 8382 6468
rect 3910 6300 3948 6356
rect 4004 6300 4014 6356
rect 12338 6300 12348 6356
rect 12404 6300 13804 6356
rect 13860 6300 13870 6356
rect 9518 6244 9528 6300
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9792 6244 9802 6300
rect 17834 6244 17844 6300
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 18108 6244 18118 6300
rect 26150 6244 26160 6300
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26424 6244 26434 6300
rect 34466 6244 34476 6300
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34740 6244 34750 6300
rect 6514 6188 6524 6244
rect 6580 6188 7084 6244
rect 7140 6188 8540 6244
rect 8596 6188 8606 6244
rect 11106 6188 11116 6244
rect 11172 6188 13860 6244
rect 14130 6188 14140 6244
rect 14196 6188 14812 6244
rect 14868 6188 14878 6244
rect 15092 6188 16044 6244
rect 16100 6188 16110 6244
rect 29922 6188 29932 6244
rect 29988 6188 30156 6244
rect 30212 6188 33068 6244
rect 33124 6188 33134 6244
rect 13804 6132 13860 6188
rect 15092 6132 15148 6188
rect 2930 6076 2940 6132
rect 2996 6076 3276 6132
rect 3332 6076 7868 6132
rect 7924 6076 7934 6132
rect 8194 6076 8204 6132
rect 8260 6076 13580 6132
rect 13636 6076 13646 6132
rect 13804 6076 15148 6132
rect 15474 6076 15484 6132
rect 15540 6076 17948 6132
rect 18004 6076 18956 6132
rect 19012 6076 19022 6132
rect 19506 6076 19516 6132
rect 19572 6076 21308 6132
rect 21364 6076 21374 6132
rect 7868 6020 7924 6076
rect 5282 5964 5292 6020
rect 5348 5964 6188 6020
rect 6244 5964 6254 6020
rect 7868 5964 8428 6020
rect 8484 5964 8494 6020
rect 11106 5964 11116 6020
rect 11172 5964 11452 6020
rect 11508 5964 11788 6020
rect 12450 5964 12460 6020
rect 12516 5964 13692 6020
rect 13748 5964 13758 6020
rect 14690 5964 14700 6020
rect 14756 5964 17388 6020
rect 17444 5964 17454 6020
rect 20066 5964 20076 6020
rect 20132 5964 20524 6020
rect 20580 5964 20972 6020
rect 21028 5964 21420 6020
rect 21476 5964 21486 6020
rect 21634 5964 21644 6020
rect 21700 5964 22988 6020
rect 23044 5964 23054 6020
rect 24210 5964 24220 6020
rect 24276 5964 25452 6020
rect 25508 5964 26908 6020
rect 26964 5964 26974 6020
rect 30930 5964 30940 6020
rect 30996 5964 33404 6020
rect 33460 5964 33470 6020
rect 2594 5852 2604 5908
rect 2660 5852 3052 5908
rect 3108 5852 3118 5908
rect 4386 5852 4396 5908
rect 4452 5852 7644 5908
rect 7700 5852 8764 5908
rect 8820 5852 9324 5908
rect 9380 5852 9390 5908
rect 11732 5796 11788 5964
rect 12786 5852 12796 5908
rect 12852 5852 14252 5908
rect 14308 5852 14318 5908
rect 14578 5852 14588 5908
rect 14644 5852 14654 5908
rect 14802 5852 14812 5908
rect 14868 5852 16156 5908
rect 16212 5852 16222 5908
rect 19282 5852 19292 5908
rect 19348 5852 21532 5908
rect 21588 5852 21598 5908
rect 24098 5852 24108 5908
rect 24164 5852 25228 5908
rect 25284 5852 25294 5908
rect 25564 5852 26796 5908
rect 26852 5852 26862 5908
rect 27356 5852 27468 5908
rect 27524 5852 27534 5908
rect 29810 5852 29820 5908
rect 29876 5852 31164 5908
rect 31220 5852 32956 5908
rect 33012 5852 33022 5908
rect 14588 5796 14644 5852
rect 25564 5796 25620 5852
rect 27356 5796 27412 5852
rect 4050 5740 4060 5796
rect 4116 5740 5964 5796
rect 6020 5740 8204 5796
rect 8260 5740 8876 5796
rect 8932 5740 8942 5796
rect 11732 5740 12628 5796
rect 14588 5740 17500 5796
rect 17556 5740 17566 5796
rect 24322 5740 24332 5796
rect 24388 5740 25564 5796
rect 25620 5740 25630 5796
rect 26002 5740 26012 5796
rect 26068 5740 27412 5796
rect 27570 5740 27580 5796
rect 27636 5740 27646 5796
rect 31714 5740 31724 5796
rect 31780 5740 33180 5796
rect 33236 5740 33246 5796
rect 12572 5684 12628 5740
rect 27580 5684 27636 5740
rect 5842 5628 5852 5684
rect 5908 5628 8092 5684
rect 8148 5628 8158 5684
rect 9314 5628 9324 5684
rect 9380 5628 11564 5684
rect 11620 5628 11630 5684
rect 12572 5628 16268 5684
rect 16324 5628 16334 5684
rect 26786 5628 26796 5684
rect 26852 5628 27636 5684
rect 8530 5516 8540 5572
rect 8596 5516 10668 5572
rect 10724 5516 11452 5572
rect 11508 5516 11518 5572
rect 5360 5460 5370 5516
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5634 5460 5644 5516
rect 13676 5460 13686 5516
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13950 5460 13960 5516
rect 21992 5460 22002 5516
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22266 5460 22276 5516
rect 30308 5460 30318 5516
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30582 5460 30592 5516
rect 5730 5404 5740 5460
rect 5796 5404 7980 5460
rect 8036 5404 10108 5460
rect 10164 5404 10174 5460
rect 10518 5404 10556 5460
rect 10612 5404 10622 5460
rect 4610 5292 4620 5348
rect 4676 5292 5180 5348
rect 5236 5292 5246 5348
rect 8418 5292 8428 5348
rect 8484 5292 10220 5348
rect 10276 5292 13692 5348
rect 13748 5292 13758 5348
rect 5058 5180 5068 5236
rect 5124 5180 6188 5236
rect 6244 5180 8652 5236
rect 8708 5180 11396 5236
rect 11778 5180 11788 5236
rect 11844 5180 12460 5236
rect 12516 5180 12526 5236
rect 18274 5180 18284 5236
rect 18340 5180 19180 5236
rect 19236 5180 19246 5236
rect 21634 5180 21644 5236
rect 21700 5180 23772 5236
rect 23828 5180 26908 5236
rect 26964 5180 27804 5236
rect 27860 5180 27870 5236
rect 30594 5180 30604 5236
rect 30660 5180 31836 5236
rect 31892 5180 31902 5236
rect 33506 5180 33516 5236
rect 33572 5180 34188 5236
rect 34244 5180 34254 5236
rect 11340 5124 11396 5180
rect 2482 5068 2492 5124
rect 2548 5068 4284 5124
rect 4340 5068 4676 5124
rect 4834 5068 4844 5124
rect 4900 5068 5964 5124
rect 6020 5068 6030 5124
rect 8866 5068 8876 5124
rect 8932 5068 11004 5124
rect 11060 5068 11070 5124
rect 11330 5068 11340 5124
rect 11396 5068 12124 5124
rect 12180 5068 12190 5124
rect 12674 5068 12684 5124
rect 12740 5068 13132 5124
rect 13188 5068 13916 5124
rect 13972 5068 13982 5124
rect 16930 5068 16940 5124
rect 16996 5068 18172 5124
rect 18228 5068 18732 5124
rect 18788 5068 18798 5124
rect 27010 5068 27020 5124
rect 27076 5068 28756 5124
rect 29698 5068 29708 5124
rect 29764 5068 30380 5124
rect 30436 5068 30446 5124
rect 4620 5012 4676 5068
rect 28700 5012 28756 5068
rect 4620 4956 6076 5012
rect 6132 4956 6860 5012
rect 6916 4956 6926 5012
rect 7298 4956 7308 5012
rect 7364 4956 8204 5012
rect 8260 4956 8270 5012
rect 8530 4956 8540 5012
rect 8596 4956 11788 5012
rect 11844 4956 13356 5012
rect 13412 4956 13422 5012
rect 15092 4956 17724 5012
rect 17780 4956 18620 5012
rect 18676 4956 18686 5012
rect 18834 4956 18844 5012
rect 18900 4956 19516 5012
rect 19572 4956 19582 5012
rect 22754 4956 22764 5012
rect 22820 4956 23436 5012
rect 23492 4956 23502 5012
rect 26226 4956 26236 5012
rect 26292 4956 26908 5012
rect 28690 4956 28700 5012
rect 28756 4956 31276 5012
rect 31332 4956 31948 5012
rect 32004 4956 32014 5012
rect 15092 4900 15148 4956
rect 6626 4844 6636 4900
rect 6692 4844 7644 4900
rect 7700 4844 7710 4900
rect 13570 4844 13580 4900
rect 13636 4844 14476 4900
rect 14532 4844 15148 4900
rect 26852 4900 26908 4956
rect 26852 4844 27468 4900
rect 27524 4844 27534 4900
rect 29586 4844 29596 4900
rect 29652 4844 31164 4900
rect 31220 4844 31230 4900
rect 9518 4676 9528 4732
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9792 4676 9802 4732
rect 17834 4676 17844 4732
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 18108 4676 18118 4732
rect 26150 4676 26160 4732
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26424 4676 26434 4732
rect 34466 4676 34476 4732
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34740 4676 34750 4732
rect 4694 4508 4732 4564
rect 4788 4508 4798 4564
rect 7606 4508 7644 4564
rect 7700 4508 8540 4564
rect 8596 4508 8606 4564
rect 8978 4508 8988 4564
rect 9044 4508 11228 4564
rect 11284 4508 12124 4564
rect 12180 4508 13468 4564
rect 13524 4508 13534 4564
rect 16258 4508 16268 4564
rect 16324 4508 17276 4564
rect 17332 4508 17342 4564
rect 18050 4508 18060 4564
rect 18116 4508 19068 4564
rect 19124 4508 19134 4564
rect 21858 4508 21868 4564
rect 21924 4508 22764 4564
rect 22820 4508 22830 4564
rect 3602 4396 3612 4452
rect 3668 4396 6972 4452
rect 7028 4396 14924 4452
rect 14980 4396 14990 4452
rect 1810 4284 1820 4340
rect 1876 4284 5740 4340
rect 5796 4284 6748 4340
rect 6804 4284 6814 4340
rect 8754 4284 8764 4340
rect 8820 4284 10668 4340
rect 10724 4284 10734 4340
rect 12562 4284 12572 4340
rect 12628 4284 15036 4340
rect 15092 4284 15102 4340
rect 16818 4284 16828 4340
rect 16884 4284 17612 4340
rect 17668 4284 17678 4340
rect 21746 4284 21756 4340
rect 21812 4284 23100 4340
rect 23156 4284 23166 4340
rect 1586 4172 1596 4228
rect 1652 4172 3612 4228
rect 3668 4172 3678 4228
rect 6822 4172 6860 4228
rect 6916 4172 6926 4228
rect 20290 4172 20300 4228
rect 20356 4172 23660 4228
rect 23716 4172 23726 4228
rect 6402 4060 6412 4116
rect 6468 4060 6972 4116
rect 7028 4060 7038 4116
rect 7858 4060 7868 4116
rect 7924 4060 10220 4116
rect 10276 4060 10286 4116
rect 23314 4060 23324 4116
rect 23380 4060 25228 4116
rect 25284 4060 25294 4116
rect 5360 3892 5370 3948
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5634 3892 5644 3948
rect 13676 3892 13686 3948
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13950 3892 13960 3948
rect 21992 3892 22002 3948
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22266 3892 22276 3948
rect 30308 3892 30318 3948
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30582 3892 30592 3948
rect 14130 3724 14140 3780
rect 14196 3724 15260 3780
rect 15316 3724 15326 3780
rect 5170 3612 5180 3668
rect 5236 3612 6748 3668
rect 6804 3612 15372 3668
rect 15428 3612 15438 3668
rect 22754 3612 22764 3668
rect 22820 3612 24556 3668
rect 24612 3612 24622 3668
rect 9538 3500 9548 3556
rect 9604 3500 12572 3556
rect 12628 3500 12638 3556
rect 14354 3500 14364 3556
rect 14420 3500 15484 3556
rect 15540 3500 15550 3556
rect 19730 3500 19740 3556
rect 19796 3500 20748 3556
rect 20804 3500 20814 3556
rect 22418 3500 22428 3556
rect 22484 3500 24892 3556
rect 24948 3500 24958 3556
rect 31490 3500 31500 3556
rect 31556 3500 32172 3556
rect 32228 3500 32238 3556
rect 10770 3388 10780 3444
rect 10836 3388 13244 3444
rect 13300 3388 13310 3444
rect 25106 3388 25116 3444
rect 25172 3388 26908 3444
rect 26964 3388 26974 3444
rect 30034 3388 30044 3444
rect 30100 3388 32284 3444
rect 32340 3388 32350 3444
rect 8194 3276 8204 3332
rect 8260 3276 11900 3332
rect 11956 3276 11966 3332
rect 9518 3108 9528 3164
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9792 3108 9802 3164
rect 17834 3108 17844 3164
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 18108 3108 18118 3164
rect 26150 3108 26160 3164
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26424 3108 26434 3164
rect 34466 3108 34476 3164
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34740 3108 34750 3164
rect 11732 2996 11788 3108
rect 11844 3052 13132 3108
rect 13188 3052 13198 3108
rect 6402 2940 6412 2996
rect 6468 2940 11788 2996
<< via3 >>
rect 5370 32116 5426 32172
rect 5474 32116 5530 32172
rect 5578 32116 5634 32172
rect 13686 32116 13742 32172
rect 13790 32116 13846 32172
rect 13894 32116 13950 32172
rect 22002 32116 22058 32172
rect 22106 32116 22162 32172
rect 22210 32116 22266 32172
rect 30318 32116 30374 32172
rect 30422 32116 30478 32172
rect 30526 32116 30582 32172
rect 9528 31332 9584 31388
rect 9632 31332 9688 31388
rect 9736 31332 9792 31388
rect 17844 31332 17900 31388
rect 17948 31332 18004 31388
rect 18052 31332 18108 31388
rect 26160 31332 26216 31388
rect 26264 31332 26320 31388
rect 26368 31332 26424 31388
rect 34476 31332 34532 31388
rect 34580 31332 34636 31388
rect 34684 31332 34740 31388
rect 5370 30548 5426 30604
rect 5474 30548 5530 30604
rect 5578 30548 5634 30604
rect 13686 30548 13742 30604
rect 13790 30548 13846 30604
rect 13894 30548 13950 30604
rect 22002 30548 22058 30604
rect 22106 30548 22162 30604
rect 22210 30548 22266 30604
rect 30318 30548 30374 30604
rect 30422 30548 30478 30604
rect 30526 30548 30582 30604
rect 9528 29764 9584 29820
rect 9632 29764 9688 29820
rect 9736 29764 9792 29820
rect 17844 29764 17900 29820
rect 17948 29764 18004 29820
rect 18052 29764 18108 29820
rect 26160 29764 26216 29820
rect 26264 29764 26320 29820
rect 26368 29764 26424 29820
rect 34476 29764 34532 29820
rect 34580 29764 34636 29820
rect 34684 29764 34740 29820
rect 5370 28980 5426 29036
rect 5474 28980 5530 29036
rect 5578 28980 5634 29036
rect 13686 28980 13742 29036
rect 13790 28980 13846 29036
rect 13894 28980 13950 29036
rect 22002 28980 22058 29036
rect 22106 28980 22162 29036
rect 22210 28980 22266 29036
rect 30318 28980 30374 29036
rect 30422 28980 30478 29036
rect 30526 28980 30582 29036
rect 9528 28196 9584 28252
rect 9632 28196 9688 28252
rect 9736 28196 9792 28252
rect 17844 28196 17900 28252
rect 17948 28196 18004 28252
rect 18052 28196 18108 28252
rect 26160 28196 26216 28252
rect 26264 28196 26320 28252
rect 26368 28196 26424 28252
rect 34476 28196 34532 28252
rect 34580 28196 34636 28252
rect 34684 28196 34740 28252
rect 5370 27412 5426 27468
rect 5474 27412 5530 27468
rect 5578 27412 5634 27468
rect 13686 27412 13742 27468
rect 13790 27412 13846 27468
rect 13894 27412 13950 27468
rect 22002 27412 22058 27468
rect 22106 27412 22162 27468
rect 22210 27412 22266 27468
rect 30318 27412 30374 27468
rect 30422 27412 30478 27468
rect 30526 27412 30582 27468
rect 9528 26628 9584 26684
rect 9632 26628 9688 26684
rect 9736 26628 9792 26684
rect 17844 26628 17900 26684
rect 17948 26628 18004 26684
rect 18052 26628 18108 26684
rect 26160 26628 26216 26684
rect 26264 26628 26320 26684
rect 26368 26628 26424 26684
rect 34476 26628 34532 26684
rect 34580 26628 34636 26684
rect 34684 26628 34740 26684
rect 5370 25844 5426 25900
rect 5474 25844 5530 25900
rect 5578 25844 5634 25900
rect 13686 25844 13742 25900
rect 13790 25844 13846 25900
rect 13894 25844 13950 25900
rect 22002 25844 22058 25900
rect 22106 25844 22162 25900
rect 22210 25844 22266 25900
rect 30318 25844 30374 25900
rect 30422 25844 30478 25900
rect 30526 25844 30582 25900
rect 12348 25452 12404 25508
rect 12460 25340 12516 25396
rect 9528 25060 9584 25116
rect 9632 25060 9688 25116
rect 9736 25060 9792 25116
rect 17844 25060 17900 25116
rect 17948 25060 18004 25116
rect 18052 25060 18108 25116
rect 26160 25060 26216 25116
rect 26264 25060 26320 25116
rect 26368 25060 26424 25116
rect 34476 25060 34532 25116
rect 34580 25060 34636 25116
rect 34684 25060 34740 25116
rect 12236 24668 12292 24724
rect 12460 24668 12516 24724
rect 14588 24668 14644 24724
rect 5370 24276 5426 24332
rect 5474 24276 5530 24332
rect 5578 24276 5634 24332
rect 13686 24276 13742 24332
rect 13790 24276 13846 24332
rect 13894 24276 13950 24332
rect 22002 24276 22058 24332
rect 22106 24276 22162 24332
rect 22210 24276 22266 24332
rect 30318 24276 30374 24332
rect 30422 24276 30478 24332
rect 30526 24276 30582 24332
rect 11900 23996 11956 24052
rect 13468 23996 13524 24052
rect 12236 23772 12292 23828
rect 12572 23772 12628 23828
rect 9528 23492 9584 23548
rect 9632 23492 9688 23548
rect 9736 23492 9792 23548
rect 11900 23548 11956 23604
rect 12348 23548 12404 23604
rect 12572 23548 12628 23604
rect 13468 23548 13524 23604
rect 17844 23492 17900 23548
rect 17948 23492 18004 23548
rect 18052 23492 18108 23548
rect 26160 23492 26216 23548
rect 26264 23492 26320 23548
rect 26368 23492 26424 23548
rect 34476 23492 34532 23548
rect 34580 23492 34636 23548
rect 34684 23492 34740 23548
rect 11228 23436 11284 23492
rect 11228 22764 11284 22820
rect 5370 22708 5426 22764
rect 5474 22708 5530 22764
rect 5578 22708 5634 22764
rect 13686 22708 13742 22764
rect 13790 22708 13846 22764
rect 13894 22708 13950 22764
rect 22002 22708 22058 22764
rect 22106 22708 22162 22764
rect 22210 22708 22266 22764
rect 30318 22708 30374 22764
rect 30422 22708 30478 22764
rect 30526 22708 30582 22764
rect 9528 21924 9584 21980
rect 9632 21924 9688 21980
rect 9736 21924 9792 21980
rect 17844 21924 17900 21980
rect 17948 21924 18004 21980
rect 18052 21924 18108 21980
rect 26160 21924 26216 21980
rect 26264 21924 26320 21980
rect 26368 21924 26424 21980
rect 34476 21924 34532 21980
rect 34580 21924 34636 21980
rect 34684 21924 34740 21980
rect 5370 21140 5426 21196
rect 5474 21140 5530 21196
rect 5578 21140 5634 21196
rect 13686 21140 13742 21196
rect 13790 21140 13846 21196
rect 13894 21140 13950 21196
rect 22002 21140 22058 21196
rect 22106 21140 22162 21196
rect 22210 21140 22266 21196
rect 30318 21140 30374 21196
rect 30422 21140 30478 21196
rect 30526 21140 30582 21196
rect 9528 20356 9584 20412
rect 9632 20356 9688 20412
rect 9736 20356 9792 20412
rect 17844 20356 17900 20412
rect 17948 20356 18004 20412
rect 18052 20356 18108 20412
rect 26160 20356 26216 20412
rect 26264 20356 26320 20412
rect 26368 20356 26424 20412
rect 34476 20356 34532 20412
rect 34580 20356 34636 20412
rect 34684 20356 34740 20412
rect 14588 19852 14644 19908
rect 5370 19572 5426 19628
rect 5474 19572 5530 19628
rect 5578 19572 5634 19628
rect 13686 19572 13742 19628
rect 13790 19572 13846 19628
rect 13894 19572 13950 19628
rect 22002 19572 22058 19628
rect 22106 19572 22162 19628
rect 22210 19572 22266 19628
rect 30318 19572 30374 19628
rect 30422 19572 30478 19628
rect 30526 19572 30582 19628
rect 9528 18788 9584 18844
rect 9632 18788 9688 18844
rect 9736 18788 9792 18844
rect 17844 18788 17900 18844
rect 17948 18788 18004 18844
rect 18052 18788 18108 18844
rect 26160 18788 26216 18844
rect 26264 18788 26320 18844
rect 26368 18788 26424 18844
rect 34476 18788 34532 18844
rect 34580 18788 34636 18844
rect 34684 18788 34740 18844
rect 11116 18732 11172 18788
rect 5370 18004 5426 18060
rect 5474 18004 5530 18060
rect 5578 18004 5634 18060
rect 13686 18004 13742 18060
rect 13790 18004 13846 18060
rect 13894 18004 13950 18060
rect 22002 18004 22058 18060
rect 22106 18004 22162 18060
rect 22210 18004 22266 18060
rect 30318 18004 30374 18060
rect 30422 18004 30478 18060
rect 30526 18004 30582 18060
rect 11116 17724 11172 17780
rect 17052 17724 17108 17780
rect 9528 17220 9584 17276
rect 9632 17220 9688 17276
rect 9736 17220 9792 17276
rect 17844 17220 17900 17276
rect 17948 17220 18004 17276
rect 18052 17220 18108 17276
rect 26160 17220 26216 17276
rect 26264 17220 26320 17276
rect 26368 17220 26424 17276
rect 34476 17220 34532 17276
rect 34580 17220 34636 17276
rect 34684 17220 34740 17276
rect 17052 16828 17108 16884
rect 5370 16436 5426 16492
rect 5474 16436 5530 16492
rect 5578 16436 5634 16492
rect 13686 16436 13742 16492
rect 13790 16436 13846 16492
rect 13894 16436 13950 16492
rect 22002 16436 22058 16492
rect 22106 16436 22162 16492
rect 22210 16436 22266 16492
rect 30318 16436 30374 16492
rect 30422 16436 30478 16492
rect 30526 16436 30582 16492
rect 9528 15652 9584 15708
rect 9632 15652 9688 15708
rect 9736 15652 9792 15708
rect 17844 15652 17900 15708
rect 17948 15652 18004 15708
rect 18052 15652 18108 15708
rect 26160 15652 26216 15708
rect 26264 15652 26320 15708
rect 26368 15652 26424 15708
rect 34476 15652 34532 15708
rect 34580 15652 34636 15708
rect 34684 15652 34740 15708
rect 5370 14868 5426 14924
rect 5474 14868 5530 14924
rect 5578 14868 5634 14924
rect 13686 14868 13742 14924
rect 13790 14868 13846 14924
rect 13894 14868 13950 14924
rect 22002 14868 22058 14924
rect 22106 14868 22162 14924
rect 22210 14868 22266 14924
rect 30318 14868 30374 14924
rect 30422 14868 30478 14924
rect 30526 14868 30582 14924
rect 9528 14084 9584 14140
rect 9632 14084 9688 14140
rect 9736 14084 9792 14140
rect 17844 14084 17900 14140
rect 17948 14084 18004 14140
rect 18052 14084 18108 14140
rect 26160 14084 26216 14140
rect 26264 14084 26320 14140
rect 26368 14084 26424 14140
rect 34476 14084 34532 14140
rect 34580 14084 34636 14140
rect 34684 14084 34740 14140
rect 5370 13300 5426 13356
rect 5474 13300 5530 13356
rect 5578 13300 5634 13356
rect 13686 13300 13742 13356
rect 13790 13300 13846 13356
rect 13894 13300 13950 13356
rect 22002 13300 22058 13356
rect 22106 13300 22162 13356
rect 22210 13300 22266 13356
rect 30318 13300 30374 13356
rect 30422 13300 30478 13356
rect 30526 13300 30582 13356
rect 9528 12516 9584 12572
rect 9632 12516 9688 12572
rect 9736 12516 9792 12572
rect 17844 12516 17900 12572
rect 17948 12516 18004 12572
rect 18052 12516 18108 12572
rect 26160 12516 26216 12572
rect 26264 12516 26320 12572
rect 26368 12516 26424 12572
rect 34476 12516 34532 12572
rect 34580 12516 34636 12572
rect 34684 12516 34740 12572
rect 5370 11732 5426 11788
rect 5474 11732 5530 11788
rect 5578 11732 5634 11788
rect 13686 11732 13742 11788
rect 13790 11732 13846 11788
rect 13894 11732 13950 11788
rect 22002 11732 22058 11788
rect 22106 11732 22162 11788
rect 22210 11732 22266 11788
rect 30318 11732 30374 11788
rect 30422 11732 30478 11788
rect 30526 11732 30582 11788
rect 4732 11676 4788 11732
rect 9528 10948 9584 11004
rect 9632 10948 9688 11004
rect 9736 10948 9792 11004
rect 17844 10948 17900 11004
rect 17948 10948 18004 11004
rect 18052 10948 18108 11004
rect 26160 10948 26216 11004
rect 26264 10948 26320 11004
rect 26368 10948 26424 11004
rect 34476 10948 34532 11004
rect 34580 10948 34636 11004
rect 34684 10948 34740 11004
rect 3276 10892 3332 10948
rect 8876 10892 8932 10948
rect 9884 10556 9940 10612
rect 4732 10444 4788 10500
rect 10108 10332 10164 10388
rect 5370 10164 5426 10220
rect 5474 10164 5530 10220
rect 5578 10164 5634 10220
rect 7420 10108 7476 10164
rect 13686 10164 13742 10220
rect 13790 10164 13846 10220
rect 13894 10164 13950 10220
rect 22002 10164 22058 10220
rect 22106 10164 22162 10220
rect 22210 10164 22266 10220
rect 30318 10164 30374 10220
rect 30422 10164 30478 10220
rect 30526 10164 30582 10220
rect 4956 9996 5012 10052
rect 3276 9772 3332 9828
rect 10556 9772 10612 9828
rect 9528 9380 9584 9436
rect 9632 9380 9688 9436
rect 9736 9380 9792 9436
rect 17844 9380 17900 9436
rect 17948 9380 18004 9436
rect 18052 9380 18108 9436
rect 26160 9380 26216 9436
rect 26264 9380 26320 9436
rect 26368 9380 26424 9436
rect 34476 9380 34532 9436
rect 34580 9380 34636 9436
rect 34684 9380 34740 9436
rect 9996 8988 10052 9044
rect 4172 8764 4228 8820
rect 6860 8652 6916 8708
rect 8876 8652 8932 8708
rect 5370 8596 5426 8652
rect 5474 8596 5530 8652
rect 5578 8596 5634 8652
rect 13686 8596 13742 8652
rect 13790 8596 13846 8652
rect 13894 8596 13950 8652
rect 7196 8540 7252 8596
rect 6636 8428 6692 8484
rect 22002 8596 22058 8652
rect 22106 8596 22162 8652
rect 22210 8596 22266 8652
rect 30318 8596 30374 8652
rect 30422 8596 30478 8652
rect 30526 8596 30582 8652
rect 4956 8204 5012 8260
rect 9884 7980 9940 8036
rect 5068 7868 5124 7924
rect 7196 7868 7252 7924
rect 13132 7868 13188 7924
rect 9528 7812 9584 7868
rect 9632 7812 9688 7868
rect 9736 7812 9792 7868
rect 17844 7812 17900 7868
rect 17948 7812 18004 7868
rect 18052 7812 18108 7868
rect 26160 7812 26216 7868
rect 26264 7812 26320 7868
rect 26368 7812 26424 7868
rect 34476 7812 34532 7868
rect 34580 7812 34636 7868
rect 34684 7812 34740 7868
rect 3948 7644 4004 7700
rect 11452 7420 11508 7476
rect 4172 7196 4228 7252
rect 5740 7084 5796 7140
rect 7644 7084 7700 7140
rect 5370 7028 5426 7084
rect 5474 7028 5530 7084
rect 5578 7028 5634 7084
rect 5068 6972 5124 7028
rect 13686 7028 13742 7084
rect 13790 7028 13846 7084
rect 13894 7028 13950 7084
rect 22002 7028 22058 7084
rect 22106 7028 22162 7084
rect 22210 7028 22266 7084
rect 30318 7028 30374 7084
rect 30422 7028 30478 7084
rect 30526 7028 30582 7084
rect 9996 6748 10052 6804
rect 7420 6412 7476 6468
rect 3948 6300 4004 6356
rect 9528 6244 9584 6300
rect 9632 6244 9688 6300
rect 9736 6244 9792 6300
rect 17844 6244 17900 6300
rect 17948 6244 18004 6300
rect 18052 6244 18108 6300
rect 26160 6244 26216 6300
rect 26264 6244 26320 6300
rect 26368 6244 26424 6300
rect 34476 6244 34532 6300
rect 34580 6244 34636 6300
rect 34684 6244 34740 6300
rect 11452 5964 11508 6020
rect 5370 5460 5426 5516
rect 5474 5460 5530 5516
rect 5578 5460 5634 5516
rect 13686 5460 13742 5516
rect 13790 5460 13846 5516
rect 13894 5460 13950 5516
rect 22002 5460 22058 5516
rect 22106 5460 22162 5516
rect 22210 5460 22266 5516
rect 30318 5460 30374 5516
rect 30422 5460 30478 5516
rect 30526 5460 30582 5516
rect 5740 5404 5796 5460
rect 10108 5404 10164 5460
rect 10556 5404 10612 5460
rect 6636 4844 6692 4900
rect 9528 4676 9584 4732
rect 9632 4676 9688 4732
rect 9736 4676 9792 4732
rect 17844 4676 17900 4732
rect 17948 4676 18004 4732
rect 18052 4676 18108 4732
rect 26160 4676 26216 4732
rect 26264 4676 26320 4732
rect 26368 4676 26424 4732
rect 34476 4676 34532 4732
rect 34580 4676 34636 4732
rect 34684 4676 34740 4732
rect 4732 4508 4788 4564
rect 7644 4508 7700 4564
rect 6860 4172 6916 4228
rect 5370 3892 5426 3948
rect 5474 3892 5530 3948
rect 5578 3892 5634 3948
rect 13686 3892 13742 3948
rect 13790 3892 13846 3948
rect 13894 3892 13950 3948
rect 22002 3892 22058 3948
rect 22106 3892 22162 3948
rect 22210 3892 22266 3948
rect 30318 3892 30374 3948
rect 30422 3892 30478 3948
rect 30526 3892 30582 3948
rect 9528 3108 9584 3164
rect 9632 3108 9688 3164
rect 9736 3108 9792 3164
rect 17844 3108 17900 3164
rect 17948 3108 18004 3164
rect 18052 3108 18108 3164
rect 26160 3108 26216 3164
rect 26264 3108 26320 3164
rect 26368 3108 26424 3164
rect 34476 3108 34532 3164
rect 34580 3108 34636 3164
rect 34684 3108 34740 3164
rect 13132 3052 13188 3108
<< metal4 >>
rect 5342 32172 5662 32204
rect 5342 32116 5370 32172
rect 5426 32116 5474 32172
rect 5530 32116 5578 32172
rect 5634 32116 5662 32172
rect 5342 30604 5662 32116
rect 5342 30548 5370 30604
rect 5426 30548 5474 30604
rect 5530 30548 5578 30604
rect 5634 30548 5662 30604
rect 5342 29036 5662 30548
rect 5342 28980 5370 29036
rect 5426 28980 5474 29036
rect 5530 28980 5578 29036
rect 5634 28980 5662 29036
rect 5342 27468 5662 28980
rect 5342 27412 5370 27468
rect 5426 27412 5474 27468
rect 5530 27412 5578 27468
rect 5634 27412 5662 27468
rect 5342 25900 5662 27412
rect 5342 25844 5370 25900
rect 5426 25844 5474 25900
rect 5530 25844 5578 25900
rect 5634 25844 5662 25900
rect 5342 24332 5662 25844
rect 5342 24276 5370 24332
rect 5426 24276 5474 24332
rect 5530 24276 5578 24332
rect 5634 24276 5662 24332
rect 5342 22764 5662 24276
rect 5342 22708 5370 22764
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5634 22708 5662 22764
rect 5342 21196 5662 22708
rect 5342 21140 5370 21196
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5634 21140 5662 21196
rect 5342 19628 5662 21140
rect 5342 19572 5370 19628
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5634 19572 5662 19628
rect 5342 18060 5662 19572
rect 5342 18004 5370 18060
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5634 18004 5662 18060
rect 5342 16492 5662 18004
rect 5342 16436 5370 16492
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5634 16436 5662 16492
rect 5342 14924 5662 16436
rect 5342 14868 5370 14924
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5634 14868 5662 14924
rect 5342 13356 5662 14868
rect 5342 13300 5370 13356
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5634 13300 5662 13356
rect 5342 11788 5662 13300
rect 4732 11732 4788 11742
rect 3276 10948 3332 10958
rect 3276 9828 3332 10892
rect 3276 9762 3332 9772
rect 4732 10500 4788 11676
rect 4172 8820 4228 8830
rect 3948 7700 4004 7710
rect 3948 6356 4004 7644
rect 4172 7252 4228 8764
rect 4172 7186 4228 7196
rect 3948 6290 4004 6300
rect 4732 4564 4788 10444
rect 5342 11732 5370 11788
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5634 11732 5662 11788
rect 5342 10220 5662 11732
rect 9500 31388 9820 32204
rect 9500 31332 9528 31388
rect 9584 31332 9632 31388
rect 9688 31332 9736 31388
rect 9792 31332 9820 31388
rect 9500 29820 9820 31332
rect 9500 29764 9528 29820
rect 9584 29764 9632 29820
rect 9688 29764 9736 29820
rect 9792 29764 9820 29820
rect 9500 28252 9820 29764
rect 9500 28196 9528 28252
rect 9584 28196 9632 28252
rect 9688 28196 9736 28252
rect 9792 28196 9820 28252
rect 9500 26684 9820 28196
rect 9500 26628 9528 26684
rect 9584 26628 9632 26684
rect 9688 26628 9736 26684
rect 9792 26628 9820 26684
rect 9500 25116 9820 26628
rect 13658 32172 13978 32204
rect 13658 32116 13686 32172
rect 13742 32116 13790 32172
rect 13846 32116 13894 32172
rect 13950 32116 13978 32172
rect 13658 30604 13978 32116
rect 13658 30548 13686 30604
rect 13742 30548 13790 30604
rect 13846 30548 13894 30604
rect 13950 30548 13978 30604
rect 13658 29036 13978 30548
rect 13658 28980 13686 29036
rect 13742 28980 13790 29036
rect 13846 28980 13894 29036
rect 13950 28980 13978 29036
rect 13658 27468 13978 28980
rect 13658 27412 13686 27468
rect 13742 27412 13790 27468
rect 13846 27412 13894 27468
rect 13950 27412 13978 27468
rect 13658 25900 13978 27412
rect 13658 25844 13686 25900
rect 13742 25844 13790 25900
rect 13846 25844 13894 25900
rect 13950 25844 13978 25900
rect 9500 25060 9528 25116
rect 9584 25060 9632 25116
rect 9688 25060 9736 25116
rect 9792 25060 9820 25116
rect 9500 23548 9820 25060
rect 12348 25508 12404 25518
rect 12236 24724 12292 24734
rect 9500 23492 9528 23548
rect 9584 23492 9632 23548
rect 9688 23492 9736 23548
rect 9792 23492 9820 23548
rect 11900 24052 11956 24062
rect 11900 23604 11956 23996
rect 12236 23828 12292 24668
rect 12236 23762 12292 23772
rect 11900 23538 11956 23548
rect 12348 23604 12404 25452
rect 12460 25396 12516 25406
rect 12460 24724 12516 25340
rect 12460 24658 12516 24668
rect 13658 24332 13978 25844
rect 17816 31388 18136 32204
rect 17816 31332 17844 31388
rect 17900 31332 17948 31388
rect 18004 31332 18052 31388
rect 18108 31332 18136 31388
rect 17816 29820 18136 31332
rect 17816 29764 17844 29820
rect 17900 29764 17948 29820
rect 18004 29764 18052 29820
rect 18108 29764 18136 29820
rect 17816 28252 18136 29764
rect 17816 28196 17844 28252
rect 17900 28196 17948 28252
rect 18004 28196 18052 28252
rect 18108 28196 18136 28252
rect 17816 26684 18136 28196
rect 17816 26628 17844 26684
rect 17900 26628 17948 26684
rect 18004 26628 18052 26684
rect 18108 26628 18136 26684
rect 17816 25116 18136 26628
rect 17816 25060 17844 25116
rect 17900 25060 17948 25116
rect 18004 25060 18052 25116
rect 18108 25060 18136 25116
rect 13658 24276 13686 24332
rect 13742 24276 13790 24332
rect 13846 24276 13894 24332
rect 13950 24276 13978 24332
rect 13468 24052 13524 24062
rect 12348 23538 12404 23548
rect 12572 23828 12628 23838
rect 12572 23604 12628 23772
rect 12572 23538 12628 23548
rect 13468 23604 13524 23996
rect 13468 23538 13524 23548
rect 9500 21980 9820 23492
rect 11228 23492 11284 23502
rect 11228 22820 11284 23436
rect 11228 22754 11284 22764
rect 13658 22764 13978 24276
rect 9500 21924 9528 21980
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9792 21924 9820 21980
rect 9500 20412 9820 21924
rect 9500 20356 9528 20412
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9792 20356 9820 20412
rect 9500 18844 9820 20356
rect 9500 18788 9528 18844
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9792 18788 9820 18844
rect 13658 22708 13686 22764
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13950 22708 13978 22764
rect 13658 21196 13978 22708
rect 13658 21140 13686 21196
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13950 21140 13978 21196
rect 13658 19628 13978 21140
rect 14588 24724 14644 24734
rect 14588 19908 14644 24668
rect 14588 19842 14644 19852
rect 17816 23548 18136 25060
rect 17816 23492 17844 23548
rect 17900 23492 17948 23548
rect 18004 23492 18052 23548
rect 18108 23492 18136 23548
rect 17816 21980 18136 23492
rect 17816 21924 17844 21980
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 18108 21924 18136 21980
rect 17816 20412 18136 21924
rect 17816 20356 17844 20412
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 18108 20356 18136 20412
rect 13658 19572 13686 19628
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13950 19572 13978 19628
rect 9500 17276 9820 18788
rect 11116 18788 11172 18798
rect 11116 17780 11172 18732
rect 11116 17714 11172 17724
rect 13658 18060 13978 19572
rect 13658 18004 13686 18060
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13950 18004 13978 18060
rect 9500 17220 9528 17276
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9792 17220 9820 17276
rect 9500 15708 9820 17220
rect 9500 15652 9528 15708
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9792 15652 9820 15708
rect 9500 14140 9820 15652
rect 9500 14084 9528 14140
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9792 14084 9820 14140
rect 9500 12572 9820 14084
rect 9500 12516 9528 12572
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9792 12516 9820 12572
rect 9500 11004 9820 12516
rect 5342 10164 5370 10220
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5634 10164 5662 10220
rect 8876 10948 8932 10958
rect 4956 10052 5012 10062
rect 4956 8260 5012 9996
rect 4956 8194 5012 8204
rect 5342 8652 5662 10164
rect 7420 10164 7476 10174
rect 5342 8596 5370 8652
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5634 8596 5662 8652
rect 5068 7924 5124 7934
rect 5068 7028 5124 7868
rect 5068 6962 5124 6972
rect 5342 7084 5662 8596
rect 6860 8708 6916 8718
rect 6636 8484 6692 8494
rect 5342 7028 5370 7084
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5634 7028 5662 7084
rect 4732 4498 4788 4508
rect 5342 5516 5662 7028
rect 5342 5460 5370 5516
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5634 5460 5662 5516
rect 5342 3948 5662 5460
rect 5740 7140 5796 7150
rect 5740 5460 5796 7084
rect 5740 5394 5796 5404
rect 6636 4900 6692 8428
rect 6636 4834 6692 4844
rect 6860 4228 6916 8652
rect 7196 8596 7252 8606
rect 7196 7924 7252 8540
rect 7196 7858 7252 7868
rect 7420 6468 7476 10108
rect 8876 8708 8932 10892
rect 8876 8642 8932 8652
rect 9500 10948 9528 11004
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9792 10948 9820 11004
rect 9500 9436 9820 10948
rect 13658 16492 13978 18004
rect 17816 18844 18136 20356
rect 17816 18788 17844 18844
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 18108 18788 18136 18844
rect 17052 17780 17108 17790
rect 17052 16884 17108 17724
rect 17052 16818 17108 16828
rect 17816 17276 18136 18788
rect 17816 17220 17844 17276
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 18108 17220 18136 17276
rect 13658 16436 13686 16492
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13950 16436 13978 16492
rect 13658 14924 13978 16436
rect 13658 14868 13686 14924
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13950 14868 13978 14924
rect 13658 13356 13978 14868
rect 13658 13300 13686 13356
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13950 13300 13978 13356
rect 13658 11788 13978 13300
rect 13658 11732 13686 11788
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13950 11732 13978 11788
rect 9500 9380 9528 9436
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9792 9380 9820 9436
rect 9500 7868 9820 9380
rect 9884 10612 9940 10622
rect 9884 8036 9940 10556
rect 10108 10388 10164 10398
rect 9884 7970 9940 7980
rect 9996 9044 10052 9054
rect 9500 7812 9528 7868
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9792 7812 9820 7868
rect 7420 6402 7476 6412
rect 7644 7140 7700 7150
rect 7644 4564 7700 7084
rect 7644 4498 7700 4508
rect 9500 6300 9820 7812
rect 9996 6804 10052 8988
rect 9996 6738 10052 6748
rect 9500 6244 9528 6300
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9792 6244 9820 6300
rect 9500 4732 9820 6244
rect 10108 5460 10164 10332
rect 13658 10220 13978 11732
rect 13658 10164 13686 10220
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13950 10164 13978 10220
rect 10108 5394 10164 5404
rect 10556 9828 10612 9838
rect 10556 5460 10612 9772
rect 13658 8652 13978 10164
rect 13658 8596 13686 8652
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13950 8596 13978 8652
rect 13132 7924 13188 7934
rect 11452 7476 11508 7486
rect 11452 6020 11508 7420
rect 11452 5954 11508 5964
rect 10556 5394 10612 5404
rect 9500 4676 9528 4732
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9792 4676 9820 4732
rect 6860 4162 6916 4172
rect 5342 3892 5370 3948
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5634 3892 5662 3948
rect 5342 3076 5662 3892
rect 9500 3164 9820 4676
rect 9500 3108 9528 3164
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9792 3108 9820 3164
rect 9500 3076 9820 3108
rect 13132 3108 13188 7868
rect 13658 7084 13978 8596
rect 13658 7028 13686 7084
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13950 7028 13978 7084
rect 13658 5516 13978 7028
rect 13658 5460 13686 5516
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13950 5460 13978 5516
rect 13658 3948 13978 5460
rect 13658 3892 13686 3948
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13950 3892 13978 3948
rect 13658 3076 13978 3892
rect 17816 15708 18136 17220
rect 17816 15652 17844 15708
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 18108 15652 18136 15708
rect 17816 14140 18136 15652
rect 17816 14084 17844 14140
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 18108 14084 18136 14140
rect 17816 12572 18136 14084
rect 17816 12516 17844 12572
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 18108 12516 18136 12572
rect 17816 11004 18136 12516
rect 17816 10948 17844 11004
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 18108 10948 18136 11004
rect 17816 9436 18136 10948
rect 17816 9380 17844 9436
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 18108 9380 18136 9436
rect 17816 7868 18136 9380
rect 17816 7812 17844 7868
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 18108 7812 18136 7868
rect 17816 6300 18136 7812
rect 17816 6244 17844 6300
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 18108 6244 18136 6300
rect 17816 4732 18136 6244
rect 17816 4676 17844 4732
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 18108 4676 18136 4732
rect 17816 3164 18136 4676
rect 17816 3108 17844 3164
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 18108 3108 18136 3164
rect 17816 3076 18136 3108
rect 21974 32172 22294 32204
rect 21974 32116 22002 32172
rect 22058 32116 22106 32172
rect 22162 32116 22210 32172
rect 22266 32116 22294 32172
rect 21974 30604 22294 32116
rect 21974 30548 22002 30604
rect 22058 30548 22106 30604
rect 22162 30548 22210 30604
rect 22266 30548 22294 30604
rect 21974 29036 22294 30548
rect 21974 28980 22002 29036
rect 22058 28980 22106 29036
rect 22162 28980 22210 29036
rect 22266 28980 22294 29036
rect 21974 27468 22294 28980
rect 21974 27412 22002 27468
rect 22058 27412 22106 27468
rect 22162 27412 22210 27468
rect 22266 27412 22294 27468
rect 21974 25900 22294 27412
rect 21974 25844 22002 25900
rect 22058 25844 22106 25900
rect 22162 25844 22210 25900
rect 22266 25844 22294 25900
rect 21974 24332 22294 25844
rect 21974 24276 22002 24332
rect 22058 24276 22106 24332
rect 22162 24276 22210 24332
rect 22266 24276 22294 24332
rect 21974 22764 22294 24276
rect 21974 22708 22002 22764
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22266 22708 22294 22764
rect 21974 21196 22294 22708
rect 21974 21140 22002 21196
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22266 21140 22294 21196
rect 21974 19628 22294 21140
rect 21974 19572 22002 19628
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22266 19572 22294 19628
rect 21974 18060 22294 19572
rect 21974 18004 22002 18060
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22266 18004 22294 18060
rect 21974 16492 22294 18004
rect 21974 16436 22002 16492
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22266 16436 22294 16492
rect 21974 14924 22294 16436
rect 21974 14868 22002 14924
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22266 14868 22294 14924
rect 21974 13356 22294 14868
rect 21974 13300 22002 13356
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22266 13300 22294 13356
rect 21974 11788 22294 13300
rect 21974 11732 22002 11788
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22266 11732 22294 11788
rect 21974 10220 22294 11732
rect 21974 10164 22002 10220
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22266 10164 22294 10220
rect 21974 8652 22294 10164
rect 21974 8596 22002 8652
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22266 8596 22294 8652
rect 21974 7084 22294 8596
rect 21974 7028 22002 7084
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22266 7028 22294 7084
rect 21974 5516 22294 7028
rect 21974 5460 22002 5516
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22266 5460 22294 5516
rect 21974 3948 22294 5460
rect 21974 3892 22002 3948
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22266 3892 22294 3948
rect 21974 3076 22294 3892
rect 26132 31388 26452 32204
rect 26132 31332 26160 31388
rect 26216 31332 26264 31388
rect 26320 31332 26368 31388
rect 26424 31332 26452 31388
rect 26132 29820 26452 31332
rect 26132 29764 26160 29820
rect 26216 29764 26264 29820
rect 26320 29764 26368 29820
rect 26424 29764 26452 29820
rect 26132 28252 26452 29764
rect 26132 28196 26160 28252
rect 26216 28196 26264 28252
rect 26320 28196 26368 28252
rect 26424 28196 26452 28252
rect 26132 26684 26452 28196
rect 26132 26628 26160 26684
rect 26216 26628 26264 26684
rect 26320 26628 26368 26684
rect 26424 26628 26452 26684
rect 26132 25116 26452 26628
rect 26132 25060 26160 25116
rect 26216 25060 26264 25116
rect 26320 25060 26368 25116
rect 26424 25060 26452 25116
rect 26132 23548 26452 25060
rect 26132 23492 26160 23548
rect 26216 23492 26264 23548
rect 26320 23492 26368 23548
rect 26424 23492 26452 23548
rect 26132 21980 26452 23492
rect 26132 21924 26160 21980
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26424 21924 26452 21980
rect 26132 20412 26452 21924
rect 26132 20356 26160 20412
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26424 20356 26452 20412
rect 26132 18844 26452 20356
rect 26132 18788 26160 18844
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26424 18788 26452 18844
rect 26132 17276 26452 18788
rect 26132 17220 26160 17276
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26424 17220 26452 17276
rect 26132 15708 26452 17220
rect 26132 15652 26160 15708
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26424 15652 26452 15708
rect 26132 14140 26452 15652
rect 26132 14084 26160 14140
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26424 14084 26452 14140
rect 26132 12572 26452 14084
rect 26132 12516 26160 12572
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26424 12516 26452 12572
rect 26132 11004 26452 12516
rect 26132 10948 26160 11004
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26424 10948 26452 11004
rect 26132 9436 26452 10948
rect 26132 9380 26160 9436
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 26424 9380 26452 9436
rect 26132 7868 26452 9380
rect 26132 7812 26160 7868
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26424 7812 26452 7868
rect 26132 6300 26452 7812
rect 26132 6244 26160 6300
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26424 6244 26452 6300
rect 26132 4732 26452 6244
rect 26132 4676 26160 4732
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26424 4676 26452 4732
rect 26132 3164 26452 4676
rect 26132 3108 26160 3164
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26424 3108 26452 3164
rect 26132 3076 26452 3108
rect 30290 32172 30610 32204
rect 30290 32116 30318 32172
rect 30374 32116 30422 32172
rect 30478 32116 30526 32172
rect 30582 32116 30610 32172
rect 30290 30604 30610 32116
rect 30290 30548 30318 30604
rect 30374 30548 30422 30604
rect 30478 30548 30526 30604
rect 30582 30548 30610 30604
rect 30290 29036 30610 30548
rect 30290 28980 30318 29036
rect 30374 28980 30422 29036
rect 30478 28980 30526 29036
rect 30582 28980 30610 29036
rect 30290 27468 30610 28980
rect 30290 27412 30318 27468
rect 30374 27412 30422 27468
rect 30478 27412 30526 27468
rect 30582 27412 30610 27468
rect 30290 25900 30610 27412
rect 30290 25844 30318 25900
rect 30374 25844 30422 25900
rect 30478 25844 30526 25900
rect 30582 25844 30610 25900
rect 30290 24332 30610 25844
rect 30290 24276 30318 24332
rect 30374 24276 30422 24332
rect 30478 24276 30526 24332
rect 30582 24276 30610 24332
rect 30290 22764 30610 24276
rect 30290 22708 30318 22764
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30582 22708 30610 22764
rect 30290 21196 30610 22708
rect 30290 21140 30318 21196
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30582 21140 30610 21196
rect 30290 19628 30610 21140
rect 30290 19572 30318 19628
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30582 19572 30610 19628
rect 30290 18060 30610 19572
rect 30290 18004 30318 18060
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30582 18004 30610 18060
rect 30290 16492 30610 18004
rect 30290 16436 30318 16492
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30582 16436 30610 16492
rect 30290 14924 30610 16436
rect 30290 14868 30318 14924
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30582 14868 30610 14924
rect 30290 13356 30610 14868
rect 30290 13300 30318 13356
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30582 13300 30610 13356
rect 30290 11788 30610 13300
rect 30290 11732 30318 11788
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30582 11732 30610 11788
rect 30290 10220 30610 11732
rect 30290 10164 30318 10220
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30582 10164 30610 10220
rect 30290 8652 30610 10164
rect 30290 8596 30318 8652
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30582 8596 30610 8652
rect 30290 7084 30610 8596
rect 30290 7028 30318 7084
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30582 7028 30610 7084
rect 30290 5516 30610 7028
rect 30290 5460 30318 5516
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30582 5460 30610 5516
rect 30290 3948 30610 5460
rect 30290 3892 30318 3948
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30582 3892 30610 3948
rect 30290 3076 30610 3892
rect 34448 31388 34768 32204
rect 34448 31332 34476 31388
rect 34532 31332 34580 31388
rect 34636 31332 34684 31388
rect 34740 31332 34768 31388
rect 34448 29820 34768 31332
rect 34448 29764 34476 29820
rect 34532 29764 34580 29820
rect 34636 29764 34684 29820
rect 34740 29764 34768 29820
rect 34448 28252 34768 29764
rect 34448 28196 34476 28252
rect 34532 28196 34580 28252
rect 34636 28196 34684 28252
rect 34740 28196 34768 28252
rect 34448 26684 34768 28196
rect 34448 26628 34476 26684
rect 34532 26628 34580 26684
rect 34636 26628 34684 26684
rect 34740 26628 34768 26684
rect 34448 25116 34768 26628
rect 34448 25060 34476 25116
rect 34532 25060 34580 25116
rect 34636 25060 34684 25116
rect 34740 25060 34768 25116
rect 34448 23548 34768 25060
rect 34448 23492 34476 23548
rect 34532 23492 34580 23548
rect 34636 23492 34684 23548
rect 34740 23492 34768 23548
rect 34448 21980 34768 23492
rect 34448 21924 34476 21980
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34740 21924 34768 21980
rect 34448 20412 34768 21924
rect 34448 20356 34476 20412
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34740 20356 34768 20412
rect 34448 18844 34768 20356
rect 34448 18788 34476 18844
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34740 18788 34768 18844
rect 34448 17276 34768 18788
rect 34448 17220 34476 17276
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34740 17220 34768 17276
rect 34448 15708 34768 17220
rect 34448 15652 34476 15708
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34740 15652 34768 15708
rect 34448 14140 34768 15652
rect 34448 14084 34476 14140
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34740 14084 34768 14140
rect 34448 12572 34768 14084
rect 34448 12516 34476 12572
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34740 12516 34768 12572
rect 34448 11004 34768 12516
rect 34448 10948 34476 11004
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34740 10948 34768 11004
rect 34448 9436 34768 10948
rect 34448 9380 34476 9436
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34740 9380 34768 9436
rect 34448 7868 34768 9380
rect 34448 7812 34476 7868
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34740 7812 34768 7868
rect 34448 6300 34768 7812
rect 34448 6244 34476 6300
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34740 6244 34768 6300
rect 34448 4732 34768 6244
rect 34448 4676 34476 4732
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34740 4676 34768 4732
rect 34448 3164 34768 4676
rect 34448 3108 34476 3164
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34740 3108 34768 3164
rect 34448 3076 34768 3108
rect 13132 3042 13188 3052
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _428_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12432 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _429_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _430_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _431_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18816 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _432_
timestamp 1698431365
transform 1 0 16576 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_4  _433_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24192 0 1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and4_4  _434_
timestamp 1698431365
transform -1 0 24864 0 -1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _435_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24192 0 1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and3_4  _436_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24976 0 1 26656
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _437_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _438_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17248 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _439_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23632 0 -1 25088
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _440_
timestamp 1698431365
transform 1 0 4816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _441_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6944 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _442_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5264 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _443_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _444_
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _445_
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _446_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _447_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _448_
timestamp 1698431365
transform -1 0 20720 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _449_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22400 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _450_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19712 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _451_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18032 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _452_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _453_
timestamp 1698431365
transform -1 0 18032 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _454_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _455_
timestamp 1698431365
transform -1 0 12320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _456_
timestamp 1698431365
transform -1 0 18144 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_4  _457_
timestamp 1698431365
transform -1 0 17024 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _458_
timestamp 1698431365
transform -1 0 16912 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _459_
timestamp 1698431365
transform -1 0 12096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _460_
timestamp 1698431365
transform 1 0 10976 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _461_
timestamp 1698431365
transform 1 0 10192 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _462_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7728 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _463_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8512 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _464_
timestamp 1698431365
transform -1 0 13104 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _465_
timestamp 1698431365
transform -1 0 14000 0 -1 7840
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _466_
timestamp 1698431365
transform 1 0 10416 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _467_
timestamp 1698431365
transform -1 0 11200 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _468_
timestamp 1698431365
transform 1 0 11088 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _469_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14112 0 -1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _470_
timestamp 1698431365
transform 1 0 18032 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _471_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18816 0 1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _472_
timestamp 1698431365
transform 1 0 11872 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _473_
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _474_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14112 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _475_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15120 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _476_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14784 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _477_
timestamp 1698431365
transform -1 0 8624 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _478_
timestamp 1698431365
transform 1 0 7168 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _479_
timestamp 1698431365
transform 1 0 18592 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _480_
timestamp 1698431365
transform 1 0 15008 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _481_
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _482_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11872 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _483_
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _484_
timestamp 1698431365
transform -1 0 11088 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _485_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4816 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _486_
timestamp 1698431365
transform -1 0 7616 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _487_
timestamp 1698431365
transform 1 0 7616 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _488_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11760 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _489_
timestamp 1698431365
transform -1 0 18592 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _490_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _491_
timestamp 1698431365
transform -1 0 11312 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _492_
timestamp 1698431365
transform -1 0 3696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _493_
timestamp 1698431365
transform -1 0 2800 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _494_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15680 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _495_
timestamp 1698431365
transform -1 0 7168 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _496_
timestamp 1698431365
transform -1 0 12320 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _497_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7056 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _498_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6608 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _499_
timestamp 1698431365
transform -1 0 5152 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _500_
timestamp 1698431365
transform 1 0 9408 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _501_
timestamp 1698431365
transform 1 0 6272 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _502_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _503_
timestamp 1698431365
transform 1 0 9856 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _504_
timestamp 1698431365
transform 1 0 7616 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _505_
timestamp 1698431365
transform 1 0 2800 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _506_
timestamp 1698431365
transform 1 0 3584 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _507_
timestamp 1698431365
transform -1 0 12992 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _508_
timestamp 1698431365
transform 1 0 8064 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _509_
timestamp 1698431365
transform -1 0 8288 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _510_
timestamp 1698431365
transform 1 0 13776 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _511_
timestamp 1698431365
transform 1 0 5152 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _512_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6832 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _513_
timestamp 1698431365
transform -1 0 10976 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _514_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7392 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _515_
timestamp 1698431365
transform 1 0 7280 0 -1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _516_
timestamp 1698431365
transform 1 0 8288 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _517_
timestamp 1698431365
transform 1 0 2688 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _518_
timestamp 1698431365
transform -1 0 10976 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _519_
timestamp 1698431365
transform 1 0 10192 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _520_
timestamp 1698431365
transform -1 0 8512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _521_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3248 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _522_
timestamp 1698431365
transform 1 0 10640 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _523_
timestamp 1698431365
transform 1 0 6608 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _524_
timestamp 1698431365
transform -1 0 12096 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _525_
timestamp 1698431365
transform -1 0 9968 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _526_
timestamp 1698431365
transform -1 0 6832 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _527_
timestamp 1698431365
transform -1 0 10304 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _528_
timestamp 1698431365
transform -1 0 10080 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _529_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _530_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8624 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _531_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _532_
timestamp 1698431365
transform 1 0 8288 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _533_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10976 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _534_
timestamp 1698431365
transform 1 0 13328 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _535_
timestamp 1698431365
transform -1 0 5936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _536_
timestamp 1698431365
transform -1 0 6944 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _537_
timestamp 1698431365
transform -1 0 5264 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _538_
timestamp 1698431365
transform 1 0 2352 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _539_
timestamp 1698431365
transform -1 0 3024 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _540_
timestamp 1698431365
transform 1 0 4704 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _541_
timestamp 1698431365
transform 1 0 11312 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _542_
timestamp 1698431365
transform -1 0 11424 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _543_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7616 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _544_
timestamp 1698431365
transform 1 0 7504 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _545_
timestamp 1698431365
transform -1 0 7840 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _546_
timestamp 1698431365
transform 1 0 6272 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _547_
timestamp 1698431365
transform 1 0 7504 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _548_
timestamp 1698431365
transform 1 0 4144 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _549_
timestamp 1698431365
transform 1 0 6496 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _550_
timestamp 1698431365
transform 1 0 2016 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _551_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3584 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _552_
timestamp 1698431365
transform -1 0 6720 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _553_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _554_
timestamp 1698431365
transform -1 0 10416 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _555_
timestamp 1698431365
transform 1 0 3360 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _556_
timestamp 1698431365
transform -1 0 3360 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _557_
timestamp 1698431365
transform 1 0 2688 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _558_
timestamp 1698431365
transform -1 0 5264 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _559_
timestamp 1698431365
transform -1 0 3024 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _560_
timestamp 1698431365
transform -1 0 5264 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _561_
timestamp 1698431365
transform 1 0 3024 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _562_
timestamp 1698431365
transform 1 0 3472 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _563_
timestamp 1698431365
transform 1 0 2688 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _564_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3024 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _565_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1904 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _566_
timestamp 1698431365
transform -1 0 6384 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _567_
timestamp 1698431365
transform 1 0 3360 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _568_
timestamp 1698431365
transform -1 0 5152 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _569_
timestamp 1698431365
transform -1 0 7728 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _570_
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _571_
timestamp 1698431365
transform 1 0 5824 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _572_
timestamp 1698431365
transform 1 0 2912 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _573_
timestamp 1698431365
transform -1 0 5264 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _574_
timestamp 1698431365
transform 1 0 4032 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _575_
timestamp 1698431365
transform 1 0 3472 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _576_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _577_
timestamp 1698431365
transform 1 0 6720 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _578_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _579_
timestamp 1698431365
transform -1 0 7056 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _580_
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _581_
timestamp 1698431365
transform -1 0 32704 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _582_
timestamp 1698431365
transform 1 0 13664 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _583_
timestamp 1698431365
transform -1 0 27664 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _584_
timestamp 1698431365
transform -1 0 23072 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _585_
timestamp 1698431365
transform -1 0 33824 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _586_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22064 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _587_
timestamp 1698431365
transform -1 0 30800 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _588_
timestamp 1698431365
transform -1 0 30576 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _589_
timestamp 1698431365
transform -1 0 30352 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _590_
timestamp 1698431365
transform 1 0 26768 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _591_
timestamp 1698431365
transform -1 0 27888 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _592_
timestamp 1698431365
transform 1 0 27664 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _593_
timestamp 1698431365
transform 1 0 30576 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _594_
timestamp 1698431365
transform -1 0 31920 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _595_
timestamp 1698431365
transform -1 0 26432 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _596_
timestamp 1698431365
transform 1 0 27776 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _597_
timestamp 1698431365
transform -1 0 28560 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _598_
timestamp 1698431365
transform 1 0 23072 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _599_
timestamp 1698431365
transform 1 0 23408 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _600_
timestamp 1698431365
transform 1 0 25200 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _601_
timestamp 1698431365
transform -1 0 26768 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _602_
timestamp 1698431365
transform -1 0 22288 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _603_
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _604_
timestamp 1698431365
transform 1 0 19376 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _605_
timestamp 1698431365
transform -1 0 22512 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _606_
timestamp 1698431365
transform -1 0 22064 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _607_
timestamp 1698431365
transform -1 0 28224 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _608_
timestamp 1698431365
transform -1 0 23520 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _609_
timestamp 1698431365
transform 1 0 23184 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _610_
timestamp 1698431365
transform -1 0 22288 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _611_
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _612_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21840 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _613_
timestamp 1698431365
transform 1 0 26096 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _614_
timestamp 1698431365
transform -1 0 24416 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _615_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23408 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _616_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _617_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _618_
timestamp 1698431365
transform 1 0 26656 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _619_
timestamp 1698431365
transform 1 0 27216 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _620_
timestamp 1698431365
transform 1 0 27328 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _621_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _622_
timestamp 1698431365
transform 1 0 26432 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _623_
timestamp 1698431365
transform 1 0 28000 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _624_
timestamp 1698431365
transform 1 0 28560 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _625_
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _626_
timestamp 1698431365
transform -1 0 30352 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _627_
timestamp 1698431365
transform -1 0 29904 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _628_
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _629_
timestamp 1698431365
transform 1 0 29904 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _630_
timestamp 1698431365
transform -1 0 31360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _631_
timestamp 1698431365
transform 1 0 30240 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _632_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _633_
timestamp 1698431365
transform 1 0 30016 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _634_
timestamp 1698431365
transform 1 0 31360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _635_
timestamp 1698431365
transform 1 0 29120 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _636_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _637_
timestamp 1698431365
transform -1 0 32368 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _638_
timestamp 1698431365
transform 1 0 31696 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _639_
timestamp 1698431365
transform -1 0 31472 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _640_
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _641_
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _642_
timestamp 1698431365
transform -1 0 29904 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _643_
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _644_
timestamp 1698431365
transform 1 0 30240 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _645_
timestamp 1698431365
transform -1 0 31136 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _646_
timestamp 1698431365
transform 1 0 31248 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _647_
timestamp 1698431365
transform -1 0 31584 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _648_
timestamp 1698431365
transform 1 0 31584 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _649_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _650_
timestamp 1698431365
transform -1 0 33824 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _651_
timestamp 1698431365
transform -1 0 30800 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _652_
timestamp 1698431365
transform 1 0 32480 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _653_
timestamp 1698431365
transform 1 0 31024 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _654_
timestamp 1698431365
transform -1 0 32368 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _655_
timestamp 1698431365
transform 1 0 31920 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _656_
timestamp 1698431365
transform -1 0 28784 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _657_
timestamp 1698431365
transform 1 0 28336 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _658_
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _659_
timestamp 1698431365
transform -1 0 27328 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _660_
timestamp 1698431365
transform -1 0 26208 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _661_
timestamp 1698431365
transform -1 0 26768 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _662_
timestamp 1698431365
transform 1 0 27104 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _663_
timestamp 1698431365
transform -1 0 27664 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _664_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _665_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _666_
timestamp 1698431365
transform -1 0 27664 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _667_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _668_
timestamp 1698431365
transform -1 0 29904 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _669_
timestamp 1698431365
transform -1 0 27776 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _670_
timestamp 1698431365
transform 1 0 25648 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _671_
timestamp 1698431365
transform -1 0 26544 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _672_
timestamp 1698431365
transform 1 0 22400 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _673_
timestamp 1698431365
transform -1 0 17920 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _674_
timestamp 1698431365
transform 1 0 17248 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _675_
timestamp 1698431365
transform 1 0 19376 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _676_
timestamp 1698431365
transform 1 0 20048 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _677_
timestamp 1698431365
transform -1 0 18816 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _678_
timestamp 1698431365
transform 1 0 20496 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _679_
timestamp 1698431365
transform -1 0 22960 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _680_
timestamp 1698431365
transform 1 0 24192 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _681_
timestamp 1698431365
transform -1 0 16912 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _682_
timestamp 1698431365
transform -1 0 15904 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _683_
timestamp 1698431365
transform 1 0 11088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _684_
timestamp 1698431365
transform -1 0 13664 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _685_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _686_
timestamp 1698431365
transform -1 0 14000 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _687_
timestamp 1698431365
transform 1 0 13888 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _688_
timestamp 1698431365
transform 1 0 15680 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _689_
timestamp 1698431365
transform -1 0 15904 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _690_
timestamp 1698431365
transform 1 0 17920 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _691_
timestamp 1698431365
transform -1 0 18480 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _692_
timestamp 1698431365
transform -1 0 19376 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _693_
timestamp 1698431365
transform 1 0 19152 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _694_
timestamp 1698431365
transform -1 0 19376 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _695_
timestamp 1698431365
transform 1 0 14560 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _696_
timestamp 1698431365
transform -1 0 15344 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _697_
timestamp 1698431365
transform -1 0 12880 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _698_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _699_
timestamp 1698431365
transform 1 0 6720 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _700_
timestamp 1698431365
transform 1 0 7056 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _701_
timestamp 1698431365
transform 1 0 7392 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _702_
timestamp 1698431365
transform 1 0 6608 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _703_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _704_
timestamp 1698431365
transform -1 0 11424 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _705_
timestamp 1698431365
transform 1 0 6160 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _706_
timestamp 1698431365
transform 1 0 7504 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _707_
timestamp 1698431365
transform 1 0 8512 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _708_
timestamp 1698431365
transform 1 0 10416 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _709_
timestamp 1698431365
transform 1 0 11984 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _710_
timestamp 1698431365
transform -1 0 18816 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _711_
timestamp 1698431365
transform -1 0 18032 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _712_
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _713_
timestamp 1698431365
transform 1 0 11984 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _714_
timestamp 1698431365
transform -1 0 14672 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _715_
timestamp 1698431365
transform 1 0 9408 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _716_
timestamp 1698431365
transform -1 0 9184 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _717_
timestamp 1698431365
transform 1 0 6048 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _718_
timestamp 1698431365
transform 1 0 7952 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _719_
timestamp 1698431365
transform 1 0 8624 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _720_
timestamp 1698431365
transform 1 0 9968 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _721_
timestamp 1698431365
transform 1 0 11200 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _722_
timestamp 1698431365
transform 1 0 11872 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _723_
timestamp 1698431365
transform -1 0 11984 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _724_
timestamp 1698431365
transform -1 0 18480 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _725_
timestamp 1698431365
transform 1 0 10864 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _726_
timestamp 1698431365
transform -1 0 10192 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _727_
timestamp 1698431365
transform 1 0 11088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _728_
timestamp 1698431365
transform 1 0 7616 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _729_
timestamp 1698431365
transform -1 0 12992 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _730_
timestamp 1698431365
transform -1 0 12320 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _731_
timestamp 1698431365
transform 1 0 9744 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _732_
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _733_
timestamp 1698431365
transform 1 0 10752 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _734_
timestamp 1698431365
transform -1 0 9184 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _735_
timestamp 1698431365
transform 1 0 7056 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _736_
timestamp 1698431365
transform 1 0 12320 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _737_
timestamp 1698431365
transform 1 0 12544 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _738_
timestamp 1698431365
transform 1 0 14000 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _739_
timestamp 1698431365
transform 1 0 15120 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _740_
timestamp 1698431365
transform -1 0 14560 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _741_
timestamp 1698431365
transform -1 0 13104 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _742_
timestamp 1698431365
transform -1 0 9072 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _743_
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _744_
timestamp 1698431365
transform 1 0 11984 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _745_
timestamp 1698431365
transform 1 0 10080 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _746_
timestamp 1698431365
transform -1 0 12544 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _747_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _748_
timestamp 1698431365
transform -1 0 15120 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _749_
timestamp 1698431365
transform -1 0 14000 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _750_
timestamp 1698431365
transform -1 0 8624 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _751_
timestamp 1698431365
transform -1 0 9408 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _752_
timestamp 1698431365
transform 1 0 6832 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _753_
timestamp 1698431365
transform -1 0 10192 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _754_
timestamp 1698431365
transform -1 0 9296 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _755_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _756_
timestamp 1698431365
transform -1 0 15456 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _757_
timestamp 1698431365
transform -1 0 18704 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _758_
timestamp 1698431365
transform 1 0 16016 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _759_
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _760_
timestamp 1698431365
transform 1 0 11312 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _761_
timestamp 1698431365
transform -1 0 11088 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _762_
timestamp 1698431365
transform 1 0 10080 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _763_
timestamp 1698431365
transform -1 0 12768 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _764_
timestamp 1698431365
transform 1 0 16016 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _765_
timestamp 1698431365
transform 1 0 14224 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _766_
timestamp 1698431365
transform -1 0 18816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _767_
timestamp 1698431365
transform -1 0 23744 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _768_
timestamp 1698431365
transform 1 0 18592 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _769_
timestamp 1698431365
transform 1 0 17696 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _770_
timestamp 1698431365
transform -1 0 24080 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _771_
timestamp 1698431365
transform 1 0 18704 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _772_
timestamp 1698431365
transform 1 0 19152 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _773_
timestamp 1698431365
transform -1 0 19376 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _774_
timestamp 1698431365
transform 1 0 19376 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _775_
timestamp 1698431365
transform 1 0 20384 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _776_
timestamp 1698431365
transform 1 0 21728 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _777_
timestamp 1698431365
transform -1 0 22848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _778_
timestamp 1698431365
transform 1 0 20160 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _779_
timestamp 1698431365
transform -1 0 22176 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _780_
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _781_
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _782_
timestamp 1698431365
transform 1 0 16352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _783_
timestamp 1698431365
transform 1 0 26880 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _784_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _785_
timestamp 1698431365
transform -1 0 26880 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _786_
timestamp 1698431365
transform 1 0 24192 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _787_
timestamp 1698431365
transform 1 0 27776 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _788_
timestamp 1698431365
transform -1 0 27776 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _789_
timestamp 1698431365
transform 1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _790_
timestamp 1698431365
transform -1 0 25984 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _791_
timestamp 1698431365
transform -1 0 27104 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _792_
timestamp 1698431365
transform -1 0 28112 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _793_
timestamp 1698431365
transform 1 0 25424 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _794_
timestamp 1698431365
transform 1 0 26880 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _795_
timestamp 1698431365
transform -1 0 25760 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _796_
timestamp 1698431365
transform -1 0 27776 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _797_
timestamp 1698431365
transform -1 0 26432 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _798_
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _799_
timestamp 1698431365
transform -1 0 19712 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _800_
timestamp 1698431365
transform 1 0 19712 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _801_
timestamp 1698431365
transform -1 0 20720 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _802_
timestamp 1698431365
transform -1 0 18704 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _803_
timestamp 1698431365
transform -1 0 17920 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _804_
timestamp 1698431365
transform 1 0 15680 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _805_
timestamp 1698431365
transform 1 0 15568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _806_
timestamp 1698431365
transform -1 0 18032 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _807_
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _808_
timestamp 1698431365
transform 1 0 15792 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _809_
timestamp 1698431365
transform 1 0 14784 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _810_
timestamp 1698431365
transform -1 0 16128 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _811_
timestamp 1698431365
transform -1 0 15568 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _812_
timestamp 1698431365
transform -1 0 14560 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _813_
timestamp 1698431365
transform -1 0 12544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _814_
timestamp 1698431365
transform 1 0 14672 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _815_
timestamp 1698431365
transform 1 0 15344 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _816_
timestamp 1698431365
transform -1 0 15344 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _817_
timestamp 1698431365
transform -1 0 14672 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _818_
timestamp 1698431365
transform -1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _819_
timestamp 1698431365
transform -1 0 17024 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _820_
timestamp 1698431365
transform -1 0 19488 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _821_
timestamp 1698431365
transform 1 0 16464 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _822_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _823_
timestamp 1698431365
transform 1 0 18816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _824_
timestamp 1698431365
transform -1 0 23184 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _825_
timestamp 1698431365
transform -1 0 23184 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _826_
timestamp 1698431365
transform 1 0 21504 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _827_
timestamp 1698431365
transform 1 0 19936 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _828_
timestamp 1698431365
transform 1 0 21392 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _829_
timestamp 1698431365
transform -1 0 20272 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _830_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _831_
timestamp 1698431365
transform -1 0 22736 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _832_
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _833_
timestamp 1698431365
transform -1 0 16240 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _834_
timestamp 1698431365
transform 1 0 18256 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _835_
timestamp 1698431365
transform 1 0 19600 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _836_
timestamp 1698431365
transform -1 0 3472 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _837_
timestamp 1698431365
transform -1 0 18144 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _838_
timestamp 1698431365
transform -1 0 4592 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _839_
timestamp 1698431365
transform -1 0 2800 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _840_
timestamp 1698431365
transform -1 0 4144 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _841_
timestamp 1698431365
transform 1 0 4144 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _842_
timestamp 1698431365
transform 1 0 4816 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _843_
timestamp 1698431365
transform 1 0 4144 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _844_
timestamp 1698431365
transform 1 0 3248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _845_
timestamp 1698431365
transform -1 0 6384 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _846_
timestamp 1698431365
transform 1 0 4816 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _847_
timestamp 1698431365
transform -1 0 5264 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _848_
timestamp 1698431365
transform 1 0 5712 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _849_
timestamp 1698431365
transform 1 0 6496 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _850_
timestamp 1698431365
transform -1 0 5488 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _851_
timestamp 1698431365
transform 1 0 5600 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _852_
timestamp 1698431365
transform -1 0 5264 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _853_
timestamp 1698431365
transform -1 0 3808 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _854_
timestamp 1698431365
transform -1 0 5376 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _855_
timestamp 1698431365
transform -1 0 4816 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _856_
timestamp 1698431365
transform -1 0 3136 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _857_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12096 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _858_
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _859_
timestamp 1698431365
transform 1 0 3024 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _860_
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _861_
timestamp 1698431365
transform 1 0 2016 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _862_
timestamp 1698431365
transform 1 0 5488 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _863_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _864_
timestamp 1698431365
transform 1 0 18592 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _865_
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _866_
timestamp 1698431365
transform 1 0 19376 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _867_
timestamp 1698431365
transform 1 0 22848 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _868_
timestamp 1698431365
transform -1 0 27216 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _869_
timestamp 1698431365
transform -1 0 28896 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _870_
timestamp 1698431365
transform -1 0 32144 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _871_
timestamp 1698431365
transform 1 0 30912 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _872_
timestamp 1698431365
transform 1 0 31136 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _873_
timestamp 1698431365
transform 1 0 31136 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _874_
timestamp 1698431365
transform -1 0 34384 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _875_
timestamp 1698431365
transform 1 0 26880 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _876_
timestamp 1698431365
transform -1 0 34384 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _877_
timestamp 1698431365
transform -1 0 34384 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _878_
timestamp 1698431365
transform 1 0 31136 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _879_
timestamp 1698431365
transform 1 0 30240 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _880_
timestamp 1698431365
transform -1 0 30912 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _881_
timestamp 1698431365
transform 1 0 24304 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _882_
timestamp 1698431365
transform 1 0 23856 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _883_
timestamp 1698431365
transform 1 0 25536 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _884_
timestamp 1698431365
transform -1 0 30912 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _885_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _886_
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _887_
timestamp 1698431365
transform 1 0 9296 0 1 3136
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _888_
timestamp 1698431365
transform 1 0 12432 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _889_
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _890_
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _891_
timestamp 1698431365
transform 1 0 7728 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _892_
timestamp 1698431365
transform -1 0 24864 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _893_
timestamp 1698431365
transform 1 0 18592 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _894_
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _895_
timestamp 1698431365
transform 1 0 8176 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _896_
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _897_
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _898_
timestamp 1698431365
transform 1 0 6944 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _899_
timestamp 1698431365
transform 1 0 14112 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _900_
timestamp 1698431365
transform -1 0 16016 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _901_
timestamp 1698431365
transform 1 0 17360 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _902_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 -1 23520
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _903_
timestamp 1698431365
transform 1 0 21392 0 1 18816
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _904_
timestamp 1698431365
transform 1 0 21280 0 1 21952
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _905_
timestamp 1698431365
transform -1 0 30128 0 -1 23520
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _906_
timestamp 1698431365
transform -1 0 29680 0 -1 25088
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _907_
timestamp 1698431365
transform -1 0 26208 0 1 25088
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _908_
timestamp 1698431365
transform -1 0 29792 0 -1 21952
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _909_
timestamp 1698431365
transform 1 0 22848 0 1 20384
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _910_
timestamp 1698431365
transform 1 0 19488 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _911_
timestamp 1698431365
transform 1 0 13776 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _912_
timestamp 1698431365
transform 1 0 9856 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _913_
timestamp 1698431365
transform 1 0 10976 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _914_
timestamp 1698431365
transform -1 0 21616 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _915_
timestamp 1698431365
transform 1 0 21168 0 -1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _916_
timestamp 1698431365
transform -1 0 24416 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _917_
timestamp 1698431365
transform 1 0 18256 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _918_
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _919_
timestamp 1698431365
transform -1 0 18144 0 1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _920_
timestamp 1698431365
transform -1 0 20048 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _921_
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _922_
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _923_
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _924_
timestamp 1698431365
transform 1 0 1792 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _925_
timestamp 1698431365
transform -1 0 8288 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _926_
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _927_
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__B
timestamp 1698431365
transform 1 0 20272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__I
timestamp 1698431365
transform -1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__B
timestamp 1698431365
transform -1 0 18816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A2
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A3
timestamp 1698431365
transform 1 0 14112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A1
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__A1
timestamp 1698431365
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A2
timestamp 1698431365
transform 1 0 19712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__A1
timestamp 1698431365
transform 1 0 19040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__A1
timestamp 1698431365
transform -1 0 3472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__I
timestamp 1698431365
transform 1 0 32928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__A1
timestamp 1698431365
transform 1 0 24192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__603__I
timestamp 1698431365
transform 1 0 18816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__606__A1
timestamp 1698431365
transform 1 0 20944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__A1
timestamp 1698431365
transform 1 0 18368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__A1
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__I
timestamp 1698431365
transform 1 0 15008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__695__I
timestamp 1698431365
transform 1 0 16128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__724__I
timestamp 1698431365
transform 1 0 17584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__767__I
timestamp 1698431365
transform 1 0 22848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__780__C
timestamp 1698431365
transform 1 0 21392 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__783__B
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__787__B
timestamp 1698431365
transform -1 0 28224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__795__A1
timestamp 1698431365
transform 1 0 26656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__822__C
timestamp 1698431365
transform 1 0 17024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__830__A1
timestamp 1698431365
transform 1 0 21392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__835__A1
timestamp 1698431365
transform 1 0 20496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__837__A1
timestamp 1698431365
transform -1 0 18592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__859__CLK
timestamp 1698431365
transform 1 0 6272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__860__CLK
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__861__CLK
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__862__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__889__CLK
timestamp 1698431365
transform -1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__890__CLK
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__891__CLK
timestamp 1698431365
transform 1 0 12544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__912__CLK
timestamp 1698431365
transform 1 0 9632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 18032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 13552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 19040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 12320 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 19936 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 22512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 25424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 13216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_rebuffer1_I
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18032 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1698431365
transform -1 0 12880 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1698431365
transform -1 0 13104 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1698431365
transform -1 0 19152 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1698431365
transform -1 0 28000 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1698431365
transform 1 0 27104 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1698431365
transform -1 0 28336 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1698431365
transform 1 0 26992 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout5
timestamp 1698431365
transform 1 0 22624 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_40 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_65
timestamp 1698431365
transform 1 0 8624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_128 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15680 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_167
timestamp 1698431365
transform 1 0 20048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_240 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_244
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_280
timestamp 1698431365
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_284
timestamp 1698431365
transform 1 0 33152 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_292
timestamp 1698431365
transform 1 0 34048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_294
timestamp 1698431365
transform 1 0 34272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_90
timestamp 1698431365
transform 1 0 11424 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_128
timestamp 1698431365
transform 1 0 15680 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_156
timestamp 1698431365
transform 1 0 18816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_160
timestamp 1698431365
transform 1 0 19264 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_216
timestamp 1698431365
transform 1 0 25536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_275
timestamp 1698431365
transform 1 0 32144 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_290
timestamp 1698431365
transform 1 0 33824 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_294
timestamp 1698431365
transform 1 0 34272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_6
timestamp 1698431365
transform 1 0 2016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_8
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_39
timestamp 1698431365
transform 1 0 5712 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_148
timestamp 1698431365
transform 1 0 17920 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_187
timestamp 1698431365
transform 1 0 22288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_189
timestamp 1698431365
transform 1 0 22512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_198
timestamp 1698431365
transform 1 0 23520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_239
timestamp 1698431365
transform 1 0 28112 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698431365
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_255
timestamp 1698431365
transform 1 0 29904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_257
timestamp 1698431365
transform 1 0 30128 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_4
timestamp 1698431365
transform 1 0 1792 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_19
timestamp 1698431365
transform 1 0 3472 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_51
timestamp 1698431365
transform 1 0 7056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_120
timestamp 1698431365
transform 1 0 14784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_169
timestamp 1698431365
transform 1 0 20272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_173
timestamp 1698431365
transform 1 0 20720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_195
timestamp 1698431365
transform 1 0 23184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_222
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_238
timestamp 1698431365
transform 1 0 28000 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_242
timestamp 1698431365
transform 1 0 28448 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_249
timestamp 1698431365
transform 1 0 29232 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_259
timestamp 1698431365
transform 1 0 30352 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_290
timestamp 1698431365
transform 1 0 33824 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_294
timestamp 1698431365
transform 1 0 34272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_10
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_14
timestamp 1698431365
transform 1 0 2912 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_16
timestamp 1698431365
transform 1 0 3136 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_21
timestamp 1698431365
transform 1 0 3696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_25
timestamp 1698431365
transform 1 0 4144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_50
timestamp 1698431365
transform 1 0 6944 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_54
timestamp 1698431365
transform 1 0 7392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_71
timestamp 1698431365
transform 1 0 9296 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_80
timestamp 1698431365
transform 1 0 10304 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_102
timestamp 1698431365
transform 1 0 12768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_109
timestamp 1698431365
transform 1 0 13552 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_162
timestamp 1698431365
transform 1 0 19488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_166
timestamp 1698431365
transform 1 0 19936 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_179
timestamp 1698431365
transform 1 0 21392 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_240
timestamp 1698431365
transform 1 0 28224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_255
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_293
timestamp 1698431365
transform 1 0 34160 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_41
timestamp 1698431365
transform 1 0 5936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_45
timestamp 1698431365
transform 1 0 6384 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_77
timestamp 1698431365
transform 1 0 9968 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_113
timestamp 1698431365
transform 1 0 14000 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_194
timestamp 1698431365
transform 1 0 23072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_201
timestamp 1698431365
transform 1 0 23856 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_243
timestamp 1698431365
transform 1 0 28560 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_247
timestamp 1698431365
transform 1 0 29008 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_277
timestamp 1698431365
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_288
timestamp 1698431365
transform 1 0 33600 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_292
timestamp 1698431365
transform 1 0 34048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_294
timestamp 1698431365
transform 1 0 34272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_6
timestamp 1698431365
transform 1 0 2016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_8
timestamp 1698431365
transform 1 0 2240 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_33
timestamp 1698431365
transform 1 0 5040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_57
timestamp 1698431365
transform 1 0 7728 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_61
timestamp 1698431365
transform 1 0 8176 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_164
timestamp 1698431365
transform 1 0 19712 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_189
timestamp 1698431365
transform 1 0 22512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_191
timestamp 1698431365
transform 1 0 22736 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_233
timestamp 1698431365
transform 1 0 27440 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_242
timestamp 1698431365
transform 1 0 28448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_263
timestamp 1698431365
transform 1 0 30800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_265
timestamp 1698431365
transform 1 0 31024 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_6
timestamp 1698431365
transform 1 0 2016 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_40
timestamp 1698431365
transform 1 0 5824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_52
timestamp 1698431365
transform 1 0 7168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_54
timestamp 1698431365
transform 1 0 7392 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_63
timestamp 1698431365
transform 1 0 8400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_205
timestamp 1698431365
transform 1 0 24304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_207
timestamp 1698431365
transform 1 0 24528 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_218
timestamp 1698431365
transform 1 0 25760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_220
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_227
timestamp 1698431365
transform 1 0 26768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_229
timestamp 1698431365
transform 1 0 26992 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_290
timestamp 1698431365
transform 1 0 33824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_294
timestamp 1698431365
transform 1 0 34272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_6
timestamp 1698431365
transform 1 0 2016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_26
timestamp 1698431365
transform 1 0 4256 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_62
timestamp 1698431365
transform 1 0 8288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_64
timestamp 1698431365
transform 1 0 8512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_75
timestamp 1698431365
transform 1 0 9744 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_93
timestamp 1698431365
transform 1 0 11760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_170
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_183
timestamp 1698431365
transform 1 0 21840 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_187
timestamp 1698431365
transform 1 0 22288 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_255
timestamp 1698431365
transform 1 0 29904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_257
timestamp 1698431365
transform 1 0 30128 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_10
timestamp 1698431365
transform 1 0 2464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_25
timestamp 1698431365
transform 1 0 4144 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_29
timestamp 1698431365
transform 1 0 4592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_35
timestamp 1698431365
transform 1 0 5264 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_43
timestamp 1698431365
transform 1 0 6160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_58
timestamp 1698431365
transform 1 0 7840 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_91
timestamp 1698431365
transform 1 0 11536 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_95
timestamp 1698431365
transform 1 0 11984 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_125
timestamp 1698431365
transform 1 0 15344 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_133
timestamp 1698431365
transform 1 0 16240 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_150
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_180
timestamp 1698431365
transform 1 0 21504 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_187
timestamp 1698431365
transform 1 0 22288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_191 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22736 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_222
timestamp 1698431365
transform 1 0 26208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_226
timestamp 1698431365
transform 1 0 26656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_257
timestamp 1698431365
transform 1 0 30128 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_277
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_290
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_294
timestamp 1698431365
transform 1 0 34272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_4
timestamp 1698431365
transform 1 0 1792 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_58
timestamp 1698431365
transform 1 0 7840 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_92
timestamp 1698431365
transform 1 0 11648 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_100
timestamp 1698431365
transform 1 0 12544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_102
timestamp 1698431365
transform 1 0 12768 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_149
timestamp 1698431365
transform 1 0 18032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_153
timestamp 1698431365
transform 1 0 18480 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_156
timestamp 1698431365
transform 1 0 18816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_195
timestamp 1698431365
transform 1 0 23184 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_203
timestamp 1698431365
transform 1 0 24080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_234
timestamp 1698431365
transform 1 0 27552 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1698431365
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_261
timestamp 1698431365
transform 1 0 30576 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_265
timestamp 1698431365
transform 1 0 31024 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_10
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_42
timestamp 1698431365
transform 1 0 6048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_52
timestamp 1698431365
transform 1 0 7168 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_76
timestamp 1698431365
transform 1 0 9856 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_78
timestamp 1698431365
transform 1 0 10080 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_87
timestamp 1698431365
transform 1 0 11088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_89
timestamp 1698431365
transform 1 0 11312 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_208
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_216
timestamp 1698431365
transform 1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_218
timestamp 1698431365
transform 1 0 25760 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_232
timestamp 1698431365
transform 1 0 27328 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_264
timestamp 1698431365
transform 1 0 30912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_266
timestamp 1698431365
transform 1 0 31136 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_275
timestamp 1698431365
transform 1 0 32144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_290
timestamp 1698431365
transform 1 0 33824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_294
timestamp 1698431365
transform 1 0 34272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_10
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_14
timestamp 1698431365
transform 1 0 2912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_16
timestamp 1698431365
transform 1 0 3136 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_47
timestamp 1698431365
transform 1 0 6608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_98
timestamp 1698431365
transform 1 0 12320 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_109
timestamp 1698431365
transform 1 0 13552 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_140
timestamp 1698431365
transform 1 0 17024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_148
timestamp 1698431365
transform 1 0 17920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_195
timestamp 1698431365
transform 1 0 23184 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_199
timestamp 1698431365
transform 1 0 23632 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_235
timestamp 1698431365
transform 1 0 27664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_255
timestamp 1698431365
transform 1 0 29904 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_263
timestamp 1698431365
transform 1 0 30800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_265
timestamp 1698431365
transform 1 0 31024 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_18
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_26
timestamp 1698431365
transform 1 0 4256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_30
timestamp 1698431365
transform 1 0 4704 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_62
timestamp 1698431365
transform 1 0 8288 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_96
timestamp 1698431365
transform 1 0 12096 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_112
timestamp 1698431365
transform 1 0 13888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_116
timestamp 1698431365
transform 1 0 14336 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_132
timestamp 1698431365
transform 1 0 16128 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_154
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_158
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_160
timestamp 1698431365
transform 1 0 19264 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_173
timestamp 1698431365
transform 1 0 20720 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_177
timestamp 1698431365
transform 1 0 21168 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_194
timestamp 1698431365
transform 1 0 23072 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_196
timestamp 1698431365
transform 1 0 23296 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_202
timestamp 1698431365
transform 1 0 23968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_294
timestamp 1698431365
transform 1 0 34272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_31
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_43
timestamp 1698431365
transform 1 0 6160 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_51
timestamp 1698431365
transform 1 0 7056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698431365
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_127
timestamp 1698431365
transform 1 0 15568 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_133
timestamp 1698431365
transform 1 0 16240 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_206
timestamp 1698431365
transform 1 0 24416 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_222
timestamp 1698431365
transform 1 0 26208 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_253
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_286
timestamp 1698431365
transform 1 0 33376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_294
timestamp 1698431365
transform 1 0 34272 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_34
timestamp 1698431365
transform 1 0 5152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_36
timestamp 1698431365
transform 1 0 5376 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_84
timestamp 1698431365
transform 1 0 10752 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_115
timestamp 1698431365
transform 1 0 14224 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_146
timestamp 1698431365
transform 1 0 17696 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_199
timestamp 1698431365
transform 1 0 23632 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698431365
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_218
timestamp 1698431365
transform 1 0 25760 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_225
timestamp 1698431365
transform 1 0 26544 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_247
timestamp 1698431365
transform 1 0 29008 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_255
timestamp 1698431365
transform 1 0 29904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_290
timestamp 1698431365
transform 1 0 33824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_294
timestamp 1698431365
transform 1 0 34272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_41
timestamp 1698431365
transform 1 0 5936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_43
timestamp 1698431365
transform 1 0 6160 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_46
timestamp 1698431365
transform 1 0 6496 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_62
timestamp 1698431365
transform 1 0 8288 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_70
timestamp 1698431365
transform 1 0 9184 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_119
timestamp 1698431365
transform 1 0 14672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_162
timestamp 1698431365
transform 1 0 19488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_170
timestamp 1698431365
transform 1 0 20384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_193
timestamp 1698431365
transform 1 0 22960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_195
timestamp 1698431365
transform 1 0 23184 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_210
timestamp 1698431365
transform 1 0 24864 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_224
timestamp 1698431365
transform 1 0 26432 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_228
timestamp 1698431365
transform 1 0 26880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_230
timestamp 1698431365
transform 1 0 27104 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_259
timestamp 1698431365
transform 1 0 30352 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_263
timestamp 1698431365
transform 1 0 30800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_265
timestamp 1698431365
transform 1 0 31024 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_10
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_14
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_44
timestamp 1698431365
transform 1 0 6272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_46
timestamp 1698431365
transform 1 0 6496 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_53
timestamp 1698431365
transform 1 0 7280 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_78
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_94
timestamp 1698431365
transform 1 0 11872 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698431365
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_118
timestamp 1698431365
transform 1 0 14560 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_241
timestamp 1698431365
transform 1 0 28336 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_245
timestamp 1698431365
transform 1 0 28784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_261
timestamp 1698431365
transform 1 0 30576 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_290
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_294
timestamp 1698431365
transform 1 0 34272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_31
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_65
timestamp 1698431365
transform 1 0 8624 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_90
timestamp 1698431365
transform 1 0 11424 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_98
timestamp 1698431365
transform 1 0 12320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_102
timestamp 1698431365
transform 1 0 12768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_123
timestamp 1698431365
transform 1 0 15120 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_127
timestamp 1698431365
transform 1 0 15568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_137
timestamp 1698431365
transform 1 0 16688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_139
timestamp 1698431365
transform 1 0 16912 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_142
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_155
timestamp 1698431365
transform 1 0 18704 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_160
timestamp 1698431365
transform 1 0 19264 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_168
timestamp 1698431365
transform 1 0 20160 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698431365
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_256
timestamp 1698431365
transform 1 0 30016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_287
timestamp 1698431365
transform 1 0 33488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_34
timestamp 1698431365
transform 1 0 5152 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_103
timestamp 1698431365
transform 1 0 12880 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_191
timestamp 1698431365
transform 1 0 22736 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_200
timestamp 1698431365
transform 1 0 23744 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_214
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_290
timestamp 1698431365
transform 1 0 33824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_294
timestamp 1698431365
transform 1 0 34272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_31
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_45
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_61
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_79
timestamp 1698431365
transform 1 0 10192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_90
timestamp 1698431365
transform 1 0 11424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698431365
transform 1 0 14224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_119
timestamp 1698431365
transform 1 0 14672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_121
timestamp 1698431365
transform 1 0 14896 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_124
timestamp 1698431365
transform 1 0 15232 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_140
timestamp 1698431365
transform 1 0 17024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_150
timestamp 1698431365
transform 1 0 18144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_154
timestamp 1698431365
transform 1 0 18592 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_170
timestamp 1698431365
transform 1 0 20384 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_215
timestamp 1698431365
transform 1 0 25424 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_255
timestamp 1698431365
transform 1 0 29904 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_287
timestamp 1698431365
transform 1 0 33488 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_39
timestamp 1698431365
transform 1 0 5712 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_47
timestamp 1698431365
transform 1 0 6608 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_63
timestamp 1698431365
transform 1 0 8400 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_103
timestamp 1698431365
transform 1 0 12880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_111
timestamp 1698431365
transform 1 0 13776 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_130
timestamp 1698431365
transform 1 0 15904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698431365
transform 1 0 17472 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_161
timestamp 1698431365
transform 1 0 19376 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_169
timestamp 1698431365
transform 1 0 20272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_188
timestamp 1698431365
transform 1 0 22400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_190
timestamp 1698431365
transform 1 0 22624 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_224
timestamp 1698431365
transform 1 0 26432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_228
timestamp 1698431365
transform 1 0 26880 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_264
timestamp 1698431365
transform 1 0 30912 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_290
timestamp 1698431365
transform 1 0 33824 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_294
timestamp 1698431365
transform 1 0 34272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_6
timestamp 1698431365
transform 1 0 2016 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_33
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_74
timestamp 1698431365
transform 1 0 9632 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_93
timestamp 1698431365
transform 1 0 11760 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_97
timestamp 1698431365
transform 1 0 12208 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_118
timestamp 1698431365
transform 1 0 14560 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_126
timestamp 1698431365
transform 1 0 15456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_136
timestamp 1698431365
transform 1 0 16576 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_140
timestamp 1698431365
transform 1 0 17024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_154
timestamp 1698431365
transform 1 0 18592 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_170
timestamp 1698431365
transform 1 0 20384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_181
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_185
timestamp 1698431365
transform 1 0 22064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_187
timestamp 1698431365
transform 1 0 22288 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_236
timestamp 1698431365
transform 1 0 27776 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_279
timestamp 1698431365
transform 1 0 32592 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_10
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_14
timestamp 1698431365
transform 1 0 2912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_16
timestamp 1698431365
transform 1 0 3136 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_40
timestamp 1698431365
transform 1 0 5824 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_56
timestamp 1698431365
transform 1 0 7616 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698431365
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_80
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_87
timestamp 1698431365
transform 1 0 11088 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_95
timestamp 1698431365
transform 1 0 11984 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_130
timestamp 1698431365
transform 1 0 15904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_132
timestamp 1698431365
transform 1 0 16128 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698431365
transform 1 0 17472 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_153
timestamp 1698431365
transform 1 0 18480 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_157
timestamp 1698431365
transform 1 0 18928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_164
timestamp 1698431365
transform 1 0 19712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_254
timestamp 1698431365
transform 1 0 29792 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698431365
transform 1 0 31584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698431365
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_290
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_294
timestamp 1698431365
transform 1 0 34272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_33
timestamp 1698431365
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_45
timestamp 1698431365
transform 1 0 6384 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_53
timestamp 1698431365
transform 1 0 7280 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_214
timestamp 1698431365
transform 1 0 25312 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_239
timestamp 1698431365
transform 1 0 28112 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698431365
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_279
timestamp 1698431365
transform 1 0 32592 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_47
timestamp 1698431365
transform 1 0 6608 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_55
timestamp 1698431365
transform 1 0 7504 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_59
timestamp 1698431365
transform 1 0 7952 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_74
timestamp 1698431365
transform 1 0 9632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_105
timestamp 1698431365
transform 1 0 13104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_107
timestamp 1698431365
transform 1 0 13328 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698431365
transform 1 0 16240 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698431365
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_257
timestamp 1698431365
transform 1 0 30128 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_294
timestamp 1698431365
transform 1 0 34272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_18
timestamp 1698431365
transform 1 0 3360 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_26
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_45
timestamp 1698431365
transform 1 0 6384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_49
timestamp 1698431365
transform 1 0 6832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_79
timestamp 1698431365
transform 1 0 10192 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_83
timestamp 1698431365
transform 1 0 10640 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_99
timestamp 1698431365
transform 1 0 12432 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_116
timestamp 1698431365
transform 1 0 14336 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_118
timestamp 1698431365
transform 1 0 14560 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_150
timestamp 1698431365
transform 1 0 18144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_154
timestamp 1698431365
transform 1 0 18592 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_167
timestamp 1698431365
transform 1 0 20048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_179
timestamp 1698431365
transform 1 0 21392 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_253
timestamp 1698431365
transform 1 0 29680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_257
timestamp 1698431365
transform 1 0 30128 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_289
timestamp 1698431365
transform 1 0 33712 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_293
timestamp 1698431365
transform 1 0 34160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_18
timestamp 1698431365
transform 1 0 3360 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_22
timestamp 1698431365
transform 1 0 3808 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_50
timestamp 1698431365
transform 1 0 6944 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_84
timestamp 1698431365
transform 1 0 10752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_110
timestamp 1698431365
transform 1 0 13664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_112
timestamp 1698431365
transform 1 0 13888 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_130
timestamp 1698431365
transform 1 0 15904 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698431365
transform 1 0 16800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_161
timestamp 1698431365
transform 1 0 19376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_163
timestamp 1698431365
transform 1 0 19600 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_199
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_203
timestamp 1698431365
transform 1 0 24080 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_216
timestamp 1698431365
transform 1 0 25536 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_253
timestamp 1698431365
transform 1 0 29680 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_269
timestamp 1698431365
transform 1 0 31472 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_294
timestamp 1698431365
transform 1 0 34272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_22
timestamp 1698431365
transform 1 0 3808 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_78
timestamp 1698431365
transform 1 0 10080 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_102
timestamp 1698431365
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_139
timestamp 1698431365
transform 1 0 16912 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_147
timestamp 1698431365
transform 1 0 17808 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_151
timestamp 1698431365
transform 1 0 18256 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698431365
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_236
timestamp 1698431365
transform 1 0 27776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698431365
transform 1 0 28224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_279
timestamp 1698431365
transform 1 0 32592 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_31
timestamp 1698431365
transform 1 0 4816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_62
timestamp 1698431365
transform 1 0 8288 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_74
timestamp 1698431365
transform 1 0 9632 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_79
timestamp 1698431365
transform 1 0 10192 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_87
timestamp 1698431365
transform 1 0 11088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_101
timestamp 1698431365
transform 1 0 12656 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_191
timestamp 1698431365
transform 1 0 22736 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_252
timestamp 1698431365
transform 1 0 29568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_268
timestamp 1698431365
transform 1 0 31360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_290
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_294
timestamp 1698431365
transform 1 0 34272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_52
timestamp 1698431365
transform 1 0 7168 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_82
timestamp 1698431365
transform 1 0 10528 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_90
timestamp 1698431365
transform 1 0 11424 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_94
timestamp 1698431365
transform 1 0 11872 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698431365
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_113
timestamp 1698431365
transform 1 0 14000 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698431365
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_185
timestamp 1698431365
transform 1 0 22064 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_189
timestamp 1698431365
transform 1 0 22512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_211
timestamp 1698431365
transform 1 0 24976 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_279
timestamp 1698431365
transform 1 0 32592 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_36
timestamp 1698431365
transform 1 0 5376 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_76
timestamp 1698431365
transform 1 0 9856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_107
timestamp 1698431365
transform 1 0 13328 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_158
timestamp 1698431365
transform 1 0 19040 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_162
timestamp 1698431365
transform 1 0 19488 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_164
timestamp 1698431365
transform 1 0 19712 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_173
timestamp 1698431365
transform 1 0 20720 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_205
timestamp 1698431365
transform 1 0 24304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_290
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_294
timestamp 1698431365
transform 1 0 34272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_53
timestamp 1698431365
transform 1 0 7280 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_90
timestamp 1698431365
transform 1 0 11424 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_98
timestamp 1698431365
transform 1 0 12320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_102
timestamp 1698431365
transform 1 0 12768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_279
timestamp 1698431365
transform 1 0 32592 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_290
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_294
timestamp 1698431365
transform 1 0 34272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_279
timestamp 1698431365
transform 1 0 32592 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_294
timestamp 1698431365
transform 1 0 34272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_36
timestamp 1698431365
transform 1 0 5376 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_70
timestamp 1698431365
transform 1 0 9184 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_138
timestamp 1698431365
transform 1 0 16800 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_172
timestamp 1698431365
transform 1 0 20608 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_206
timestamp 1698431365
transform 1 0 24416 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_240
timestamp 1698431365
transform 1 0 28224 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_274
timestamp 1698431365
transform 1 0 32032 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_290
timestamp 1698431365
transform 1 0 33824 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_294
timestamp 1698431365
transform 1 0 34272 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18032 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698431365
transform 1 0 25088 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698431365
transform -1 0 31808 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_37 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 34608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_38
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 34608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_39
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 34608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_40
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 34608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_41
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 34608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_42
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 34608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_43
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 34608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_44
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 34608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_45
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 34608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_46
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 34608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_47
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 34608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_48
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 34608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_49
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 34608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_50
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 34608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_51
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 34608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_52
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 34608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_53
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 34608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 34608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 34608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 34608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 34608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 34608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 34608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 34608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 34608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 34608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 34608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 34608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 34608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 34608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 34608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 34608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 34608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 34608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 34608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 34608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer1
timestamp 1698431365
transform -1 0 20384 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer2
timestamp 1698431365
transform 1 0 17920 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer3
timestamp 1698431365
transform -1 0 5040 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer4
timestamp 1698431365
transform 1 0 10304 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer5
timestamp 1698431365
transform -1 0 11648 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlya_2  rebuffer6 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24192 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_74 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_75
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_76
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_77
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_78
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_79
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_80
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_81
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_82
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_83
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_84
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_85
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_86
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_87
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_88
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_89
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_90
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_91
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_92
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_93
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_94
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_95
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_96
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_97
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_98
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_99
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_100
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_101
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_102
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_103
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_104
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_105
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_106
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_107
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_108
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_109
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_110
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_111
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_112
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_113
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_114
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_115
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_116
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_117
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_118
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_119
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_120
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_121
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_122
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_123
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_124
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_125
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_126
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_127
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_128
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_129
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_130
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_131
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_132
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_133
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_134
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_135
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_136
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_137
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_138
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_139
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_140
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_141
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_142
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_143
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_144
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_145
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_146
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_147
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_148
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_149
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_150
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_151
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_152
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_153
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_154
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_155
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_156
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_157
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_158
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_159
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_160
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_161
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_162
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_163
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_164
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_165
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_166
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_167
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_168
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_169
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_170
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_171
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_172
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_173
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_174
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_175
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_176
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_177
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_178
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_179
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_180
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_181
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_182
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_183
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_184
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_185
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_186
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_187
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_188
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_189
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_190
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_191
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_192
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_193
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_194
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_195
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_196
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_197
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_198
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_199
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_200
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_201
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_202
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_203
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_204
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_205
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_206
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_207
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_208
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_209
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_210
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_211
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_212
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_213
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_214
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_215
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_216
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_217
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_218
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_219
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_220
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_221
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_222
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_223
timestamp 1698431365
transform 1 0 8960 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_224
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_225
timestamp 1698431365
transform 1 0 16576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_226
timestamp 1698431365
transform 1 0 20384 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_227
timestamp 1698431365
transform 1 0 24192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_228
timestamp 1698431365
transform 1 0 28000 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_229
timestamp 1698431365
transform 1 0 31808 0 1 31360
box -86 -86 310 870
<< labels >>
flabel metal2 s 17920 0 18032 800 0 FreeSans 448 90 0 0 io_out[0]
port 0 nsew signal tristate
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 io_out[1]
port 1 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 io_out[2]
port 2 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 rst_n
port 3 nsew signal input
flabel metal4 s 5342 3076 5662 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 13658 3076 13978 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 21974 3076 22294 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 30290 3076 30610 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 9500 3076 9820 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 17816 3076 18136 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 26132 3076 26452 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 34448 3076 34768 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal2 s 3584 0 3696 800 0 FreeSans 448 90 0 0 wb_clk_i
port 6 nsew signal input
rlabel metal1 17976 32144 17976 32144 0 vdd
rlabel via1 18056 31360 18056 31360 0 vss
rlabel metal3 12768 26264 12768 26264 0 LFSR\[0\]
rlabel metal2 11704 27832 11704 27832 0 LFSR\[1\]
rlabel metal2 11144 24192 11144 24192 0 LFSR\[2\]
rlabel metal2 9912 24416 9912 24416 0 LFSR\[3\]
rlabel metal2 11648 23016 11648 23016 0 LFSR\[4\]
rlabel metal3 16800 27160 16800 27160 0 LFSR\[5\]
rlabel metal2 16408 25088 16408 25088 0 LFSR\[6\]
rlabel metal2 21672 17248 21672 17248 0 OP_reg
rlabel metal2 17976 8624 17976 8624 0 PC\[0\]
rlabel metal2 13832 6440 13832 6440 0 PC\[1\]
rlabel metal3 18480 6104 18480 6104 0 PC\[2\]
rlabel metal2 3416 12488 3416 12488 0 PC\[3\]
rlabel metal2 5656 13944 5656 13944 0 PC\[4\]
rlabel metal2 10808 13328 10808 13328 0 PC\[5\]
rlabel metal2 13048 11144 13048 11144 0 _000_
rlabel metal3 12824 11480 12824 11480 0 _001_
rlabel metal3 4928 16856 4928 16856 0 _002_
rlabel metal2 2408 14504 2408 14504 0 _003_
rlabel metal2 2968 15120 2968 15120 0 _004_
rlabel metal2 6440 15148 6440 15148 0 _005_
rlabel metal2 21784 9744 21784 9744 0 _006_
rlabel metal2 21336 6048 21336 6048 0 _007_
rlabel metal2 21560 4312 21560 4312 0 _008_
rlabel metal3 22008 4200 22008 4200 0 _009_
rlabel metal2 23800 8624 23800 8624 0 _010_
rlabel metal3 26572 4984 26572 4984 0 _011_
rlabel metal2 27944 4536 27944 4536 0 _012_
rlabel metal2 31192 4648 31192 4648 0 _013_
rlabel metal2 30520 5152 30520 5152 0 _014_
rlabel metal2 32088 5432 32088 5432 0 _015_
rlabel metal2 32088 7896 32088 7896 0 _016_
rlabel metal2 33208 9464 33208 9464 0 _017_
rlabel metal2 29512 9744 29512 9744 0 _018_
rlabel metal2 33432 11704 33432 11704 0 _019_
rlabel metal2 33432 13384 33432 13384 0 _020_
rlabel metal2 32424 15960 32424 15960 0 _021_
rlabel metal2 32424 15456 32424 15456 0 _022_
rlabel metal2 29736 13384 29736 13384 0 _023_
rlabel metal2 25704 10864 25704 10864 0 _024_
rlabel metal2 24808 13272 24808 13272 0 _025_
rlabel metal2 27160 19544 27160 19544 0 _026_
rlabel metal2 29624 17360 29624 17360 0 _027_
rlabel metal2 25984 15176 25984 15176 0 _028_
rlabel metal2 16072 6384 16072 6384 0 _029_
rlabel metal2 10248 3864 10248 3864 0 _030_
rlabel metal2 11928 6328 11928 6328 0 _031_
rlabel metal2 2912 5208 2912 5208 0 _032_
rlabel metal2 2520 12992 2520 12992 0 _033_
rlabel metal3 9856 12264 9856 12264 0 _034_
rlabel metal2 24472 16464 24472 16464 0 _035_
rlabel metal2 19544 18816 19544 18816 0 _036_
rlabel metal2 12264 27440 12264 27440 0 _037_
rlabel metal2 9520 28504 9520 28504 0 _038_
rlabel metal2 8904 25704 8904 25704 0 _039_
rlabel metal2 8792 23744 8792 23744 0 _040_
rlabel metal2 8344 23576 8344 23576 0 _041_
rlabel metal2 15400 25984 15400 25984 0 _042_
rlabel metal2 14504 25872 14504 25872 0 _043_
rlabel metal2 18200 26488 18200 26488 0 _044_
rlabel metal2 20328 23296 20328 23296 0 _045_
rlabel metal2 22400 19320 22400 19320 0 _046_
rlabel metal3 21448 22232 21448 22232 0 _047_
rlabel metal2 29232 23240 29232 23240 0 _048_
rlabel metal2 28728 24864 28728 24864 0 _049_
rlabel metal3 25984 25256 25984 25256 0 _050_
rlabel metal2 27496 21168 27496 21168 0 _051_
rlabel metal2 24360 20272 24360 20272 0 _052_
rlabel metal2 20384 26376 20384 26376 0 _053_
rlabel metal2 16072 18032 16072 18032 0 _054_
rlabel metal2 10808 16520 10808 16520 0 _055_
rlabel metal2 11928 15624 11928 15624 0 _056_
rlabel metal2 20664 17192 20664 17192 0 _057_
rlabel metal2 22120 12488 22120 12488 0 _058_
rlabel metal3 22568 14616 22568 14616 0 _059_
rlabel metal3 20328 9912 20328 9912 0 _060_
rlabel metal2 18200 12488 18200 12488 0 _061_
rlabel metal2 15960 23576 15960 23576 0 _062_
rlabel metal2 19768 3304 19768 3304 0 _063_
rlabel metal2 2520 20328 2520 20328 0 _064_
rlabel metal2 2520 19600 2520 19600 0 _065_
rlabel metal2 2520 22792 2520 22792 0 _066_
rlabel metal2 2744 22680 2744 22680 0 _067_
rlabel metal3 6832 26376 6832 26376 0 _068_
rlabel metal2 3304 26040 3304 26040 0 _069_
rlabel metal2 2632 25928 2632 25928 0 _070_
rlabel metal2 11704 3220 11704 3220 0 _071_
rlabel metal2 8568 12824 8568 12824 0 _072_
rlabel metal2 13552 9576 13552 9576 0 _073_
rlabel metal2 16072 8848 16072 8848 0 _074_
rlabel metal2 16856 10472 16856 10472 0 _075_
rlabel metal2 23464 23856 23464 23856 0 _076_
rlabel metal2 22792 22680 22792 22680 0 _077_
rlabel metal2 22456 24304 22456 24304 0 _078_
rlabel metal2 23464 25760 23464 25760 0 _079_
rlabel metal2 16968 14784 16968 14784 0 _080_
rlabel metal2 16184 19040 16184 19040 0 _081_
rlabel metal3 19488 19320 19488 19320 0 _082_
rlabel metal2 4648 25424 4648 25424 0 _083_
rlabel metal2 6216 22680 6216 22680 0 _084_
rlabel metal2 5768 21112 5768 21112 0 _085_
rlabel metal2 16296 13328 16296 13328 0 _086_
rlabel metal2 17640 20720 17640 20720 0 _087_
rlabel metal3 17976 15400 17976 15400 0 _088_
rlabel metal3 18704 15848 18704 15848 0 _089_
rlabel metal2 18200 14056 18200 14056 0 _090_
rlabel metal2 19880 12208 19880 12208 0 _091_
rlabel metal2 19544 13216 19544 13216 0 _092_
rlabel metal2 18312 12600 18312 12600 0 _093_
rlabel metal2 17304 11648 17304 11648 0 _094_
rlabel metal2 17752 9296 17752 9296 0 _095_
rlabel metal2 15848 11536 15848 11536 0 _096_
rlabel metal3 10640 13832 10640 13832 0 _097_
rlabel metal3 11704 12712 11704 12712 0 _098_
rlabel metal3 12824 8232 12824 8232 0 _099_
rlabel metal2 16184 7000 16184 7000 0 _100_
rlabel metal2 11928 9072 11928 9072 0 _101_
rlabel metal2 11704 13216 11704 13216 0 _102_
rlabel metal2 11256 13384 11256 13384 0 _103_
rlabel metal2 9912 11816 9912 11816 0 _104_
rlabel metal2 2856 10696 2856 10696 0 _105_
rlabel metal2 15736 7448 15736 7448 0 _106_
rlabel metal2 11200 7448 11200 7448 0 _107_
rlabel metal2 4872 7504 4872 7504 0 _108_
rlabel metal2 5656 8344 5656 8344 0 _109_
rlabel metal2 12488 6384 12488 6384 0 _110_
rlabel metal2 6328 5936 6328 5936 0 _111_
rlabel metal2 18312 8904 18312 8904 0 _112_
rlabel metal2 17192 7336 17192 7336 0 _113_
rlabel metal3 10080 3304 10080 3304 0 _114_
rlabel metal3 18200 4984 18200 4984 0 _115_
rlabel metal2 15960 6720 15960 6720 0 _116_
rlabel metal2 14056 5880 14056 5880 0 _117_
rlabel metal2 8456 4480 8456 4480 0 _118_
rlabel metal2 7448 3976 7448 3976 0 _119_
rlabel metal3 18200 23016 18200 23016 0 _120_
rlabel metal2 16744 5040 16744 5040 0 _121_
rlabel metal2 12656 6552 12656 6552 0 _122_
rlabel metal2 12152 6720 12152 6720 0 _123_
rlabel metal2 10248 6608 10248 6608 0 _124_
rlabel metal3 11032 9800 11032 9800 0 _125_
rlabel metal3 6664 13832 6664 13832 0 _126_
rlabel metal2 7448 13496 7448 13496 0 _127_
rlabel metal2 7952 12152 7952 12152 0 _128_
rlabel metal2 10136 9520 10136 9520 0 _129_
rlabel metal2 17472 7336 17472 7336 0 _130_
rlabel metal2 16296 5096 16296 5096 0 _131_
rlabel metal2 8904 7504 8904 7504 0 _132_
rlabel metal2 3080 6160 3080 6160 0 _133_
rlabel metal2 2520 5432 2520 5432 0 _134_
rlabel metal3 10976 4424 10976 4424 0 _135_
rlabel metal2 7672 8848 7672 8848 0 _136_
rlabel metal2 11704 6104 11704 6104 0 _137_
rlabel metal2 6440 5096 6440 5096 0 _138_
rlabel metal2 6104 3304 6104 3304 0 _139_
rlabel metal3 6048 5880 6048 5880 0 _140_
rlabel metal3 9856 6776 9856 6776 0 _141_
rlabel metal2 7560 11760 7560 11760 0 _142_
rlabel metal2 10024 9520 10024 9520 0 _143_
rlabel metal2 10360 9968 10360 9968 0 _144_
rlabel metal2 4984 11312 4984 11312 0 _145_
rlabel metal3 3136 6104 3136 6104 0 _146_
rlabel metal2 8232 5824 8232 5824 0 _147_
rlabel metal2 11312 4312 11312 4312 0 _148_
rlabel metal2 8120 9044 8120 9044 0 _149_
rlabel metal2 8008 10696 8008 10696 0 _150_
rlabel metal2 15400 4256 15400 4256 0 _151_
rlabel metal2 5880 6888 5880 6888 0 _152_
rlabel metal2 6552 6384 6552 6384 0 _153_
rlabel metal2 8400 8008 8400 8008 0 _154_
rlabel metal2 8064 6104 8064 6104 0 _155_
rlabel metal2 9184 8344 9184 8344 0 _156_
rlabel metal2 3192 11984 3192 11984 0 _157_
rlabel metal2 10752 11480 10752 11480 0 _158_
rlabel metal2 8792 10864 8792 10864 0 _159_
rlabel metal2 3976 5824 3976 5824 0 _160_
rlabel metal2 10472 10752 10472 10752 0 _161_
rlabel metal3 7112 10528 7112 10528 0 _162_
rlabel metal3 10640 8232 10640 8232 0 _163_
rlabel metal3 6496 7560 6496 7560 0 _164_
rlabel metal2 5600 7448 5600 7448 0 _165_
rlabel metal4 9912 9296 9912 9296 0 _166_
rlabel metal3 5488 8232 5488 8232 0 _167_
rlabel metal2 10360 10976 10360 10976 0 _168_
rlabel metal2 8680 10136 8680 10136 0 _169_
rlabel metal2 8456 10920 8456 10920 0 _170_
rlabel metal2 9016 10976 9016 10976 0 _171_
rlabel metal2 8232 6384 8232 6384 0 _172_
rlabel metal2 5096 6832 5096 6832 0 _173_
rlabel metal2 3304 9520 3304 9520 0 _174_
rlabel metal2 4984 7112 4984 7112 0 _175_
rlabel metal2 3640 7840 3640 7840 0 _176_
rlabel metal2 5152 7672 5152 7672 0 _177_
rlabel metal2 9352 5376 9352 5376 0 _178_
rlabel metal2 6664 8736 6664 8736 0 _179_
rlabel metal3 5208 9016 5208 9016 0 _180_
rlabel metal3 6048 9128 6048 9128 0 _181_
rlabel metal2 2968 9632 2968 9632 0 _182_
rlabel metal2 5880 8792 5880 8792 0 _183_
rlabel metal2 6776 7728 6776 7728 0 _184_
rlabel metal3 4424 9912 4424 9912 0 _185_
rlabel metal2 4536 7616 4536 7616 0 _186_
rlabel metal2 5208 8512 5208 8512 0 _187_
rlabel metal2 2856 7336 2856 7336 0 _188_
rlabel metal2 3080 10304 3080 10304 0 _189_
rlabel metal2 2296 10304 2296 10304 0 _190_
rlabel metal2 2520 11032 2520 11032 0 _191_
rlabel metal2 4648 12768 4648 12768 0 _192_
rlabel metal2 2744 8372 2744 8372 0 _193_
rlabel metal2 3752 7672 3752 7672 0 _194_
rlabel metal2 3920 9240 3920 9240 0 _195_
rlabel metal2 3696 10808 3696 10808 0 _196_
rlabel metal2 2968 7952 2968 7952 0 _197_
rlabel metal3 3024 8344 3024 8344 0 _198_
rlabel metal3 6048 12936 6048 12936 0 _199_
rlabel metal3 5320 12152 5320 12152 0 _200_
rlabel metal2 3864 12544 3864 12544 0 _201_
rlabel metal2 7168 11928 7168 11928 0 _202_
rlabel metal2 5432 12544 5432 12544 0 _203_
rlabel metal2 6328 10416 6328 10416 0 _204_
rlabel metal2 3920 11368 3920 11368 0 _205_
rlabel metal2 4760 10920 4760 10920 0 _206_
rlabel metal2 4312 12208 4312 12208 0 _207_
rlabel metal2 6608 13160 6608 13160 0 _208_
rlabel metal2 5992 11312 5992 11312 0 _209_
rlabel metal2 6328 12824 6328 12824 0 _210_
rlabel metal2 24024 15568 24024 15568 0 _211_
rlabel metal2 23632 18424 23632 18424 0 _212_
rlabel metal2 22232 6720 22232 6720 0 _213_
rlabel metal3 23912 6552 23912 6552 0 _214_
rlabel metal2 30184 6440 30184 6440 0 _215_
rlabel metal2 23072 5992 23072 5992 0 _216_
rlabel metal3 30128 8232 30128 8232 0 _217_
rlabel metal2 30632 9576 30632 9576 0 _218_
rlabel metal3 28728 8120 28728 8120 0 _219_
rlabel metal2 24248 5936 24248 5936 0 _220_
rlabel metal2 27608 7952 27608 7952 0 _221_
rlabel metal2 28168 8008 28168 8008 0 _222_
rlabel metal2 30856 14896 30856 14896 0 _223_
rlabel metal2 28168 15624 28168 15624 0 _224_
rlabel metal3 27048 15960 27048 15960 0 _225_
rlabel metal2 28448 15512 28448 15512 0 _226_
rlabel metal2 24136 6888 24136 6888 0 _227_
rlabel metal2 23800 7000 23800 7000 0 _228_
rlabel metal2 25480 14056 25480 14056 0 _229_
rlabel metal2 26824 11760 26824 11760 0 _230_
rlabel metal2 25816 12544 25816 12544 0 _231_
rlabel metal2 19656 13776 19656 13776 0 _232_
rlabel metal2 21448 18592 21448 18592 0 _233_
rlabel metal2 23352 7784 23352 7784 0 _234_
rlabel metal2 23800 4760 23800 4760 0 _235_
rlabel metal3 22344 4536 22344 4536 0 _236_
rlabel metal2 21952 5320 21952 5320 0 _237_
rlabel metal2 24696 3752 24696 3752 0 _238_
rlabel metal3 24640 7448 24640 7448 0 _239_
rlabel metal2 24360 5040 24360 5040 0 _240_
rlabel metal2 25256 8008 25256 8008 0 _241_
rlabel metal3 27440 5880 27440 5880 0 _242_
rlabel metal2 27384 5488 27384 5488 0 _243_
rlabel metal3 27608 5712 27608 5712 0 _244_
rlabel metal2 26712 6552 26712 6552 0 _245_
rlabel metal2 29288 7448 29288 7448 0 _246_
rlabel metal2 29288 5096 29288 5096 0 _247_
rlabel via2 30072 6776 30072 6776 0 _248_
rlabel metal3 32088 5880 32088 5880 0 _249_
rlabel metal2 30072 18144 30072 18144 0 _250_
rlabel metal2 30408 16856 30408 16856 0 _251_
rlabel metal2 31024 5096 31024 5096 0 _252_
rlabel metal3 32480 5768 32480 5768 0 _253_
rlabel metal2 30744 6776 30744 6776 0 _254_
rlabel metal2 30968 10640 30968 10640 0 _255_
rlabel metal2 32928 7560 32928 7560 0 _256_
rlabel metal3 32760 9016 32760 9016 0 _257_
rlabel metal3 29456 9800 29456 9800 0 _258_
rlabel metal2 29288 10472 29288 10472 0 _259_
rlabel metal2 29624 13720 29624 13720 0 _260_
rlabel metal2 31640 11368 31640 11368 0 _261_
rlabel metal2 30856 10080 30856 10080 0 _262_
rlabel metal2 31304 13552 31304 13552 0 _263_
rlabel metal3 31584 15176 31584 15176 0 _264_
rlabel metal2 32536 16856 32536 16856 0 _265_
rlabel metal2 32760 14840 32760 14840 0 _266_
rlabel metal2 32256 14728 32256 14728 0 _267_
rlabel metal2 32032 15400 32032 15400 0 _268_
rlabel metal2 26712 12880 26712 12880 0 _269_
rlabel metal2 28840 14000 28840 14000 0 _270_
rlabel metal2 26040 11424 26040 11424 0 _271_
rlabel metal3 26880 13608 26880 13608 0 _272_
rlabel metal2 29064 15960 29064 15960 0 _273_
rlabel metal2 29176 19600 29176 19600 0 _274_
rlabel metal2 29176 16184 29176 16184 0 _275_
rlabel metal2 29288 17920 29288 17920 0 _276_
rlabel metal2 25816 17304 25816 17304 0 _277_
rlabel metal2 26488 15400 26488 15400 0 _278_
rlabel metal2 22232 20048 22232 20048 0 _279_
rlabel metal2 19320 22400 19320 22400 0 _280_
rlabel metal2 18536 17304 18536 17304 0 _281_
rlabel metal2 18648 12768 18648 12768 0 _282_
rlabel metal3 22568 12936 22568 12936 0 _283_
rlabel metal3 19600 12376 19600 12376 0 _284_
rlabel metal2 22232 15540 22232 15540 0 _285_
rlabel metal3 23520 15960 23520 15960 0 _286_
rlabel metal3 16072 21784 16072 21784 0 _287_
rlabel metal2 15624 24192 15624 24192 0 _288_
rlabel metal3 12320 23912 12320 23912 0 _289_
rlabel metal2 13440 23912 13440 23912 0 _290_
rlabel metal2 13832 23688 13832 23688 0 _291_
rlabel metal3 13048 21784 13048 21784 0 _292_
rlabel metal2 14392 20720 14392 20720 0 _293_
rlabel metal2 18312 19936 18312 19936 0 _294_
rlabel metal2 16632 20048 16632 20048 0 _295_
rlabel metal2 16632 25592 16632 25592 0 _296_
rlabel metal3 18424 19992 18424 19992 0 _297_
rlabel metal2 19656 22568 19656 22568 0 _298_
rlabel metal3 15120 27048 15120 27048 0 _299_
rlabel metal3 17248 15512 17248 15512 0 _300_
rlabel metal2 15848 23408 15848 23408 0 _301_
rlabel metal3 12824 21672 12824 21672 0 _302_
rlabel metal2 7112 17864 7112 17864 0 _303_
rlabel metal2 11424 18424 11424 18424 0 _304_
rlabel metal2 7672 17248 7672 17248 0 _305_
rlabel metal2 10472 17192 10472 17192 0 _306_
rlabel metal2 8232 18704 8232 18704 0 _307_
rlabel metal2 11256 17304 11256 17304 0 _308_
rlabel metal2 10920 19208 10920 19208 0 _309_
rlabel metal2 7280 19880 7280 19880 0 _310_
rlabel metal2 8680 19488 8680 19488 0 _311_
rlabel metal2 9464 18536 9464 18536 0 _312_
rlabel metal2 12208 20216 12208 20216 0 _313_
rlabel metal3 12320 24920 12320 24920 0 _314_
rlabel metal2 18312 22456 18312 22456 0 _315_
rlabel metal2 17528 24976 17528 24976 0 _316_
rlabel metal3 13160 25592 13160 25592 0 _317_
rlabel metal2 14168 23520 14168 23520 0 _318_
rlabel metal2 9912 17920 9912 17920 0 _319_
rlabel metal3 8456 18536 8456 18536 0 _320_
rlabel metal2 7672 19208 7672 19208 0 _321_
rlabel metal2 8680 18536 8680 18536 0 _322_
rlabel metal3 9520 18200 9520 18200 0 _323_
rlabel metal2 10696 18928 10696 18928 0 _324_
rlabel metal2 11480 21280 11480 21280 0 _325_
rlabel metal2 12040 24136 12040 24136 0 _326_
rlabel metal2 11312 23128 11312 23128 0 _327_
rlabel metal3 17248 23240 17248 23240 0 _328_
rlabel metal2 10024 25536 10024 25536 0 _329_
rlabel metal2 11536 18648 11536 18648 0 _330_
rlabel metal2 8232 18200 8232 18200 0 _331_
rlabel metal2 12712 19488 12712 19488 0 _332_
rlabel metal2 12040 20776 12040 20776 0 _333_
rlabel metal2 10248 23184 10248 23184 0 _334_
rlabel metal3 11032 23912 11032 23912 0 _335_
rlabel metal2 9016 24304 9016 24304 0 _336_
rlabel metal2 10248 20328 10248 20328 0 _337_
rlabel metal2 12768 20216 12768 20216 0 _338_
rlabel metal2 15512 21280 15512 21280 0 _339_
rlabel metal2 15176 22736 15176 22736 0 _340_
rlabel metal2 12488 22848 12488 22848 0 _341_
rlabel metal2 13160 22344 13160 22344 0 _342_
rlabel metal3 10752 23016 10752 23016 0 _343_
rlabel metal2 9912 18368 9912 18368 0 _344_
rlabel metal2 12656 18648 12656 18648 0 _345_
rlabel metal2 10864 17864 10864 17864 0 _346_
rlabel metal2 12264 19264 12264 19264 0 _347_
rlabel metal2 13832 20832 13832 20832 0 _348_
rlabel metal3 14168 21672 14168 21672 0 _349_
rlabel metal2 13720 22008 13720 22008 0 _350_
rlabel metal2 8904 19152 8904 19152 0 _351_
rlabel metal2 8008 19600 8008 19600 0 _352_
rlabel metal2 9240 19264 9240 19264 0 _353_
rlabel metal3 9800 19320 9800 19320 0 _354_
rlabel metal2 10360 19992 10360 19992 0 _355_
rlabel metal2 15176 25200 15176 25200 0 _356_
rlabel metal2 16128 25368 16128 25368 0 _357_
rlabel metal2 15904 25480 15904 25480 0 _358_
rlabel metal2 12544 25480 12544 25480 0 _359_
rlabel metal2 10584 21112 10584 21112 0 _360_
rlabel metal2 11032 21336 11032 21336 0 _361_
rlabel metal2 14280 25368 14280 25368 0 _362_
rlabel metal3 15708 25256 15708 25256 0 _363_
rlabel metal2 18536 25760 18536 25760 0 _364_
rlabel metal2 23240 18368 23240 18368 0 _365_
rlabel metal3 18592 26264 18592 26264 0 _366_
rlabel metal3 22624 21672 22624 21672 0 _367_
rlabel metal2 19488 24024 19488 24024 0 _368_
rlabel metal2 19656 20776 19656 20776 0 _369_
rlabel metal2 18872 23576 18872 23576 0 _370_
rlabel metal3 21728 19880 21728 19880 0 _371_
rlabel metal3 21504 21000 21504 21000 0 _372_
rlabel metal2 20888 22008 20888 22008 0 _373_
rlabel metal2 25480 23184 25480 23184 0 _374_
rlabel metal2 25816 23688 25816 23688 0 _375_
rlabel metal2 26712 21000 26712 21000 0 _376_
rlabel metal3 28168 23800 28168 23800 0 _377_
rlabel metal2 26152 22848 26152 22848 0 _378_
rlabel metal2 25816 25816 25816 25816 0 _379_
rlabel metal2 28056 24696 28056 24696 0 _380_
rlabel metal2 26600 25088 26600 25088 0 _381_
rlabel metal2 26376 25984 26376 25984 0 _382_
rlabel metal2 27384 21224 27384 21224 0 _383_
rlabel metal2 25928 21672 25928 21672 0 _384_
rlabel metal2 25704 21672 25704 21672 0 _385_
rlabel metal2 27048 21056 27048 21056 0 _386_
rlabel metal3 24976 19992 24976 19992 0 _387_
rlabel metal3 19656 27832 19656 27832 0 _388_
rlabel metal2 19992 26712 19992 26712 0 _389_
rlabel metal2 16184 17584 16184 17584 0 _390_
rlabel metal2 15792 15512 15792 15512 0 _391_
rlabel metal2 16632 16464 16632 16464 0 _392_
rlabel metal2 15848 17360 15848 17360 0 _393_
rlabel metal2 17528 17640 17528 17640 0 _394_
rlabel metal2 16520 17976 16520 17976 0 _395_
rlabel metal2 16016 15288 16016 15288 0 _396_
rlabel metal2 15400 16016 15400 16016 0 _397_
rlabel metal2 13944 16744 13944 16744 0 _398_
rlabel metal2 12376 16800 12376 16800 0 _399_
rlabel metal2 14952 15792 14952 15792 0 _400_
rlabel metal2 15176 16016 15176 16016 0 _401_
rlabel metal3 14504 15960 14504 15960 0 _402_
rlabel metal3 13272 16184 13272 16184 0 _403_
rlabel metal2 19320 16352 19320 16352 0 _404_
rlabel metal3 17864 15960 17864 15960 0 _405_
rlabel metal2 17416 16352 17416 16352 0 _406_
rlabel metal2 18200 16912 18200 16912 0 _407_
rlabel metal2 22848 11592 22848 11592 0 _408_
rlabel metal3 22288 12824 22288 12824 0 _409_
rlabel metal2 20832 15960 20832 15960 0 _410_
rlabel metal3 20552 10024 20552 10024 0 _411_
rlabel metal2 21560 11928 21560 11928 0 _412_
rlabel metal2 19600 5768 19600 5768 0 _413_
rlabel metal3 2688 20552 2688 20552 0 _414_
rlabel metal2 17416 22736 17416 22736 0 _415_
rlabel metal2 2632 23240 2632 23240 0 _416_
rlabel metal2 4536 20272 4536 20272 0 _417_
rlabel metal2 5432 20048 5432 20048 0 _418_
rlabel metal2 5208 23464 5208 23464 0 _419_
rlabel metal2 3640 22064 3640 22064 0 _420_
rlabel metal2 5096 24808 5096 24808 0 _421_
rlabel metal2 5880 23184 5880 23184 0 _422_
rlabel metal3 6384 27048 6384 27048 0 _423_
rlabel metal3 5544 27272 5544 27272 0 _424_
rlabel metal2 3864 25368 3864 25368 0 _425_
rlabel metal2 4704 27832 4704 27832 0 _426_
rlabel metal2 2968 26712 2968 26712 0 _427_
rlabel metal2 19936 21784 19936 21784 0 clknet_0_wb_clk_i
rlabel metal2 3304 15960 3304 15960 0 clknet_3_0__leaf_wb_clk_i
rlabel metal3 12376 15288 12376 15288 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 1904 23128 1904 23128 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 14392 26992 14392 26992 0 clknet_3_3__leaf_wb_clk_i
rlabel metal2 24472 12152 24472 12152 0 clknet_3_4__leaf_wb_clk_i
rlabel metal2 34104 12152 34104 12152 0 clknet_3_5__leaf_wb_clk_i
rlabel metal3 22232 20776 22232 20776 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 25928 25144 25928 25144 0 clknet_3_7__leaf_wb_clk_i
rlabel metal2 23912 23632 23912 23632 0 clock_div\[0\]
rlabel metal2 24024 19712 24024 19712 0 clock_div\[1\]
rlabel metal2 24472 22120 24472 22120 0 clock_div\[2\]
rlabel metal2 26824 23352 26824 23352 0 clock_div\[3\]
rlabel metal2 26600 24584 26600 24584 0 clock_div\[4\]
rlabel metal3 23688 24920 23688 24920 0 clock_div\[5\]
rlabel metal2 26152 21504 26152 21504 0 clock_div\[6\]
rlabel metal3 25256 20888 25256 20888 0 clock_div\[7\]
rlabel metal3 23352 26152 23352 26152 0 clock_div\[8\]
rlabel metal2 22344 8400 22344 8400 0 counter\[0\]
rlabel metal2 33432 7896 33432 7896 0 counter\[10\]
rlabel metal2 31304 10248 31304 10248 0 counter\[11\]
rlabel metal2 30856 10528 30856 10528 0 counter\[12\]
rlabel metal3 30184 9800 30184 9800 0 counter\[13\]
rlabel metal2 31304 14392 31304 14392 0 counter\[14\]
rlabel metal2 33656 15736 33656 15736 0 counter\[15\]
rlabel metal2 31976 17416 31976 17416 0 counter\[16\]
rlabel metal3 30184 15288 30184 15288 0 counter\[17\]
rlabel via2 26376 13384 26376 13384 0 counter\[18\]
rlabel metal2 27384 13160 27384 13160 0 counter\[19\]
rlabel metal3 22400 7448 22400 7448 0 counter\[1\]
rlabel metal2 29176 17080 29176 17080 0 counter\[20\]
rlabel metal3 28728 16968 28728 16968 0 counter\[21\]
rlabel metal2 26096 18424 26096 18424 0 counter\[22\]
rlabel metal2 22456 3864 22456 3864 0 counter\[3\]
rlabel metal2 25928 8288 25928 8288 0 counter\[4\]
rlabel metal3 24696 5880 24696 5880 0 counter\[5\]
rlabel metal2 26040 6832 26040 6832 0 counter\[6\]
rlabel metal2 28952 5096 28952 5096 0 counter\[7\]
rlabel metal2 33432 6048 33432 6048 0 counter\[8\]
rlabel metal2 33600 5880 33600 5880 0 counter\[9\]
rlabel metal2 17976 1638 17976 1638 0 io_out[0]
rlabel metal2 25144 2086 25144 2086 0 io_out[1]
rlabel metal3 31192 3416 31192 3416 0 io_out[2]
rlabel metal3 22120 16072 22120 16072 0 just_inc
rlabel metal2 15960 16408 15960 16408 0 just_rst
rlabel metal2 4536 21280 4536 21280 0 master_clk_div\[0\]
rlabel metal3 6104 20664 6104 20664 0 master_clk_div\[1\]
rlabel metal3 4312 21672 4312 21672 0 master_clk_div\[2\]
rlabel metal2 4928 23016 4928 23016 0 master_clk_div\[3\]
rlabel metal3 6048 26936 6048 26936 0 master_clk_div\[4\]
rlabel metal2 5040 27160 5040 27160 0 master_clk_div\[5\]
rlabel metal2 4312 27356 4312 27356 0 master_clk_div\[6\]
rlabel metal2 11256 4816 11256 4816 0 net1
rlabel metal2 9800 7644 9800 7644 0 net10
rlabel metal3 22064 19992 22064 19992 0 net11
rlabel metal3 17584 5096 17584 5096 0 net2
rlabel metal2 22792 6272 22792 6272 0 net3
rlabel metal3 31864 3528 31864 3528 0 net4
rlabel metal2 23352 4144 23352 4144 0 net5
rlabel metal2 19656 9352 19656 9352 0 net6
rlabel metal3 18984 13944 18984 13944 0 net7
rlabel metal2 2296 7728 2296 7728 0 net8
rlabel metal2 10864 8120 10864 8120 0 net9
rlabel metal3 21560 26600 21560 26600 0 prev_clk_div
rlabel metal2 16856 16576 16856 16576 0 rhythm_LFSR\[0\]
rlabel metal3 17304 16968 17304 16968 0 rhythm_LFSR\[1\]
rlabel metal3 16408 15344 16408 15344 0 rhythm_LFSR\[2\]
rlabel metal2 17640 16856 17640 16856 0 rhythm_LFSR\[3\]
rlabel metal2 10808 2058 10808 2058 0 rst_n
rlabel metal2 22456 12264 22456 12264 0 tempo_LFSR\[0\]
rlabel metal3 22512 13496 22512 13496 0 tempo_LFSR\[1\]
rlabel metal2 22232 13832 22232 13832 0 tempo_LFSR\[2\]
rlabel metal2 20552 11760 20552 11760 0 tempo_LFSR\[3\]
rlabel metal2 15736 15904 15736 15904 0 tune_ROM\[0\]
rlabel metal2 15848 13552 15848 13552 0 tune_ROM\[1\]
rlabel metal2 6328 17192 6328 17192 0 tune_ROM\[2\]
rlabel metal3 6160 17640 6160 17640 0 tune_ROM\[3\]
rlabel metal3 5936 16968 5936 16968 0 tune_ROM\[4\]
rlabel metal2 8904 16016 8904 16016 0 tune_ROM\[5\]
rlabel metal2 1624 9688 1624 9688 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 36000 36000
<< end >>
