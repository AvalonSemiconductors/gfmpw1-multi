magic
tech gf180mcuD
magscale 1 10
timestamp 1702244006
<< metal1 >>
rect 41122 240494 41134 240546
rect 41186 240543 41198 240546
rect 44146 240543 44158 240546
rect 41186 240497 44158 240543
rect 41186 240494 41198 240497
rect 44146 240494 44158 240497
rect 44210 240494 44222 240546
rect 343858 196478 343870 196530
rect 343922 196527 343934 196530
rect 344978 196527 344990 196530
rect 343922 196481 344990 196527
rect 343922 196478 343934 196481
rect 344978 196478 344990 196481
rect 345042 196478 345054 196530
rect 310930 160638 310942 160690
rect 310994 160687 311006 160690
rect 311266 160687 311278 160690
rect 310994 160641 311278 160687
rect 310994 160638 311006 160641
rect 311266 160638 311278 160641
rect 311330 160638 311342 160690
<< via1 >>
rect 41134 240494 41186 240546
rect 44158 240494 44210 240546
rect 343870 196478 343922 196530
rect 344990 196478 345042 196530
rect 310942 160638 310994 160690
rect 311278 160638 311330 160690
<< metal2 >>
rect 11032 595672 11256 597000
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 11004 595560 11256 595672
rect 33068 595560 33320 595672
rect 55132 595560 55384 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 143416 595672 143640 597000
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 209608 595672 209832 597000
rect 231672 595672 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 319928 595672 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 99288 595560 99540 595672
rect 4172 388164 4228 388174
rect 4172 333396 4228 388108
rect 4172 333330 4228 333340
rect 11004 301588 11060 595560
rect 12572 573076 12628 573086
rect 12572 395668 12628 573020
rect 14252 530740 14308 530750
rect 14252 397348 14308 530684
rect 14252 397282 14308 397292
rect 15932 488404 15988 488414
rect 12572 395602 12628 395612
rect 15932 393988 15988 488348
rect 15932 393922 15988 393932
rect 33068 392308 33124 595560
rect 55132 409220 55188 595560
rect 77308 572068 77364 595560
rect 99484 590548 99540 595560
rect 99484 590482 99540 590492
rect 121324 595560 121576 595672
rect 143388 595560 143640 595672
rect 165452 595560 165704 595672
rect 187516 595560 187768 595672
rect 209580 595560 209832 595672
rect 231644 595560 231896 595672
rect 253708 595560 253960 595672
rect 275772 595560 276024 595672
rect 297836 595560 298088 595672
rect 319900 595560 320152 595672
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386120 595672 386344 597000
rect 386120 595560 386372 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 430220 595560 430472 595672
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 452312 595560 452564 595672
rect 77308 572002 77364 572012
rect 121324 570388 121380 595560
rect 121324 570322 121380 570332
rect 141932 590548 141988 590558
rect 57932 544852 57988 544862
rect 56252 502516 56308 502526
rect 56252 409892 56308 502460
rect 56252 409826 56308 409836
rect 57932 409780 57988 544796
rect 57932 409714 57988 409724
rect 55132 409154 55188 409164
rect 33068 392242 33124 392252
rect 103404 407428 103460 407438
rect 99932 386708 99988 386718
rect 38556 386596 38612 386606
rect 38444 386484 38500 386494
rect 11004 301522 11060 301532
rect 12572 383124 12628 383134
rect 4172 290836 4228 290846
rect 4172 239428 4228 290780
rect 12572 276724 12628 383068
rect 32732 380212 32788 380222
rect 29372 380100 29428 380110
rect 27692 379988 27748 379998
rect 20972 379876 21028 379886
rect 12572 276658 12628 276668
rect 14252 379316 14308 379326
rect 4172 239362 4228 239372
rect 13244 229460 13300 229470
rect 4172 208740 4228 208750
rect 4172 121716 4228 208684
rect 4172 121650 4228 121660
rect 11340 47908 11396 47918
rect 11340 480 11396 47852
rect 13244 480 13300 229404
rect 14252 192052 14308 379260
rect 14252 191986 14308 191996
rect 20860 229348 20916 229358
rect 14252 79156 14308 79166
rect 14252 50372 14308 79100
rect 14252 50306 14308 50316
rect 15372 4228 15428 4238
rect 15372 480 15428 4172
rect 17276 4228 17332 4238
rect 17276 480 17332 4172
rect 19180 4228 19236 4238
rect 19180 480 19236 4172
rect 11340 392 11592 480
rect 13244 392 13496 480
rect 11368 -960 11592 392
rect 13272 -960 13496 392
rect 15176 392 15428 480
rect 17080 392 17332 480
rect 18984 392 19236 480
rect 20860 480 20916 229292
rect 20972 65044 21028 379820
rect 20972 64978 21028 64988
rect 22764 232708 22820 232718
rect 22764 480 22820 232652
rect 26572 222628 26628 222638
rect 25116 4228 25172 4238
rect 24892 4172 25116 4228
rect 24892 480 24948 4172
rect 25116 4162 25172 4172
rect 20860 392 21112 480
rect 22764 392 23016 480
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 24696 392 24948 480
rect 26572 480 26628 222572
rect 27692 22708 27748 379932
rect 29372 107380 29428 380044
rect 29372 107314 29428 107324
rect 30380 227668 30436 227678
rect 27692 22642 27748 22652
rect 30380 480 30436 227612
rect 32284 214228 32340 214238
rect 32284 480 32340 214172
rect 32732 149716 32788 380156
rect 38332 379540 38388 379550
rect 38332 238196 38388 379484
rect 38444 238308 38500 386428
rect 38556 238532 38612 386540
rect 40908 384020 40964 384030
rect 40684 379428 40740 379438
rect 38556 238466 38612 238476
rect 40236 378644 40292 378654
rect 40236 238420 40292 378588
rect 40236 238354 40292 238364
rect 38444 238242 38500 238252
rect 38332 238130 38388 238140
rect 40684 237972 40740 379372
rect 40908 243628 40964 383964
rect 41132 380772 41188 380782
rect 41132 255388 41188 380716
rect 62412 304052 62468 304062
rect 47404 302484 47460 302494
rect 47404 299880 47460 302428
rect 62412 299880 62468 303996
rect 77420 304052 77476 304062
rect 77420 299880 77476 303996
rect 92428 304052 92484 304062
rect 92428 299880 92484 303996
rect 41132 255332 41748 255388
rect 40908 243572 41188 243628
rect 41132 240546 41188 243572
rect 41132 240494 41134 240546
rect 41186 240494 41188 240546
rect 41132 240482 41188 240494
rect 41692 240548 41748 255332
rect 60844 240772 60900 240782
rect 60844 240706 60900 240716
rect 74956 240772 75012 240782
rect 74956 240706 75012 240716
rect 44156 240548 44212 240558
rect 64876 240548 64932 240558
rect 41692 240492 42728 240548
rect 44156 240546 44744 240548
rect 44156 240494 44158 240546
rect 44210 240494 44744 240546
rect 44156 240492 44744 240494
rect 44156 240482 44212 240492
rect 64876 240482 64932 240492
rect 62860 240436 62916 240446
rect 62860 240370 62916 240380
rect 66892 240324 66948 240334
rect 66892 240258 66948 240268
rect 68908 240212 68964 240222
rect 68908 240146 68964 240156
rect 56812 240100 56868 240110
rect 46732 238532 46788 240072
rect 46732 238466 46788 238476
rect 48748 238196 48804 240072
rect 50764 238308 50820 240072
rect 52780 238420 52836 240072
rect 52780 238354 52836 238364
rect 50764 238242 50820 238252
rect 48748 238130 48804 238140
rect 40684 237906 40740 237916
rect 54796 237972 54852 240072
rect 56812 240034 56868 240044
rect 58828 239876 58884 240072
rect 58828 239810 58884 239820
rect 54796 237906 54852 237916
rect 70924 235172 70980 240072
rect 72940 238532 72996 240072
rect 72940 238466 72996 238476
rect 76972 238532 77028 240072
rect 76972 238466 77028 238476
rect 78988 237972 79044 240072
rect 81004 239764 81060 240072
rect 81004 239698 81060 239708
rect 78988 237906 79044 237916
rect 83020 237860 83076 240072
rect 85036 238084 85092 240072
rect 87052 238196 87108 240072
rect 87052 238130 87108 238140
rect 85036 238018 85092 238028
rect 83020 237794 83076 237804
rect 89068 237748 89124 240072
rect 91084 238532 91140 240072
rect 91084 238466 91140 238476
rect 93100 238308 93156 240072
rect 95116 238532 95172 240072
rect 95116 238466 95172 238476
rect 97132 238420 97188 240072
rect 99932 238532 99988 386652
rect 103292 385140 103348 385150
rect 100380 385028 100436 385038
rect 99932 238466 99988 238476
rect 100156 384804 100212 384814
rect 97132 238354 97188 238364
rect 93100 238242 93156 238252
rect 89068 237682 89124 237692
rect 96572 238196 96628 238206
rect 96572 237636 96628 238140
rect 100156 237748 100212 384748
rect 100380 237860 100436 384972
rect 103292 237972 103348 385084
rect 103404 284452 103460 407372
rect 141932 390740 141988 590492
rect 143388 410788 143444 595560
rect 143388 410722 143444 410732
rect 165452 392420 165508 595560
rect 186396 590548 186452 590558
rect 179004 587188 179060 587198
rect 175532 572068 175588 572078
rect 172172 570388 172228 570398
rect 172172 408100 172228 570332
rect 172172 408034 172228 408044
rect 173852 446068 173908 446078
rect 173852 399028 173908 446012
rect 173852 398962 173908 398972
rect 165452 392354 165508 392364
rect 141932 390674 141988 390684
rect 111692 386820 111748 386830
rect 103404 284386 103460 284396
rect 103516 384916 103572 384926
rect 103516 238196 103572 384860
rect 106652 383348 106708 383358
rect 104972 379092 105028 379102
rect 103628 286580 103684 286590
rect 103628 272804 103684 286524
rect 103628 272738 103684 272748
rect 103516 238130 103572 238140
rect 103292 237906 103348 237916
rect 100380 237794 100436 237804
rect 100156 237682 100212 237692
rect 96572 237570 96628 237580
rect 104972 237636 105028 379036
rect 106652 238420 106708 383292
rect 106652 238354 106708 238364
rect 111692 238308 111748 386764
rect 118412 383572 118468 383582
rect 115052 382116 115108 382126
rect 113372 321860 113428 321870
rect 113372 278628 113428 321804
rect 113372 278562 113428 278572
rect 115052 239876 115108 382060
rect 115164 320180 115220 320190
rect 115164 261156 115220 320124
rect 115164 261090 115220 261100
rect 115052 239810 115108 239820
rect 111692 238242 111748 238252
rect 118412 238084 118468 383516
rect 126812 381780 126868 381790
rect 120092 381668 120148 381678
rect 120092 239988 120148 381612
rect 120092 239922 120148 239932
rect 125132 381556 125188 381566
rect 125132 239764 125188 381500
rect 125244 378980 125300 378990
rect 125244 319060 125300 378924
rect 125244 318994 125300 319004
rect 126812 241108 126868 381724
rect 126812 241042 126868 241052
rect 130172 380324 130228 380334
rect 125132 239698 125188 239708
rect 118412 238018 118468 238028
rect 104972 237570 105028 237580
rect 70924 235106 70980 235116
rect 130172 234388 130228 380268
rect 130284 378756 130340 378766
rect 130284 361396 130340 378700
rect 130284 361330 130340 361340
rect 140252 322084 140308 322094
rect 140252 266980 140308 322028
rect 168028 322084 168084 322094
rect 152796 321972 152852 321982
rect 143612 321748 143668 321758
rect 143612 302484 143668 321692
rect 143612 289044 143668 302428
rect 143612 285908 143668 288988
rect 151116 288932 151172 288942
rect 151116 287252 151172 288876
rect 151116 287196 151284 287252
rect 143612 285852 144312 285908
rect 151228 285348 151284 287196
rect 152796 285880 152852 321916
rect 168028 321636 168084 322028
rect 168028 321570 168084 321580
rect 173964 301588 174020 301598
rect 161308 299908 161364 299918
rect 161308 285880 161364 299852
rect 169148 289828 169204 289838
rect 168812 286692 168868 286702
rect 151228 285282 151284 285292
rect 165452 285348 165508 285358
rect 165452 278852 165508 285292
rect 165452 278786 165508 278796
rect 168812 277956 168868 286636
rect 169148 284004 169204 289772
rect 169148 283938 169204 283948
rect 168812 277890 168868 277900
rect 173964 273028 174020 301532
rect 174636 278852 174692 278862
rect 174636 276052 174692 278796
rect 174636 275986 174692 275996
rect 173964 272962 174020 272972
rect 175532 271684 175588 572012
rect 178892 414596 178948 414606
rect 177324 410788 177380 410798
rect 176316 360388 176372 360398
rect 175532 271618 175588 271628
rect 175980 337540 176036 337550
rect 140252 266914 140308 266924
rect 174636 268772 174692 268782
rect 174636 267204 174692 268716
rect 174636 239988 174692 267148
rect 174636 239922 174692 239932
rect 130172 234322 130228 234332
rect 175980 233044 176036 337484
rect 175980 232978 176036 232988
rect 176092 333508 176148 333518
rect 40236 229572 40292 229582
rect 38556 224420 38612 224430
rect 37996 222852 38052 222862
rect 32732 149650 32788 149660
rect 33516 210868 33572 210878
rect 33516 4452 33572 210812
rect 33516 4386 33572 4396
rect 34412 4228 34468 4238
rect 34412 480 34468 4172
rect 37996 480 38052 222796
rect 38444 219268 38500 219278
rect 38332 214452 38388 214462
rect 38332 4228 38388 214396
rect 38332 4162 38388 4172
rect 38444 4116 38500 219212
rect 38556 5012 38612 224364
rect 38556 4946 38612 4956
rect 39900 222740 39956 222750
rect 38444 4050 38500 4060
rect 39900 480 39956 222684
rect 40236 4676 40292 229516
rect 176092 221060 176148 333452
rect 176092 220994 176148 221004
rect 176204 329476 176260 329486
rect 176204 217812 176260 329420
rect 176316 220948 176372 360332
rect 176428 346276 176484 346286
rect 176428 286580 176484 346220
rect 176428 286514 176484 286524
rect 177212 276052 177268 276062
rect 177212 265524 177268 275996
rect 177324 270340 177380 410732
rect 177996 357700 178052 357710
rect 177324 270274 177380 270284
rect 177884 338884 177940 338894
rect 177212 265458 177268 265468
rect 177884 234164 177940 338828
rect 177884 234098 177940 234108
rect 177996 224644 178052 357644
rect 178556 342916 178612 342926
rect 178332 336084 178388 336094
rect 178220 332836 178276 332846
rect 178220 249508 178276 332780
rect 178220 249442 178276 249452
rect 178332 255332 178388 336028
rect 178444 330148 178500 330158
rect 178444 255388 178500 330092
rect 178556 321636 178612 342860
rect 178892 321748 178948 414540
rect 179004 409332 179060 587132
rect 184716 578788 184772 578798
rect 179004 409266 179060 409276
rect 180460 577108 180516 577118
rect 179228 403732 179284 403742
rect 179004 390964 179060 390974
rect 179004 342916 179060 390908
rect 179228 390852 179284 403676
rect 179228 390786 179284 390796
rect 179676 362964 179732 362974
rect 179452 356244 179508 356254
rect 179004 342850 179060 342860
rect 179116 354452 179172 354462
rect 179116 336084 179172 354396
rect 179116 336018 179172 336028
rect 178892 321682 178948 321692
rect 178556 321570 178612 321580
rect 178444 255332 179172 255388
rect 178332 243628 178388 255276
rect 179004 249508 179060 249518
rect 178332 243572 178948 243628
rect 178892 224756 178948 243572
rect 178892 224690 178948 224700
rect 177996 224578 178052 224588
rect 179004 222964 179060 249452
rect 179116 243684 179172 255332
rect 179116 231364 179172 243628
rect 179452 232820 179508 356188
rect 179452 232754 179508 232764
rect 179564 350980 179620 350990
rect 179116 231298 179172 231308
rect 179564 223076 179620 350924
rect 179676 234724 179732 362908
rect 180460 262276 180516 577052
rect 183932 460180 183988 460190
rect 181468 417844 181524 417854
rect 181468 409556 181524 417788
rect 181468 409490 181524 409500
rect 183932 409444 183988 460124
rect 183932 409378 183988 409388
rect 182476 407652 182532 407662
rect 180908 397460 180964 397470
rect 180796 395780 180852 395790
rect 180684 385476 180740 385486
rect 180460 262210 180516 262220
rect 180572 380436 180628 380446
rect 180572 235172 180628 380380
rect 180684 240772 180740 385420
rect 180796 322756 180852 395724
rect 180908 346276 180964 397404
rect 182364 394212 182420 394222
rect 182252 379764 182308 379774
rect 182252 379540 182308 379708
rect 182252 379474 182308 379484
rect 182252 369796 182308 369806
rect 181244 361732 181300 361742
rect 181132 352324 181188 352334
rect 180908 346210 180964 346220
rect 181020 349636 181076 349646
rect 180796 322690 180852 322700
rect 180908 344260 180964 344270
rect 180684 240706 180740 240716
rect 180572 235106 180628 235116
rect 179676 234658 179732 234668
rect 180908 232932 180964 344204
rect 181020 234836 181076 349580
rect 181020 234770 181076 234780
rect 180908 232866 180964 232876
rect 181132 229684 181188 352268
rect 181132 229618 181188 229628
rect 181244 227780 181300 361676
rect 182252 299908 182308 369740
rect 182364 330260 182420 394156
rect 182476 354452 182532 407596
rect 184044 394100 184100 394110
rect 183932 385588 183988 385598
rect 182476 354386 182532 354396
rect 183820 368452 183876 368462
rect 183036 353668 183092 353678
rect 182812 348292 182868 348302
rect 182364 330194 182420 330204
rect 182588 334852 182644 334862
rect 182252 299842 182308 299852
rect 181356 272132 181412 272142
rect 181356 240660 181412 272076
rect 181468 265524 181524 265534
rect 181468 255444 181524 265468
rect 181468 255378 181524 255388
rect 181356 240594 181412 240604
rect 182588 239540 182644 334796
rect 182588 239474 182644 239484
rect 182700 330820 182756 330830
rect 182700 229908 182756 330764
rect 182700 229842 182756 229852
rect 182812 227892 182868 348236
rect 182812 227826 182868 227836
rect 182924 341572 182980 341582
rect 181244 227714 181300 227724
rect 179564 223010 179620 223020
rect 179004 222898 179060 222908
rect 176316 220882 176372 220892
rect 176204 217746 176260 217756
rect 154924 217700 154980 217710
rect 40236 4610 40292 4620
rect 41132 215908 41188 215918
rect 41132 4564 41188 215852
rect 154924 209944 154980 217644
rect 182924 217700 182980 341516
rect 183036 219380 183092 353612
rect 183820 322308 183876 368396
rect 183820 322242 183876 322252
rect 183932 240324 183988 385532
rect 184044 332836 184100 394044
rect 184044 332770 184100 332780
rect 184156 380548 184212 380558
rect 184156 240548 184212 380492
rect 184604 365764 184660 365774
rect 184492 345604 184548 345614
rect 184380 332164 184436 332174
rect 184156 240482 184212 240492
rect 184268 328132 184324 328142
rect 183932 240258 183988 240268
rect 183036 219314 183092 219324
rect 184268 217924 184324 328076
rect 184380 219492 184436 332108
rect 184492 224868 184548 345548
rect 184492 224802 184548 224812
rect 184380 219426 184436 219436
rect 184268 217858 184324 217868
rect 182924 217634 182980 217644
rect 184604 209524 184660 365708
rect 184716 263620 184772 578732
rect 186284 565124 186340 565134
rect 186172 550788 186228 550798
rect 186060 543620 186116 543630
rect 186060 388948 186116 543564
rect 186060 388882 186116 388892
rect 186172 387268 186228 550732
rect 186284 390628 186340 565068
rect 186396 404180 186452 590492
rect 187180 514948 187236 514958
rect 187180 408996 187236 514892
rect 187180 408930 187236 408940
rect 187292 507780 187348 507790
rect 186396 404114 186452 404124
rect 186284 390562 186340 390572
rect 186172 387202 186228 387212
rect 186396 359044 186452 359054
rect 186284 346948 186340 346958
rect 186172 340228 186228 340238
rect 185612 283892 185668 283902
rect 185612 278908 185668 283836
rect 185612 278852 185780 278908
rect 184716 263554 184772 263564
rect 185724 273924 185780 278852
rect 185612 255444 185668 255454
rect 185612 243572 185668 255388
rect 185612 243506 185668 243516
rect 185724 240548 185780 273868
rect 185724 240482 185780 240492
rect 186172 228004 186228 340172
rect 186284 231140 186340 346892
rect 186284 231074 186340 231084
rect 186172 227938 186228 227948
rect 186396 223188 186452 358988
rect 186508 296548 186564 296558
rect 186508 286692 186564 296492
rect 187292 289828 187348 507724
rect 187516 487284 187572 595560
rect 189644 591332 189700 591342
rect 189196 590996 189252 591006
rect 189084 575428 189140 575438
rect 187852 557956 187908 557966
rect 187516 487218 187572 487228
rect 187740 536452 187796 536462
rect 187292 289762 187348 289772
rect 187404 471940 187460 471950
rect 186508 286626 186564 286636
rect 187180 285684 187236 285694
rect 187180 280532 187236 285628
rect 187404 283892 187460 471884
rect 187628 464772 187684 464782
rect 187404 283826 187460 283836
rect 187516 450436 187572 450446
rect 187516 281428 187572 450380
rect 187628 283668 187684 464716
rect 187740 409668 187796 536396
rect 187852 410452 187908 557900
rect 188076 493444 188132 493454
rect 187852 410386 187908 410396
rect 187964 443268 188020 443278
rect 187740 409602 187796 409612
rect 187852 295652 187908 295662
rect 187852 285796 187908 295596
rect 187852 285730 187908 285740
rect 187628 283602 187684 283612
rect 187964 282212 188020 443212
rect 188076 288484 188132 493388
rect 188860 487284 188916 487294
rect 188860 407876 188916 487228
rect 189084 407988 189140 575372
rect 189084 407922 189140 407932
rect 188860 407810 188916 407820
rect 189196 407540 189252 590940
rect 189196 407474 189252 407484
rect 189308 590772 189364 590782
rect 189308 405748 189364 590716
rect 189532 572068 189588 572078
rect 189308 405682 189364 405692
rect 189420 570388 189476 570398
rect 189308 367108 189364 367118
rect 189196 355012 189252 355022
rect 189084 342916 189140 342926
rect 188860 336196 188916 336206
rect 188076 288418 188132 288428
rect 188748 326788 188804 326798
rect 187964 282146 188020 282156
rect 187516 281362 187572 281372
rect 187180 280466 187236 280476
rect 188188 243572 188244 243582
rect 188076 242116 188132 242126
rect 188076 236292 188132 242060
rect 188188 238532 188244 243516
rect 188188 238466 188244 238476
rect 188076 236226 188132 236236
rect 188748 233156 188804 326732
rect 188748 233090 188804 233100
rect 188860 231252 188916 336140
rect 188860 231186 188916 231196
rect 189084 229796 189140 342860
rect 189196 231028 189252 354956
rect 189196 230962 189252 230972
rect 189084 229730 189140 229740
rect 186396 223122 186452 223132
rect 189308 212660 189364 367052
rect 189420 266308 189476 570332
rect 189532 267652 189588 572012
rect 189644 268996 189700 591276
rect 209580 591332 209636 595560
rect 209580 591266 209636 591276
rect 190652 591220 190708 591230
rect 189644 268930 189700 268940
rect 189756 588868 189812 588878
rect 189532 267586 189588 267596
rect 189420 266242 189476 266252
rect 189756 264964 189812 588812
rect 190652 399140 190708 591164
rect 231644 591220 231700 595560
rect 231644 591154 231700 591164
rect 253708 591108 253764 595560
rect 253708 591042 253764 591052
rect 275772 572068 275828 595560
rect 297836 590996 297892 595560
rect 297836 590930 297892 590940
rect 319900 590884 319956 595560
rect 319900 590818 319956 590828
rect 275772 572002 275828 572012
rect 341964 570388 342020 595560
rect 364028 590772 364084 595560
rect 364028 590706 364084 590716
rect 386316 590772 386372 595560
rect 386316 590706 386372 590716
rect 401436 590772 401492 590782
rect 401436 587972 401492 590716
rect 408268 588868 408324 595560
rect 430220 590660 430276 595560
rect 430220 590594 430276 590604
rect 452508 590660 452564 595560
rect 452508 590594 452564 590604
rect 474348 595560 474600 595672
rect 496412 595560 496664 595672
rect 518476 595560 518728 595672
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 408268 588802 408324 588812
rect 401436 587906 401492 587916
rect 407372 587972 407428 587982
rect 341964 570322 342020 570332
rect 407372 567028 407428 587916
rect 474348 578788 474404 595560
rect 496412 590548 496468 595560
rect 496412 590482 496468 590492
rect 518476 590212 518532 595560
rect 518476 590146 518532 590156
rect 474348 578722 474404 578732
rect 540540 577108 540596 595560
rect 562604 591332 562660 595560
rect 562604 591266 562660 591276
rect 584668 590212 584724 595560
rect 584668 590146 584724 590156
rect 540540 577042 540596 577052
rect 407372 566962 407428 566972
rect 552748 560420 552804 560430
rect 551068 541604 551124 541614
rect 549948 507892 550004 507902
rect 549500 484484 549556 484494
rect 549388 423444 549444 423454
rect 341404 410452 341460 410462
rect 190652 399074 190708 399084
rect 195132 394212 195188 410088
rect 195132 394146 195188 394156
rect 200508 394100 200564 410088
rect 205884 407652 205940 410088
rect 205884 407586 205940 407596
rect 208348 407988 208404 407998
rect 204764 404068 204820 404078
rect 200508 394034 200564 394044
rect 202860 394772 202916 394782
rect 201964 393204 202020 393214
rect 197372 382228 197428 382238
rect 196476 382004 196532 382014
rect 190652 380660 190708 380670
rect 189756 264898 189812 264908
rect 190092 292628 190148 292638
rect 189308 212594 189364 212604
rect 190092 211316 190148 292572
rect 190652 250348 190708 380604
rect 196476 379988 196532 381948
rect 197372 379988 197428 382172
rect 199164 382228 199220 382238
rect 198044 382004 198100 382014
rect 198044 379988 198100 381948
rect 199164 379988 199220 382172
rect 200844 382228 200900 382238
rect 199724 382004 199780 382014
rect 199724 379988 199780 381948
rect 200844 379988 200900 382172
rect 201404 382004 201460 382014
rect 201404 379988 201460 381948
rect 195832 379932 196532 379988
rect 196728 379932 197428 379988
rect 197624 379932 198100 379988
rect 198520 379932 199220 379988
rect 199416 379932 199780 379988
rect 200312 379932 200900 379988
rect 201208 379932 201460 379988
rect 201964 379988 202020 393148
rect 202860 379988 202916 394716
rect 204764 384748 204820 404012
rect 206556 402500 206612 402510
rect 206556 384748 206612 402444
rect 208348 396508 208404 407932
rect 211036 405860 211092 405870
rect 210140 404180 210196 404190
rect 208348 396452 208516 396508
rect 204652 384692 204820 384748
rect 206444 384692 206612 384748
rect 204316 382004 204372 382014
rect 204316 379988 204372 381948
rect 201964 379932 202104 379988
rect 202860 379932 203000 379988
rect 203896 379932 204372 379988
rect 204652 379988 204708 384692
rect 206108 382004 206164 382014
rect 206108 379988 206164 381948
rect 204652 379932 204792 379988
rect 205688 379932 206164 379988
rect 206444 379988 206500 384692
rect 208236 382228 208292 382238
rect 208236 379988 208292 382172
rect 208460 379988 208516 396452
rect 210140 384748 210196 404124
rect 210028 384692 210196 384748
rect 210364 399812 210420 399822
rect 210364 398244 210420 399756
rect 209916 382228 209972 382238
rect 209916 379988 209972 382172
rect 206444 379932 206584 379988
rect 207480 379932 208292 379988
rect 208376 379932 208516 379988
rect 209272 379932 209972 379988
rect 210028 379988 210084 384692
rect 210028 379932 210168 379988
rect 210364 379764 210420 398188
rect 211036 384748 211092 405804
rect 211260 399812 211316 410088
rect 212828 407540 212884 407550
rect 211260 399746 211316 399756
rect 211932 405748 211988 405758
rect 211932 384748 211988 405692
rect 212828 384748 212884 407484
rect 213724 399140 213780 399150
rect 213724 384748 213780 399084
rect 210924 384692 211092 384748
rect 211820 384692 211988 384748
rect 212716 384692 212884 384748
rect 213612 384692 213780 384748
rect 214508 392420 214564 392430
rect 210924 379988 210980 384692
rect 211820 379988 211876 384692
rect 212716 379988 212772 384692
rect 213612 379988 213668 384692
rect 214508 379988 214564 392364
rect 216300 392308 216356 392318
rect 215404 390740 215460 390750
rect 215404 379988 215460 390684
rect 216300 379988 216356 392252
rect 216636 391412 216692 410088
rect 222012 403284 222068 410088
rect 227416 410060 227668 410116
rect 227612 406644 227668 410060
rect 232764 407428 232820 410088
rect 232764 407362 232820 407372
rect 238140 407092 238196 410088
rect 243516 407988 243572 410088
rect 243516 407922 243572 407932
rect 248892 407540 248948 410088
rect 254268 407988 254324 410088
rect 254268 407922 254324 407932
rect 259644 407652 259700 410088
rect 259644 407586 259700 407596
rect 248892 407474 248948 407484
rect 238140 407026 238196 407036
rect 227612 406578 227668 406588
rect 265020 406644 265076 410088
rect 265020 406578 265076 406588
rect 270396 409108 270452 410088
rect 275800 410060 276388 410116
rect 281176 410060 281428 410116
rect 270396 406644 270452 409052
rect 276332 407764 276388 410060
rect 270396 406578 270452 406588
rect 275548 407540 275604 407550
rect 219996 399028 220052 399038
rect 218204 397348 218260 397358
rect 216636 391346 216692 391356
rect 217196 395668 217252 395678
rect 217196 379988 217252 395612
rect 218204 384748 218260 397292
rect 218092 384692 218260 384748
rect 218988 393988 219044 393998
rect 218092 379988 218148 384692
rect 218988 379988 219044 393932
rect 219996 384748 220052 398972
rect 222012 397460 222068 403228
rect 222012 397394 222068 397404
rect 275548 396508 275604 407484
rect 276332 406644 276388 407708
rect 276332 406578 276388 406588
rect 280028 409108 280084 409118
rect 278236 400708 278292 400718
rect 275548 396452 275716 396508
rect 219884 384692 220052 384748
rect 220780 390852 220836 390862
rect 219884 379988 219940 384692
rect 220780 379988 220836 390796
rect 272188 386820 272244 386830
rect 252028 386596 252084 386606
rect 246764 385364 246820 385374
rect 240716 383684 240772 383694
rect 245196 383684 245252 383694
rect 240772 383628 240884 383684
rect 240716 383618 240772 383628
rect 235116 383236 235172 383246
rect 223468 383124 223524 383134
rect 223468 379988 223524 383068
rect 231644 382340 231700 382350
rect 231532 382284 231644 382340
rect 230076 382228 230132 382238
rect 223692 380324 223748 380334
rect 223748 380268 223860 380324
rect 223692 380258 223748 380268
rect 223804 379988 223860 380268
rect 225484 380212 225540 380222
rect 225540 380156 225652 380212
rect 225484 380146 225540 380156
rect 225596 379988 225652 380156
rect 226828 380100 226884 380110
rect 226828 379988 226884 380044
rect 228956 379988 229012 379998
rect 230076 379988 230132 382172
rect 231532 379988 231588 382284
rect 231644 382274 231700 382284
rect 231756 382228 231812 382238
rect 231756 379988 231812 382172
rect 210924 379932 211064 379988
rect 211820 379932 211960 379988
rect 212716 379932 212856 379988
rect 213612 379932 213752 379988
rect 214508 379932 214648 379988
rect 215404 379932 215544 379988
rect 216300 379932 216440 379988
rect 217196 379932 217336 379988
rect 218092 379932 218232 379988
rect 218988 379932 219128 379988
rect 219884 379932 220024 379988
rect 220780 379932 220920 379988
rect 223468 379932 223608 379988
rect 223804 379932 224504 379988
rect 225596 379932 226296 379988
rect 226828 379932 227192 379988
rect 229880 379932 230132 379988
rect 230776 379932 231588 379988
rect 231672 379932 231812 379988
rect 232204 382004 232260 382014
rect 232204 379988 232260 381948
rect 232652 381892 232708 381902
rect 232708 381836 232820 381892
rect 232652 381826 232708 381836
rect 232764 379988 232820 381836
rect 235116 379988 235172 383180
rect 240156 381892 240212 381902
rect 239484 381444 239540 381454
rect 239484 379988 239540 381388
rect 240156 379988 240212 381836
rect 232204 379932 232568 379988
rect 232764 379932 233464 379988
rect 234360 379932 235172 379988
rect 238840 379932 239540 379988
rect 239736 379932 240212 379988
rect 240828 379988 240884 383628
rect 244972 383124 245028 383134
rect 244972 379988 245028 383068
rect 245196 379988 245252 383628
rect 246652 380212 246708 380222
rect 246652 379988 246708 380156
rect 240828 379932 241528 379988
rect 244216 379932 245028 379988
rect 245112 379932 245252 379988
rect 246008 379932 246708 379988
rect 246764 379988 246820 385308
rect 250572 384020 250628 384030
rect 250628 383964 250740 384020
rect 250572 383954 250628 383964
rect 250348 380772 250404 380782
rect 248556 380100 248612 380110
rect 248556 379988 248612 380044
rect 246764 379932 246904 379988
rect 247800 379932 248612 379988
rect 248668 379988 248724 379998
rect 250348 379988 250404 380716
rect 250684 379988 250740 383964
rect 252028 379988 252084 386540
rect 253708 386484 253764 386494
rect 253708 379988 253764 386428
rect 260540 385588 260596 385598
rect 257068 382116 257124 382126
rect 256060 381668 256116 381678
rect 256060 379988 256116 381612
rect 257068 379988 257124 382060
rect 257740 381780 257796 381790
rect 257796 381724 257908 381780
rect 257740 381714 257796 381724
rect 257852 379988 257908 381724
rect 258748 380660 258804 380670
rect 258748 379988 258804 380604
rect 259532 380548 259588 380558
rect 259588 380492 259700 380548
rect 259532 380482 259588 380492
rect 259644 379988 259700 380492
rect 260540 379988 260596 385532
rect 264124 385476 264180 385486
rect 262108 383796 262164 383806
rect 262164 383740 262276 383796
rect 262108 383730 262164 383740
rect 262220 379988 262276 383740
rect 263788 383460 263844 383470
rect 250348 379932 250488 379988
rect 250684 379932 251384 379988
rect 252028 379932 252280 379988
rect 253708 379932 254072 379988
rect 256060 379932 256760 379988
rect 257068 379932 257656 379988
rect 257852 379932 258552 379988
rect 258748 379932 259448 379988
rect 259644 379932 260344 379988
rect 260540 379932 261240 379988
rect 262136 379932 262276 379988
rect 262332 380436 262388 380446
rect 262332 379988 262388 380380
rect 263788 379988 263844 383404
rect 264124 379988 264180 385420
rect 265468 385252 265524 385262
rect 265468 379988 265524 385196
rect 265916 385140 265972 385150
rect 265916 379988 265972 385084
rect 267708 385028 267764 385038
rect 267260 381556 267316 381566
rect 267260 379988 267316 381500
rect 267708 379988 267764 384972
rect 271292 384916 271348 384926
rect 270732 384804 270788 384814
rect 268828 383572 268884 383582
rect 268828 379988 268884 383516
rect 270732 379988 270788 384748
rect 271292 379988 271348 384860
rect 272188 379988 272244 386764
rect 273084 386708 273140 386718
rect 273084 379988 273140 386652
rect 273868 383348 273924 383358
rect 273924 383292 274036 383348
rect 273868 383282 273924 383292
rect 273980 379988 274036 383292
rect 275660 379988 275716 396452
rect 277228 394548 277284 394558
rect 277116 382116 277172 382126
rect 277116 379988 277172 382060
rect 262332 379932 263032 379988
rect 263788 379932 263928 379988
rect 264124 379932 264824 379988
rect 265468 379932 265720 379988
rect 265916 379932 266616 379988
rect 267260 379932 267512 379988
rect 267708 379932 268408 379988
rect 268828 379932 269304 379988
rect 270732 379932 271096 379988
rect 271292 379932 271992 379988
rect 272188 379932 272888 379988
rect 273084 379932 273784 379988
rect 273980 379932 274680 379988
rect 275576 379932 275716 379988
rect 276472 379932 277172 379988
rect 277228 379988 277284 394492
rect 278236 384748 278292 400652
rect 278124 384692 278292 384748
rect 279020 392308 279076 392318
rect 278124 379988 278180 384692
rect 279020 379988 279076 392252
rect 280028 384748 280084 409052
rect 281372 407876 281428 410060
rect 286412 410060 286552 410116
rect 291452 410060 291928 410116
rect 296492 410060 297304 410116
rect 302680 410088 303268 410116
rect 308056 410088 308308 410116
rect 302652 410060 303268 410088
rect 285516 409220 285572 409230
rect 285516 408212 285572 409164
rect 285516 408146 285572 408156
rect 281372 406644 281428 407820
rect 281372 406578 281428 406588
rect 286412 408100 286468 410060
rect 286412 406644 286468 408044
rect 286412 406578 286468 406588
rect 291452 408212 291508 410060
rect 288988 406196 289044 406206
rect 288204 406084 288260 406094
rect 285404 405972 285460 405982
rect 281820 405860 281876 405870
rect 280924 397348 280980 397358
rect 280924 384748 280980 397292
rect 281820 384748 281876 405804
rect 283612 405748 283668 405758
rect 279916 384692 280084 384748
rect 280812 384692 280980 384748
rect 281708 384692 281876 384748
rect 282604 390740 282660 390750
rect 279916 379988 279972 384692
rect 280812 379988 280868 384692
rect 281708 379988 281764 384692
rect 282604 379988 282660 390684
rect 283612 384748 283668 405692
rect 284508 401380 284564 401390
rect 284508 384748 284564 401324
rect 285404 384748 285460 405916
rect 287980 390852 288036 390862
rect 283500 384692 283668 384748
rect 284396 384692 284564 384748
rect 285292 384692 285460 384748
rect 286972 385588 287028 385598
rect 283500 379988 283556 384692
rect 284396 379988 284452 384692
rect 285292 379988 285348 384692
rect 286972 379988 287028 385532
rect 287196 382116 287252 382126
rect 277228 379932 277368 379988
rect 278124 379932 278264 379988
rect 279020 379932 279160 379988
rect 279916 379932 280056 379988
rect 280812 379932 280952 379988
rect 281708 379932 281848 379988
rect 282604 379932 282744 379988
rect 283500 379932 283640 379988
rect 284396 379932 284536 379988
rect 285292 379932 285432 379988
rect 286328 379932 287028 379988
rect 287084 382060 287196 382116
rect 287084 379988 287140 382060
rect 287196 382050 287252 382060
rect 287980 379988 288036 390796
rect 288204 382116 288260 406028
rect 288988 396508 289044 406140
rect 288988 396452 289156 396508
rect 288204 382050 288260 382060
rect 289100 379988 289156 396452
rect 290668 395668 290724 395678
rect 290556 385700 290612 385710
rect 290556 379988 290612 385644
rect 287084 379932 287224 379988
rect 287980 379932 288120 379988
rect 289016 379932 289156 379988
rect 289912 379932 290612 379988
rect 290668 379988 290724 395612
rect 291452 380548 291508 408156
rect 293468 410004 293524 410014
rect 292572 400820 292628 400830
rect 291676 397460 291732 397470
rect 291676 384748 291732 397404
rect 292572 384748 292628 400764
rect 293468 384748 293524 409948
rect 296492 409332 296548 410060
rect 302652 409780 302708 410060
rect 302652 409714 302708 409724
rect 294364 409220 294420 409230
rect 294364 384748 294420 409164
rect 295260 402836 295316 402846
rect 295260 384748 295316 402780
rect 296156 399028 296212 399038
rect 296156 384748 296212 398972
rect 296492 385812 296548 409276
rect 298844 408660 298900 408670
rect 296492 385746 296548 385756
rect 297052 404628 297108 404638
rect 297052 384748 297108 404572
rect 297948 399140 298004 399150
rect 297948 384748 298004 399084
rect 298844 384748 298900 408604
rect 300636 404516 300692 404526
rect 299740 399252 299796 399262
rect 299740 384748 299796 399196
rect 300636 384748 300692 404460
rect 302428 399588 302484 399598
rect 301532 399364 301588 399374
rect 301532 384748 301588 399308
rect 302428 396508 302484 399532
rect 302428 396452 302596 396508
rect 291452 380482 291508 380492
rect 291564 384692 291732 384748
rect 292460 384692 292628 384748
rect 293356 384692 293524 384748
rect 294252 384692 294420 384748
rect 295148 384692 295316 384748
rect 296044 384692 296212 384748
rect 296940 384692 297108 384748
rect 297836 384692 298004 384748
rect 298732 384692 298900 384748
rect 299628 384692 299796 384748
rect 300524 384692 300692 384748
rect 301420 384692 301588 384748
rect 291564 379988 291620 384692
rect 292460 379988 292516 384692
rect 293356 379988 293412 384692
rect 294252 379988 294308 384692
rect 295148 379988 295204 384692
rect 296044 379988 296100 384692
rect 296940 379988 296996 384692
rect 297836 379988 297892 384692
rect 298732 379988 298788 384692
rect 299628 379988 299684 384692
rect 300524 379988 300580 384692
rect 301420 379988 301476 384692
rect 302540 379988 302596 396452
rect 303212 385924 303268 410060
rect 308028 410060 308308 410088
rect 308028 409892 308084 410060
rect 308028 409826 308084 409836
rect 304220 408548 304276 408558
rect 303324 399476 303380 399486
rect 303324 396508 303380 399420
rect 303324 396452 303492 396508
rect 303212 385858 303268 385868
rect 303436 379988 303492 396452
rect 304220 384748 304276 408492
rect 307804 404292 307860 404302
rect 306012 402724 306068 402734
rect 306012 384748 306068 402668
rect 307804 384748 307860 404236
rect 308252 386036 308308 410060
rect 313404 409444 313460 410088
rect 313404 408268 313460 409388
rect 313292 408212 313460 408268
rect 318332 409556 318388 409566
rect 309596 406420 309652 406430
rect 308252 385970 308308 385980
rect 308700 400932 308756 400942
rect 308700 384748 308756 400876
rect 309596 384748 309652 406364
rect 311388 406308 311444 406318
rect 310492 401044 310548 401054
rect 310492 384748 310548 400988
rect 311388 384748 311444 406252
rect 312284 401268 312340 401278
rect 312284 384748 312340 401212
rect 290668 379932 290808 379988
rect 291564 379932 291704 379988
rect 292460 379932 292600 379988
rect 293356 379932 293496 379988
rect 294252 379932 294392 379988
rect 295148 379932 295288 379988
rect 296044 379932 296184 379988
rect 296940 379932 297080 379988
rect 297836 379932 297976 379988
rect 298732 379932 298872 379988
rect 299628 379932 299768 379988
rect 300524 379932 300664 379988
rect 301420 379932 301560 379988
rect 302456 379932 302596 379988
rect 303352 379932 303492 379988
rect 304108 384692 304276 384748
rect 305900 384692 306068 384748
rect 307692 384692 307860 384748
rect 308588 384692 308756 384748
rect 309484 384692 309652 384748
rect 310380 384692 310548 384748
rect 311276 384692 311444 384748
rect 312172 384692 312340 384748
rect 313068 394660 313124 394670
rect 304108 379988 304164 384692
rect 305676 382116 305732 382126
rect 305676 379988 305732 382060
rect 304108 379932 304248 379988
rect 305144 379932 305732 379988
rect 305900 379988 305956 384692
rect 307356 382116 307412 382126
rect 307356 379988 307412 382060
rect 305900 379932 306040 379988
rect 306936 379932 307412 379988
rect 307692 379988 307748 384692
rect 308588 379988 308644 384692
rect 309484 379988 309540 384692
rect 310380 379988 310436 384692
rect 311276 379988 311332 384692
rect 312172 379988 312228 384692
rect 313068 379988 313124 394604
rect 313292 380660 313348 408212
rect 315756 407652 315812 407662
rect 315756 404404 315812 407596
rect 315756 404338 315812 404348
rect 315868 404180 315924 404190
rect 314076 401156 314132 401166
rect 314076 384748 314132 401100
rect 315868 396508 315924 404124
rect 315868 396452 316036 396508
rect 313292 380594 313348 380604
rect 313964 384692 314132 384748
rect 314860 396340 314916 396350
rect 313964 379988 314020 384692
rect 314860 379988 314916 396284
rect 315980 379988 316036 396452
rect 307692 379932 307832 379988
rect 308588 379932 308728 379988
rect 309484 379932 309624 379988
rect 310380 379932 310520 379988
rect 311276 379932 311416 379988
rect 312172 379932 312312 379988
rect 313068 379932 313208 379988
rect 313964 379932 314104 379988
rect 314860 379932 315000 379988
rect 315896 379932 316036 379988
rect 316652 396228 316708 396238
rect 316652 379988 316708 396172
rect 318332 386148 318388 409500
rect 318780 409556 318836 410088
rect 318780 409490 318836 409500
rect 321244 409332 321300 409342
rect 318332 386082 318388 386092
rect 318444 396116 318500 396126
rect 318332 382116 318388 382126
rect 318332 379988 318388 382060
rect 316652 379932 316792 379988
rect 317688 379932 318388 379988
rect 318444 379988 318500 396060
rect 320236 396004 320292 396014
rect 320124 382116 320180 382126
rect 320124 379988 320180 382060
rect 318444 379932 318584 379988
rect 319480 379932 320180 379988
rect 320236 379988 320292 395948
rect 321244 384748 321300 409276
rect 324156 406644 324212 410088
rect 324156 406578 324212 406588
rect 324828 409556 324884 409566
rect 321132 384692 321300 384748
rect 322028 395892 322084 395902
rect 321132 379988 321188 384692
rect 322028 379988 322084 395836
rect 323820 394436 323876 394446
rect 323596 382116 323652 382126
rect 323596 379988 323652 382060
rect 320236 379932 320376 379988
rect 321132 379932 321272 379988
rect 322028 379932 322168 379988
rect 323064 379932 323652 379988
rect 323820 379988 323876 394380
rect 324828 384748 324884 409500
rect 326620 409444 326676 409454
rect 324716 384692 324884 384748
rect 325612 395780 325668 395790
rect 324716 379988 324772 384692
rect 325612 379988 325668 395724
rect 326620 384748 326676 409388
rect 329420 392644 329476 392654
rect 326508 384692 326676 384748
rect 327404 392420 327460 392430
rect 326508 379988 326564 384692
rect 327404 379988 327460 392364
rect 329196 382116 329252 382126
rect 329196 379988 329252 382060
rect 329420 379988 329476 392588
rect 329532 388164 329588 410088
rect 334908 406644 334964 410088
rect 334908 406578 334964 406588
rect 340172 408324 340228 408334
rect 332892 402948 332948 402958
rect 329532 388098 329588 388108
rect 330988 390964 331044 390974
rect 330876 382116 330932 382126
rect 330876 379988 330932 382060
rect 323820 379932 323960 379988
rect 324716 379932 324856 379988
rect 325612 379932 325752 379988
rect 326508 379932 326648 379988
rect 327404 379932 327544 379988
rect 328440 379932 329252 379988
rect 329336 379932 329476 379988
rect 330232 379932 330932 379988
rect 330988 379988 331044 390908
rect 332892 384748 332948 402892
rect 332780 384692 332948 384748
rect 340060 388836 340116 388846
rect 332556 382228 332612 382238
rect 332556 379988 332612 382172
rect 330988 379932 331128 379988
rect 332024 379932 332612 379988
rect 332780 379988 332836 384692
rect 339500 383684 339556 383694
rect 334236 382116 334292 382126
rect 334236 379988 334292 382060
rect 335468 381556 335524 381566
rect 335468 379988 335524 381500
rect 332780 379932 332920 379988
rect 333816 379932 334292 379988
rect 334712 379932 335524 379988
rect 228956 379922 229012 379932
rect 248668 379922 248724 379932
rect 228060 379876 228116 379886
rect 228060 379810 228116 379820
rect 240604 379876 240660 379886
rect 240604 379810 240660 379820
rect 210364 379698 210420 379708
rect 236124 379764 236180 379774
rect 236124 379698 236180 379708
rect 242396 379764 242452 379774
rect 242396 379698 242452 379708
rect 253148 379540 253204 379550
rect 253148 379474 253204 379484
rect 254940 379540 254996 379550
rect 254940 379474 254996 379484
rect 195468 379428 195524 379438
rect 194936 379372 195468 379428
rect 195468 379362 195524 379372
rect 221788 379428 221844 379438
rect 221788 379362 221844 379372
rect 222684 379428 222740 379438
rect 222684 379362 222740 379372
rect 225372 379428 225428 379438
rect 225372 379362 225428 379372
rect 235228 379428 235284 379438
rect 235228 379362 235284 379372
rect 237020 379428 237076 379438
rect 238476 379428 238532 379438
rect 237944 379372 238476 379428
rect 237020 379362 237076 379372
rect 238476 379362 238532 379372
rect 243292 379428 243348 379438
rect 249900 379428 249956 379438
rect 249592 379372 249900 379428
rect 243292 379362 243348 379372
rect 249900 379362 249956 379372
rect 255836 379428 255892 379438
rect 255836 379362 255892 379372
rect 270172 379428 270228 379438
rect 270172 379362 270228 379372
rect 339388 354564 339444 354574
rect 339276 261492 339332 261502
rect 339276 260036 339332 261436
rect 339276 259970 339332 259980
rect 190540 250292 190708 250348
rect 190540 240436 190596 250292
rect 190652 245476 190708 245486
rect 190652 241108 190708 245420
rect 190652 241042 190708 241052
rect 339276 243572 339332 243582
rect 190540 240370 190596 240380
rect 315644 240660 315700 240670
rect 315644 240436 315700 240604
rect 317884 240660 317940 240670
rect 317884 240594 317940 240604
rect 318556 240660 318612 240670
rect 318556 240594 318612 240604
rect 322588 240660 322644 240670
rect 322588 240594 322644 240604
rect 323260 240660 323316 240670
rect 323260 240594 323316 240604
rect 337148 240660 337204 240670
rect 315644 240370 315700 240380
rect 336028 240324 336084 240334
rect 317212 240212 317268 240222
rect 317212 240146 317268 240156
rect 320572 240212 320628 240222
rect 320572 240146 320628 240156
rect 214396 240100 214452 240110
rect 303100 240100 303156 240110
rect 206332 238532 206388 240072
rect 206332 234388 206388 238476
rect 206332 234322 206388 234332
rect 207004 229460 207060 240072
rect 207676 232708 207732 240072
rect 207676 232642 207732 232652
rect 207004 229394 207060 229404
rect 208348 227668 208404 240072
rect 208348 227602 208404 227612
rect 209020 222852 209076 240072
rect 209692 224420 209748 240072
rect 210364 236180 210420 240072
rect 210364 236114 210420 236124
rect 209692 224354 209748 224364
rect 209020 222786 209076 222796
rect 211036 219268 211092 240072
rect 211036 219202 211092 219212
rect 190092 211250 190148 211260
rect 211708 210868 211764 240072
rect 212380 229572 212436 240072
rect 212380 229506 212436 229516
rect 213052 217588 213108 240072
rect 213724 224532 213780 240072
rect 214396 240034 214452 240044
rect 215068 234612 215124 240072
rect 215068 234546 215124 234556
rect 215740 234500 215796 240072
rect 215740 234434 215796 234444
rect 216412 234500 216468 240072
rect 217084 234612 217140 240072
rect 217784 240044 218372 240100
rect 218316 236964 218372 240044
rect 218428 237076 218484 240072
rect 218428 237010 218484 237020
rect 218316 236898 218372 236908
rect 217084 234546 217140 234556
rect 216412 234434 216468 234444
rect 219100 231476 219156 240072
rect 219772 231700 219828 240072
rect 219772 231634 219828 231644
rect 220444 231588 220500 240072
rect 220444 231522 220500 231532
rect 219100 231410 219156 231420
rect 221116 228116 221172 240072
rect 221116 228050 221172 228060
rect 221788 227668 221844 240072
rect 222460 228228 222516 240072
rect 222460 228162 222516 228172
rect 221788 227602 221844 227612
rect 213724 224466 213780 224476
rect 223132 224420 223188 240072
rect 223804 235060 223860 240072
rect 223804 234994 223860 235004
rect 224476 224980 224532 240072
rect 225148 235172 225204 240072
rect 225148 235106 225204 235116
rect 225820 234276 225876 240072
rect 225820 234210 225876 234220
rect 226492 230916 226548 240072
rect 227164 231812 227220 240072
rect 227836 236516 227892 240072
rect 227836 236450 227892 236460
rect 227164 231746 227220 231756
rect 226492 230850 226548 230860
rect 228508 228340 228564 240072
rect 229180 236964 229236 240072
rect 229180 236898 229236 236908
rect 228508 228274 228564 228284
rect 224476 224914 224532 224924
rect 223132 224354 223188 224364
rect 213052 217522 213108 217532
rect 229852 214228 229908 240072
rect 230524 222740 230580 240072
rect 230524 222674 230580 222684
rect 231196 214452 231252 240072
rect 231196 214386 231252 214396
rect 231868 214340 231924 240072
rect 231868 214274 231924 214284
rect 229852 214162 229908 214172
rect 232540 212548 232596 240072
rect 233212 237300 233268 240072
rect 233212 237234 233268 237244
rect 233884 215908 233940 240072
rect 234556 216020 234612 240072
rect 235228 224308 235284 240072
rect 235900 237300 235956 240072
rect 236600 240044 236852 240100
rect 235900 237234 235956 237244
rect 236796 236964 236852 240044
rect 236796 236898 236852 236908
rect 237244 228452 237300 240072
rect 237244 228386 237300 228396
rect 237916 227556 237972 240072
rect 237916 227490 237972 227500
rect 235228 224242 235284 224252
rect 234556 215954 234612 215964
rect 233884 215842 233940 215852
rect 232540 212482 232596 212492
rect 211708 210802 211764 210812
rect 238588 209972 238644 240072
rect 239260 225092 239316 240072
rect 239260 225026 239316 225036
rect 239932 224196 239988 240072
rect 240604 232708 240660 240072
rect 240604 232642 240660 232652
rect 241276 224308 241332 240072
rect 241948 238532 242004 240072
rect 241948 238466 242004 238476
rect 242620 238532 242676 240072
rect 242620 238466 242676 238476
rect 243292 238420 243348 240072
rect 243292 238354 243348 238364
rect 243964 237860 244020 240072
rect 244636 238308 244692 240072
rect 244636 238242 244692 238252
rect 243964 237794 244020 237804
rect 245308 237748 245364 240072
rect 245980 237972 246036 240072
rect 245980 237906 246036 237916
rect 245308 237682 245364 237692
rect 241276 224242 241332 224252
rect 239932 224130 239988 224140
rect 246652 213332 246708 240072
rect 247324 238532 247380 240072
rect 247324 238466 247380 238476
rect 247996 237524 248052 240072
rect 248668 238084 248724 240072
rect 249340 238196 249396 240072
rect 249340 238130 249396 238140
rect 248668 238018 248724 238028
rect 247996 237458 248052 237468
rect 246652 213266 246708 213276
rect 250012 210756 250068 240072
rect 250684 236180 250740 240072
rect 251356 236404 251412 240072
rect 251356 236338 251412 236348
rect 250684 236114 250740 236124
rect 252028 214228 252084 240072
rect 252700 216020 252756 240072
rect 253372 223300 253428 240072
rect 253372 223234 253428 223244
rect 252700 215954 252756 215964
rect 252028 214162 252084 214172
rect 254044 211652 254100 240072
rect 254716 215012 254772 240072
rect 255388 221284 255444 240072
rect 256060 221396 256116 240072
rect 256060 221330 256116 221340
rect 255388 221218 255444 221228
rect 254716 214946 254772 214956
rect 256732 212548 256788 240072
rect 257404 224532 257460 240072
rect 258076 229460 258132 240072
rect 258076 229394 258132 229404
rect 257404 224466 257460 224476
rect 256732 212482 256788 212492
rect 254044 211586 254100 211596
rect 258748 211428 258804 240072
rect 259420 226548 259476 240072
rect 260092 236628 260148 240072
rect 260092 236562 260148 236572
rect 259420 226482 259476 226492
rect 260764 211540 260820 240072
rect 261436 214116 261492 240072
rect 262108 214340 262164 240072
rect 262780 214452 262836 240072
rect 263452 214900 263508 240072
rect 264124 217588 264180 240072
rect 264796 218260 264852 240072
rect 264796 218194 264852 218204
rect 264124 217522 264180 217532
rect 263452 214834 263508 214844
rect 262780 214386 262836 214396
rect 262108 214274 262164 214284
rect 261436 214050 261492 214060
rect 265468 213108 265524 240072
rect 266140 218372 266196 240072
rect 266140 218306 266196 218316
rect 266812 217476 266868 240072
rect 267484 237076 267540 240072
rect 268184 240044 268660 240100
rect 268856 240044 269332 240100
rect 267484 237010 267540 237020
rect 268604 236964 268660 240044
rect 268604 236898 268660 236908
rect 266812 217410 266868 217420
rect 265468 213042 265524 213052
rect 260764 211474 260820 211484
rect 258748 211362 258804 211372
rect 250012 210690 250068 210700
rect 238588 209906 238644 209916
rect 184604 209458 184660 209468
rect 269276 143668 269332 240044
rect 269500 237076 269556 240072
rect 270200 240044 270452 240100
rect 269500 237010 269556 237020
rect 269724 238308 269780 238318
rect 269276 143602 269332 143612
rect 269388 236516 269444 236526
rect 53228 49588 53284 49598
rect 41132 4498 41188 4508
rect 41804 42868 41860 42878
rect 41804 480 41860 42812
rect 45612 5012 45668 5022
rect 45612 480 45668 4956
rect 49420 4340 49476 4350
rect 47516 4228 47572 4238
rect 47516 480 47572 4172
rect 49420 480 49476 4284
rect 53228 480 53284 49532
rect 95116 49588 95172 49598
rect 87500 48244 87556 48254
rect 85708 37940 85764 37950
rect 57148 37828 57204 37838
rect 55132 3444 55188 3454
rect 55132 480 55188 3388
rect 57148 480 57204 37772
rect 62748 27748 62804 27758
rect 58940 4116 58996 4126
rect 58940 480 58996 4060
rect 60844 3444 60900 3454
rect 60844 480 60900 3388
rect 62748 480 62804 27692
rect 79884 24612 79940 24622
rect 68460 24500 68516 24510
rect 66556 4900 66612 4910
rect 64652 4452 64708 4462
rect 64652 480 64708 4396
rect 66556 480 66612 4844
rect 68460 480 68516 24444
rect 74172 24388 74228 24398
rect 70364 4676 70420 4686
rect 70364 480 70420 4620
rect 72268 4564 72324 4574
rect 72268 480 72324 4508
rect 74172 480 74228 24332
rect 76076 5012 76132 5022
rect 76076 480 76132 4956
rect 77980 4788 78036 4798
rect 77980 480 78036 4732
rect 79884 480 79940 24556
rect 83692 4340 83748 4350
rect 81788 4228 81844 4238
rect 81788 480 81844 4172
rect 83692 480 83748 4284
rect 85708 480 85764 37884
rect 87500 480 87556 48188
rect 93212 48132 93268 48142
rect 89404 41188 89460 41198
rect 89404 480 89460 41132
rect 91532 3444 91588 3454
rect 91532 480 91588 3388
rect 26572 392 26824 480
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 480
rect 30380 392 30632 480
rect 32284 392 32536 480
rect 30408 -960 30632 392
rect 32312 -960 32536 392
rect 34216 392 34468 480
rect 34216 -960 34440 392
rect 36120 -960 36344 480
rect 37996 392 38248 480
rect 39900 392 40152 480
rect 41804 392 42056 480
rect 38024 -960 38248 392
rect 39928 -960 40152 392
rect 41832 -960 42056 392
rect 43736 -960 43960 480
rect 45612 392 45864 480
rect 47516 392 47768 480
rect 49420 392 49672 480
rect 45640 -960 45864 392
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 -960 51576 480
rect 53228 392 53480 480
rect 55132 392 55384 480
rect 53256 -960 53480 392
rect 55160 -960 55384 392
rect 57064 -960 57288 480
rect 58940 392 59192 480
rect 60844 392 61096 480
rect 62748 392 63000 480
rect 64652 392 64904 480
rect 66556 392 66808 480
rect 68460 392 68712 480
rect 70364 392 70616 480
rect 72268 392 72520 480
rect 74172 392 74424 480
rect 76076 392 76328 480
rect 77980 392 78232 480
rect 79884 392 80136 480
rect 81788 392 82040 480
rect 83692 392 83944 480
rect 58968 -960 59192 392
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 64680 -960 64904 392
rect 66584 -960 66808 392
rect 68488 -960 68712 392
rect 70392 -960 70616 392
rect 72296 -960 72520 392
rect 74200 -960 74424 392
rect 76104 -960 76328 392
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 83720 -960 83944 392
rect 85624 -960 85848 480
rect 87500 392 87752 480
rect 89404 392 89656 480
rect 87528 -960 87752 392
rect 89432 -960 89656 392
rect 91336 392 91588 480
rect 93212 480 93268 48076
rect 95116 480 95172 49532
rect 97356 48692 97412 50120
rect 197932 49812 197988 49822
rect 97356 47908 97412 48636
rect 123676 49700 123732 49710
rect 116060 48132 116116 48142
rect 97356 47842 97412 47852
rect 98924 48020 98980 48030
rect 97020 34468 97076 34478
rect 97020 480 97076 34412
rect 98924 480 98980 47964
rect 110348 48020 110404 48030
rect 104636 47908 104692 47918
rect 100828 41300 100884 41310
rect 100828 480 100884 41244
rect 102732 34580 102788 34590
rect 102732 480 102788 34524
rect 104636 480 104692 47852
rect 106540 38052 106596 38062
rect 106540 480 106596 37996
rect 108444 34692 108500 34702
rect 108444 480 108500 34636
rect 110348 480 110404 47964
rect 114380 4676 114436 4686
rect 112476 4228 112532 4238
rect 112476 480 112532 4172
rect 114380 480 114436 4620
rect 93212 392 93464 480
rect 95116 392 95368 480
rect 97020 392 97272 480
rect 98924 392 99176 480
rect 100828 392 101080 480
rect 102732 392 102984 480
rect 104636 392 104888 480
rect 106540 392 106792 480
rect 108444 392 108696 480
rect 110348 392 110600 480
rect 91336 -960 91560 392
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 98952 -960 99176 392
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 -960 106792 392
rect 108472 -960 108696 392
rect 110376 -960 110600 392
rect 112280 392 112532 480
rect 114184 392 114436 480
rect 116060 480 116116 48076
rect 121772 44548 121828 44558
rect 117964 38164 118020 38174
rect 117964 480 118020 38108
rect 119868 31108 119924 31118
rect 119868 480 119924 31052
rect 121772 480 121828 44492
rect 123676 480 123732 49644
rect 190316 48468 190372 48478
rect 186508 48356 186564 48366
rect 138908 48244 138964 48254
rect 133196 44772 133252 44782
rect 127484 44660 127540 44670
rect 125580 34804 125636 34814
rect 125580 480 125636 34748
rect 127484 480 127540 44604
rect 129388 41412 129444 41422
rect 129388 480 129444 41356
rect 131292 31220 131348 31230
rect 131292 480 131348 31164
rect 133196 480 133252 44716
rect 135100 38388 135156 38398
rect 135100 480 135156 38332
rect 137004 38276 137060 38286
rect 137004 480 137060 38220
rect 138908 480 138964 48188
rect 184604 45332 184660 45342
rect 178892 45220 178948 45230
rect 167468 45108 167524 45118
rect 144620 44996 144676 45006
rect 140812 26068 140868 26078
rect 140812 480 140868 26012
rect 142940 3444 142996 3454
rect 142940 480 142996 3388
rect 116060 392 116312 480
rect 117964 392 118216 480
rect 119868 392 120120 480
rect 121772 392 122024 480
rect 123676 392 123928 480
rect 125580 392 125832 480
rect 127484 392 127736 480
rect 129388 392 129640 480
rect 131292 392 131544 480
rect 133196 392 133448 480
rect 135100 392 135352 480
rect 137004 392 137256 480
rect 138908 392 139160 480
rect 140812 392 141064 480
rect 112280 -960 112504 392
rect 114184 -960 114408 392
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 -960 120120 392
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 392
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 392 142996 480
rect 144620 480 144676 44940
rect 148428 44884 148484 44894
rect 146748 7588 146804 7598
rect 146748 480 146804 7532
rect 144620 392 144872 480
rect 142744 -960 142968 392
rect 144648 -960 144872 392
rect 146552 392 146804 480
rect 148428 480 148484 44828
rect 161756 41748 161812 41758
rect 156044 41636 156100 41646
rect 150332 41524 150388 41534
rect 150332 480 150388 41468
rect 152236 17668 152292 17678
rect 152236 480 152292 17612
rect 154364 4340 154420 4350
rect 154364 480 154420 4284
rect 148428 392 148680 480
rect 150332 392 150584 480
rect 152236 392 152488 480
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 392 154420 480
rect 156044 480 156100 41580
rect 159852 31332 159908 31342
rect 158172 5908 158228 5918
rect 158172 480 158228 5852
rect 156044 392 156296 480
rect 154168 -960 154392 392
rect 156072 -960 156296 392
rect 157976 392 158228 480
rect 159852 480 159908 31276
rect 161756 480 161812 41692
rect 163660 12628 163716 12638
rect 163660 480 163716 12572
rect 165788 4452 165844 4462
rect 165788 480 165844 4396
rect 159852 392 160104 480
rect 161756 392 162008 480
rect 163660 392 163912 480
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 -960 162008 392
rect 163688 -960 163912 392
rect 165592 392 165844 480
rect 167468 480 167524 45052
rect 175084 42980 175140 42990
rect 173180 41860 173236 41870
rect 169372 29428 169428 29438
rect 169372 480 169428 29372
rect 171500 4116 171556 4126
rect 171500 480 171556 4060
rect 167468 392 167720 480
rect 169372 392 169624 480
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 392 171556 480
rect 173180 480 173236 41804
rect 175084 480 175140 42924
rect 176988 38500 177044 38510
rect 176988 480 177044 38444
rect 178892 480 178948 45164
rect 181020 4900 181076 4910
rect 181020 480 181076 4844
rect 182924 4564 182980 4574
rect 182924 480 182980 4508
rect 173180 392 173432 480
rect 175084 392 175336 480
rect 176988 392 177240 480
rect 178892 392 179144 480
rect 171304 -960 171528 392
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 392 181076 480
rect 182728 392 182980 480
rect 184604 480 184660 45276
rect 186508 480 186564 48300
rect 188412 31444 188468 31454
rect 188412 480 188468 31388
rect 190316 480 190372 48412
rect 196028 41076 196084 41086
rect 192220 24724 192276 24734
rect 192220 480 192276 24668
rect 194348 4788 194404 4798
rect 194348 480 194404 4732
rect 184604 392 184856 480
rect 186508 392 186760 480
rect 188412 392 188664 480
rect 190316 392 190568 480
rect 192220 392 192472 480
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 392
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 392 194404 480
rect 196028 480 196084 41020
rect 197932 480 197988 49756
rect 201740 48580 201796 48590
rect 199948 41972 200004 41982
rect 199948 480 200004 41916
rect 201740 480 201796 48524
rect 207452 47796 207508 47806
rect 203644 44436 203700 44446
rect 203644 480 203700 44380
rect 205772 5012 205828 5022
rect 205772 480 205828 4956
rect 196028 392 196280 480
rect 197932 392 198184 480
rect 194152 -960 194376 392
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 -960 200088 480
rect 201740 392 201992 480
rect 203644 392 203896 480
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 392 205828 480
rect 207452 480 207508 47740
rect 212268 47684 212324 50120
rect 269388 48580 269444 236460
rect 269612 231812 269668 231822
rect 269388 48514 269444 48524
rect 269500 211316 269556 211326
rect 212268 47618 212324 47628
rect 269500 47684 269556 211260
rect 269500 47618 269556 47628
rect 269612 41076 269668 231756
rect 269612 41010 269668 41020
rect 269724 12628 269780 238252
rect 269836 237524 269892 237534
rect 269836 24724 269892 237468
rect 270396 236964 270452 240044
rect 270396 236898 270452 236908
rect 270732 238532 270788 238542
rect 270620 232708 270676 232718
rect 269836 24658 269892 24668
rect 270508 213332 270564 213342
rect 269724 12562 269780 12572
rect 270508 4900 270564 213276
rect 270620 41412 270676 232652
rect 270732 48356 270788 238476
rect 270844 159348 270900 240072
rect 271068 234500 271124 234510
rect 270844 159282 270900 159292
rect 270956 225092 271012 225102
rect 270732 48290 270788 48300
rect 270620 41346 270676 41356
rect 270956 38164 271012 225036
rect 271068 47908 271124 234444
rect 271068 47842 271124 47852
rect 271180 231476 271236 231486
rect 271180 44660 271236 231420
rect 271292 228340 271348 228350
rect 271292 47796 271348 228284
rect 271516 152292 271572 240072
rect 272188 210868 272244 240072
rect 272412 211316 272468 211326
rect 272188 210802 272244 210812
rect 272300 210980 272356 210990
rect 271516 152226 271572 152236
rect 272188 209972 272244 209982
rect 271292 47730 271348 47740
rect 271180 44594 271236 44604
rect 270956 38098 271012 38108
rect 270508 4834 270564 4844
rect 211484 4676 211540 4686
rect 209580 4116 209636 4126
rect 209580 480 209636 4060
rect 211484 480 211540 4620
rect 272188 4228 272244 209916
rect 272300 160468 272356 210924
rect 272412 172116 272468 211260
rect 272860 210980 272916 240072
rect 272860 210914 272916 210924
rect 272972 231476 273028 231486
rect 272636 209972 272692 209982
rect 272524 209188 272580 209198
rect 272524 175028 272580 209132
rect 272636 177940 272692 209916
rect 272748 209860 272804 209870
rect 272748 180852 272804 209804
rect 272748 180786 272804 180796
rect 272636 177874 272692 177884
rect 272524 174962 272580 174972
rect 272412 172050 272468 172060
rect 272300 160402 272356 160412
rect 272524 153636 272580 153646
rect 272300 145348 272356 145358
rect 272300 36820 272356 145292
rect 272412 142996 272468 143006
rect 272412 50372 272468 142940
rect 272524 131348 272580 153580
rect 272524 131282 272580 131292
rect 272972 99316 273028 231420
rect 273532 211092 273588 240072
rect 273868 238196 273924 238206
rect 273532 211026 273588 211036
rect 273756 236068 273812 236078
rect 273756 235172 273812 236012
rect 273084 205940 273140 205950
rect 273084 102228 273140 205884
rect 273420 154532 273476 154542
rect 273196 154308 273252 154318
rect 273196 134260 273252 154252
rect 273196 134194 273252 134204
rect 273308 145460 273364 145470
rect 273308 128436 273364 145404
rect 273420 137172 273476 154476
rect 273756 153636 273812 235116
rect 273756 153570 273812 153580
rect 273532 143780 273588 143790
rect 273532 142996 273588 143724
rect 273532 142930 273588 142940
rect 273420 137106 273476 137116
rect 273308 128370 273364 128380
rect 273756 126868 273812 126878
rect 273756 125524 273812 126812
rect 273756 125458 273812 125468
rect 273084 102162 273140 102172
rect 272972 99250 273028 99260
rect 273308 101668 273364 101678
rect 273308 73108 273364 101612
rect 273308 73042 273364 73052
rect 273084 70196 273140 70206
rect 272972 67284 273028 67294
rect 272972 50596 273028 67228
rect 273084 52836 273140 70140
rect 273084 52770 273140 52780
rect 273196 61460 273252 61470
rect 272972 50530 273028 50540
rect 272412 50306 272468 50316
rect 273196 49700 273252 61404
rect 273196 49634 273252 49644
rect 273868 44436 273924 238140
rect 273980 238084 274036 238094
rect 273980 49812 274036 238028
rect 273980 49746 274036 49756
rect 274092 228228 274148 228238
rect 273868 44370 273924 44380
rect 274092 41636 274148 228172
rect 274204 160356 274260 240072
rect 274428 231588 274484 231598
rect 274204 160290 274260 160300
rect 274316 224980 274372 224990
rect 274316 41860 274372 224924
rect 274428 48244 274484 231532
rect 274428 48178 274484 48188
rect 274540 228116 274596 228126
rect 274540 44996 274596 228060
rect 274652 210084 274708 210094
rect 274652 154420 274708 210028
rect 274876 160692 274932 240072
rect 274876 160626 274932 160636
rect 275548 160580 275604 240072
rect 275772 227668 275828 227678
rect 275548 160514 275604 160524
rect 275660 224308 275716 224318
rect 274652 154354 274708 154364
rect 274652 141988 274708 141998
rect 274652 81844 274708 141932
rect 274652 81778 274708 81788
rect 275436 58548 275492 58558
rect 275436 49812 275492 58492
rect 275548 52724 275604 52734
rect 275548 50708 275604 52668
rect 275548 50642 275604 50652
rect 275436 49746 275492 49756
rect 274540 44930 274596 44940
rect 274316 41794 274372 41804
rect 274092 41570 274148 41580
rect 275660 38388 275716 224252
rect 275772 41524 275828 227612
rect 275884 224420 275940 224430
rect 275884 41748 275940 224364
rect 276220 197204 276276 240072
rect 276220 197138 276276 197148
rect 276332 224420 276388 224430
rect 275884 41682 275940 41692
rect 275772 41458 275828 41468
rect 275660 38322 275716 38332
rect 272300 36754 272356 36764
rect 276332 24500 276388 224364
rect 276444 219268 276500 219278
rect 276444 38500 276500 219212
rect 276892 150948 276948 240072
rect 276892 150882 276948 150892
rect 277228 237860 277284 237870
rect 276556 138628 276612 138638
rect 276556 76020 276612 138572
rect 276556 75954 276612 75964
rect 276556 64372 276612 64382
rect 276556 49588 276612 64316
rect 276556 49522 276612 49532
rect 276444 38434 276500 38444
rect 276332 24434 276388 24444
rect 277228 5908 277284 237804
rect 277564 237860 277620 240072
rect 278236 238084 278292 240072
rect 278908 238196 278964 240072
rect 278908 238130 278964 238140
rect 278236 238018 278292 238028
rect 277564 237794 277620 237804
rect 279020 237972 279076 237982
rect 278908 237748 278964 237758
rect 278124 224308 278180 224318
rect 278012 219716 278068 219726
rect 277228 5842 277284 5852
rect 277340 210756 277396 210766
rect 272188 4162 272244 4172
rect 277340 4116 277396 210700
rect 278012 31444 278068 219660
rect 278124 41972 278180 224252
rect 278236 132020 278292 132030
rect 278236 78932 278292 131964
rect 278236 78866 278292 78876
rect 278124 41906 278180 41916
rect 278012 31378 278068 31388
rect 278908 29428 278964 237692
rect 279020 42980 279076 237916
rect 279580 237748 279636 240072
rect 279580 237682 279636 237692
rect 279020 42914 279076 42924
rect 279692 236292 279748 236302
rect 279692 33684 279748 236236
rect 279692 33618 279748 33628
rect 279804 227668 279860 227678
rect 279804 31332 279860 227612
rect 279916 222852 279972 222862
rect 279916 38276 279972 222796
rect 280028 219828 280084 219838
rect 280028 42868 280084 219772
rect 280252 155988 280308 240072
rect 280924 238308 280980 240072
rect 280924 238242 280980 238252
rect 280252 155922 280308 155932
rect 280364 219940 280420 219950
rect 280364 44884 280420 219884
rect 281596 152852 281652 240072
rect 282268 237972 282324 240072
rect 282268 237906 282324 237916
rect 282940 155540 282996 240072
rect 283164 226212 283220 226222
rect 282940 155474 282996 155484
rect 283052 222740 283108 222750
rect 281596 152786 281652 152796
rect 280364 44818 280420 44828
rect 280028 42802 280084 42812
rect 279916 38210 279972 38220
rect 279804 31266 279860 31276
rect 283052 31220 283108 222684
rect 283164 34804 283220 226156
rect 283612 152180 283668 240072
rect 283612 152114 283668 152124
rect 284284 150836 284340 240072
rect 284956 151060 285012 240072
rect 284956 150994 285012 151004
rect 284284 150770 284340 150780
rect 285628 149156 285684 240072
rect 286300 238532 286356 240072
rect 286300 238466 286356 238476
rect 286636 226324 286692 226334
rect 285628 149090 285684 149100
rect 286412 226100 286468 226110
rect 283164 34738 283220 34748
rect 286412 34692 286468 226044
rect 286412 34626 286468 34636
rect 286636 34468 286692 226268
rect 286860 225988 286916 225998
rect 286860 34580 286916 225932
rect 286972 159460 287028 240072
rect 286972 159394 287028 159404
rect 287644 159124 287700 240072
rect 287644 159058 287700 159068
rect 288204 239316 288260 239326
rect 286860 34514 286916 34524
rect 286636 34402 286692 34412
rect 283052 31154 283108 31164
rect 278908 29362 278964 29372
rect 288204 5012 288260 239260
rect 288316 158900 288372 240072
rect 288988 238420 289044 240072
rect 288988 238354 289044 238364
rect 289660 159012 289716 240072
rect 289660 158946 289716 158956
rect 289772 234388 289828 234398
rect 288316 158834 288372 158844
rect 288988 55636 289044 55646
rect 288988 50484 289044 55580
rect 288988 50418 289044 50428
rect 288204 4946 288260 4956
rect 289772 4676 289828 234332
rect 289884 226436 289940 226446
rect 289884 31108 289940 226380
rect 289884 31042 289940 31052
rect 289996 216468 290052 216478
rect 289996 24388 290052 216412
rect 290220 216356 290276 216366
rect 290220 48580 290276 216300
rect 290332 161924 290388 240072
rect 290332 161858 290388 161868
rect 291004 150724 291060 240072
rect 291004 150658 291060 150668
rect 291676 150388 291732 240072
rect 292348 237076 292404 240072
rect 292348 237010 292404 237020
rect 293020 162148 293076 240072
rect 293720 240044 293860 240100
rect 293244 238308 293300 238318
rect 293020 162082 293076 162092
rect 293132 211652 293188 211662
rect 291676 150322 291732 150332
rect 293132 123620 293188 211596
rect 293244 152404 293300 238252
rect 293804 236964 293860 240044
rect 293804 236898 293860 236908
rect 293244 152338 293300 152348
rect 294364 152068 294420 240072
rect 295064 240044 295652 240100
rect 294812 238532 294868 238542
rect 294812 155652 294868 238476
rect 295596 236964 295652 240044
rect 295596 236898 295652 236908
rect 294812 155586 294868 155596
rect 294364 152002 294420 152012
rect 295708 149492 295764 240072
rect 295708 149426 295764 149436
rect 296380 149268 296436 240072
rect 296380 149202 296436 149212
rect 296492 215012 296548 215022
rect 296492 123732 296548 214956
rect 297052 155428 297108 240072
rect 297724 236964 297780 240072
rect 297724 236898 297780 236908
rect 297052 155362 297108 155372
rect 298172 236404 298228 236414
rect 298172 123956 298228 236348
rect 298396 162036 298452 240072
rect 298396 161970 298452 161980
rect 299068 148708 299124 240072
rect 299740 236964 299796 240072
rect 299740 236898 299796 236908
rect 299964 238420 300020 238430
rect 299068 148642 299124 148652
rect 299852 212548 299908 212558
rect 298172 123890 298228 123900
rect 296492 123666 296548 123676
rect 293132 123554 293188 123564
rect 299852 123508 299908 212492
rect 299964 159236 300020 238364
rect 299964 159170 300020 159180
rect 300412 158788 300468 240072
rect 301084 160468 301140 240072
rect 301644 238196 301700 238206
rect 301084 160402 301140 160412
rect 301532 236180 301588 236190
rect 300412 158722 300468 158732
rect 301532 124292 301588 236124
rect 301644 155764 301700 238140
rect 301756 233492 301812 240072
rect 301756 233426 301812 233436
rect 302428 228452 302484 240072
rect 319900 240100 319956 240110
rect 303100 240034 303156 240044
rect 302428 228386 302484 228396
rect 303548 237972 303604 237982
rect 303436 221396 303492 221406
rect 303212 221284 303268 221294
rect 301644 155698 301700 155708
rect 303100 213108 303156 213118
rect 303100 133812 303156 213052
rect 303100 133746 303156 133756
rect 303212 127428 303268 221228
rect 303212 127362 303268 127372
rect 303324 216020 303380 216030
rect 301532 124226 301588 124236
rect 303324 124068 303380 215964
rect 303436 130452 303492 221340
rect 303548 149604 303604 237916
rect 303772 236292 303828 240072
rect 303772 236226 303828 236236
rect 303996 238084 304052 238094
rect 303548 149538 303604 149548
rect 303660 218372 303716 218382
rect 303660 133700 303716 218316
rect 303660 133634 303716 133644
rect 303884 217476 303940 217486
rect 303884 133588 303940 217420
rect 303996 155876 304052 238028
rect 304444 236516 304500 240072
rect 304444 236450 304500 236460
rect 304892 239428 304948 239438
rect 303996 155810 304052 155820
rect 304892 152516 304948 239372
rect 305004 237860 305060 237870
rect 305004 156212 305060 237804
rect 305116 236740 305172 240072
rect 305116 236674 305172 236684
rect 305788 236404 305844 240072
rect 306460 237636 306516 240072
rect 306460 237570 306516 237580
rect 305788 236338 305844 236348
rect 307132 236180 307188 240072
rect 307132 236114 307188 236124
rect 307356 239316 307412 239326
rect 307356 236628 307412 239260
rect 307356 236068 307412 236572
rect 307356 236002 307412 236012
rect 307804 236068 307860 240072
rect 308476 237524 308532 240072
rect 308476 237458 308532 237468
rect 308700 237748 308756 237758
rect 307804 236002 307860 236012
rect 305116 231364 305172 231374
rect 305116 204148 305172 231308
rect 305116 204082 305172 204092
rect 306572 223300 306628 223310
rect 305004 156146 305060 156156
rect 304892 152450 304948 152460
rect 303884 133522 303940 133532
rect 303436 130386 303492 130396
rect 306572 124180 306628 223244
rect 307020 218260 307076 218270
rect 306796 217588 306852 217598
rect 306684 214452 306740 214462
rect 306684 127092 306740 214396
rect 306796 130228 306852 217532
rect 306796 130162 306852 130172
rect 306908 214340 306964 214350
rect 306908 127204 306964 214284
rect 307020 133924 307076 218204
rect 307020 133858 307076 133868
rect 307132 214900 307188 214910
rect 307132 130340 307188 214844
rect 308252 214228 308308 214238
rect 307132 130274 307188 130284
rect 307244 211540 307300 211550
rect 307244 127316 307300 211484
rect 307244 127250 307300 127260
rect 306908 127138 306964 127148
rect 306684 127026 306740 127036
rect 306572 124114 306628 124124
rect 303324 124002 303380 124012
rect 299852 123442 299908 123452
rect 308252 123396 308308 214172
rect 308700 156100 308756 237692
rect 309148 230132 309204 240072
rect 309820 230916 309876 240072
rect 310492 237748 310548 240072
rect 311164 238196 311220 240072
rect 311164 238130 311220 238140
rect 311836 237860 311892 240072
rect 312508 238308 312564 240072
rect 313180 238420 313236 240072
rect 313180 238354 313236 238364
rect 312508 238242 312564 238252
rect 311836 237794 311892 237804
rect 310492 237682 310548 237692
rect 312508 237524 312564 237534
rect 312508 235060 312564 237468
rect 313852 237524 313908 240072
rect 314524 237972 314580 240072
rect 314524 237906 314580 237916
rect 313852 237458 313908 237468
rect 312508 234994 312564 235004
rect 315196 234948 315252 240072
rect 315868 238084 315924 240072
rect 315868 238018 315924 238028
rect 316540 236852 316596 240072
rect 316540 236786 316596 236796
rect 318332 239540 318388 239550
rect 315196 234882 315252 234892
rect 311164 234612 311220 234622
rect 309820 230850 309876 230860
rect 309932 232708 309988 232718
rect 309148 230066 309204 230076
rect 308700 156034 308756 156044
rect 308252 123330 308308 123340
rect 309932 116788 309988 232652
rect 311052 230244 311108 230254
rect 310156 229460 310212 229470
rect 310044 224532 310100 224542
rect 310044 123844 310100 224476
rect 310044 123778 310100 123788
rect 310156 119700 310212 229404
rect 310268 219604 310324 219614
rect 310268 157668 310324 219548
rect 310940 214676 310996 214686
rect 310380 211092 310436 211102
rect 310380 160244 310436 211036
rect 310380 160178 310436 160188
rect 310604 210980 310660 210990
rect 310604 159908 310660 210924
rect 310940 160690 310996 214620
rect 310940 160638 310942 160690
rect 310994 160638 310996 160690
rect 310940 160626 310996 160638
rect 310604 159842 310660 159852
rect 310268 157602 310324 157612
rect 310156 119634 310212 119644
rect 309932 116722 309988 116732
rect 311052 105140 311108 230188
rect 311052 105074 311108 105084
rect 311164 96404 311220 234556
rect 311612 233156 311668 233166
rect 311612 196952 311668 233100
rect 314972 229908 315028 229918
rect 312732 217924 312788 217934
rect 312732 196952 312788 217868
rect 313852 217812 313908 217822
rect 313852 196952 313908 217756
rect 314972 196952 315028 229852
rect 317212 221060 317268 221070
rect 316092 219492 316148 219502
rect 316092 196952 316148 219436
rect 317212 196952 317268 221004
rect 318332 196952 318388 239484
rect 319228 239540 319284 240072
rect 325836 240100 325892 240110
rect 319900 240034 319956 240044
rect 319228 239474 319284 239484
rect 321244 238532 321300 240072
rect 321244 238466 321300 238476
rect 321916 238532 321972 240072
rect 325836 239428 325892 240044
rect 325836 239362 325892 239372
rect 321916 238466 321972 238476
rect 330652 234836 330708 234846
rect 321692 234164 321748 234174
rect 320572 233044 320628 233054
rect 319452 231252 319508 231262
rect 319452 196952 319508 231196
rect 320572 196952 320628 232988
rect 321692 196952 321748 234108
rect 326172 232932 326228 232942
rect 325052 229796 325108 229806
rect 322812 228004 322868 228014
rect 321804 224756 321860 224766
rect 321804 214228 321860 224700
rect 321804 214162 321860 214172
rect 322812 196952 322868 227948
rect 323932 217700 323988 217710
rect 323932 196952 323988 217644
rect 325052 196952 325108 229740
rect 326172 196952 326228 232876
rect 328412 231140 328468 231150
rect 327292 224868 327348 224878
rect 327292 196952 327348 224812
rect 328412 196952 328468 231084
rect 329532 227892 329588 227902
rect 329532 196952 329588 227836
rect 330652 196952 330708 234780
rect 336028 231140 336084 240268
rect 336028 231074 336084 231084
rect 336252 232820 336308 232830
rect 335132 231028 335188 231038
rect 332892 229684 332948 229694
rect 331772 223076 331828 223086
rect 331772 196952 331828 223020
rect 331996 222964 332052 222974
rect 331996 209188 332052 222908
rect 331996 209122 332052 209132
rect 332892 196952 332948 229628
rect 334012 219380 334068 219390
rect 334012 196952 334068 219324
rect 335132 196952 335188 230972
rect 336252 196952 336308 232764
rect 337148 219940 337204 240604
rect 337148 219874 337204 219884
rect 337372 224644 337428 224654
rect 337372 196952 337428 224588
rect 338492 223188 338548 223198
rect 338492 196952 338548 223132
rect 339276 216468 339332 243516
rect 339276 216402 339332 216412
rect 339388 198212 339444 354508
rect 339388 198146 339444 198156
rect 339500 197876 339556 383628
rect 339612 381444 339668 381454
rect 339612 239428 339668 381388
rect 339948 281204 340004 281214
rect 339948 280644 340004 281148
rect 339948 280578 340004 280588
rect 339612 239362 339668 239372
rect 340060 236852 340116 388780
rect 340172 237524 340228 408268
rect 340284 360500 340340 410088
rect 341292 409668 341348 409678
rect 340284 359604 340340 360444
rect 340284 359538 340340 359548
rect 340396 396788 340452 396798
rect 340172 237458 340228 237468
rect 340060 236786 340116 236796
rect 340396 236068 340452 396732
rect 340732 389396 340788 389406
rect 340396 236002 340452 236012
rect 340508 389172 340564 389182
rect 340508 230132 340564 389116
rect 340732 234948 340788 389340
rect 340956 389284 341012 389294
rect 340956 235060 341012 389228
rect 341180 381892 341236 381902
rect 341068 252196 341124 252206
rect 341068 243572 341124 252140
rect 341068 243506 341124 243516
rect 341180 239092 341236 381836
rect 341292 291620 341348 409612
rect 341404 294868 341460 410396
rect 429660 410116 429716 410126
rect 345324 394884 345380 394894
rect 343756 393428 343812 393438
rect 343532 393316 343588 393326
rect 341852 392756 341908 392766
rect 341628 381556 341684 381566
rect 341404 294308 341460 294812
rect 341404 294242 341460 294252
rect 341516 380212 341572 380222
rect 341292 291554 341348 291564
rect 341292 282660 341348 282670
rect 341292 240660 341348 282604
rect 341292 240594 341348 240604
rect 341404 261156 341460 261166
rect 341180 239026 341236 239036
rect 340956 234994 341012 235004
rect 340732 234882 340788 234892
rect 340508 230066 340564 230076
rect 340732 227780 340788 227790
rect 339500 197810 339556 197820
rect 339612 220948 339668 220958
rect 339612 196952 339668 220892
rect 340732 196952 340788 227724
rect 341404 222740 341460 261100
rect 341404 222674 341460 222684
rect 341516 197764 341572 380156
rect 341516 197698 341572 197708
rect 341628 196532 341684 381500
rect 341740 234724 341796 234734
rect 341740 208348 341796 234668
rect 341852 233492 341908 392700
rect 342972 390628 343028 390638
rect 341852 233426 341908 233436
rect 341964 389508 342020 389518
rect 341964 230916 342020 389452
rect 342860 388948 342916 388958
rect 342076 385924 342132 385934
rect 342076 319844 342132 385868
rect 342076 319778 342132 319788
rect 342860 297388 342916 388892
rect 342748 297332 342916 297388
rect 342748 292516 342804 297332
rect 342972 295204 343028 390572
rect 342972 295138 343028 295148
rect 343084 387268 343140 387278
rect 343084 293188 343140 387212
rect 343532 371364 343588 393260
rect 343756 374052 343812 393372
rect 343756 373986 343812 373996
rect 345212 385364 345268 385374
rect 343532 371298 343588 371308
rect 344764 364196 344820 364206
rect 343532 345380 343588 345390
rect 343084 293122 343140 293132
rect 343196 340900 343252 340910
rect 342748 292450 342804 292460
rect 342076 290724 342132 290734
rect 342076 234612 342132 290668
rect 342860 273700 342916 273710
rect 342748 262948 342804 262958
rect 342748 241668 342804 262892
rect 342748 241602 342804 241612
rect 342076 234546 342132 234556
rect 342188 240772 342244 240782
rect 341964 230850 342020 230860
rect 342188 219268 342244 240716
rect 342860 234388 342916 273644
rect 342972 272804 343028 272814
rect 342972 241220 343028 272748
rect 342972 241154 343028 241164
rect 343084 266532 343140 266542
rect 343084 240996 343140 266476
rect 343084 240930 343140 240940
rect 342860 234322 342916 234332
rect 342188 219202 342244 219212
rect 341740 208292 341908 208348
rect 341852 196952 341908 208292
rect 342972 201572 343028 201582
rect 342972 196952 343028 201516
rect 341628 196466 341684 196476
rect 343196 196420 343252 340844
rect 343308 264740 343364 264750
rect 343308 241892 343364 264684
rect 343532 251188 343588 345324
rect 344092 339108 344148 339118
rect 343532 251122 343588 251132
rect 343644 338212 343700 338222
rect 343308 241826 343364 241836
rect 343420 249508 343476 249518
rect 343420 231252 343476 249452
rect 343420 231186 343476 231196
rect 343532 240436 343588 240446
rect 343532 215908 343588 240380
rect 343532 215842 343588 215852
rect 343644 208348 343700 338156
rect 343756 240884 343812 240894
rect 343756 224308 343812 240828
rect 343756 224242 343812 224252
rect 343980 209524 344036 209534
rect 343644 208292 343924 208348
rect 343868 196530 343924 208292
rect 343980 202468 344036 209468
rect 344092 208348 344148 339052
rect 344316 278852 344372 278862
rect 344316 264628 344372 278796
rect 344316 264562 344372 264572
rect 344092 208292 344372 208348
rect 343980 202412 344148 202468
rect 344092 196952 344148 202412
rect 343868 196478 343870 196530
rect 343922 196478 343924 196530
rect 343868 196466 343924 196478
rect 343196 196354 343252 196364
rect 344316 196420 344372 208292
rect 344316 196354 344372 196364
rect 344764 196420 344820 364140
rect 345100 252084 345156 252094
rect 345100 240324 345156 252028
rect 345100 240258 345156 240268
rect 345100 212660 345156 212670
rect 345100 197876 345156 212604
rect 345212 198100 345268 385308
rect 345324 237860 345380 394828
rect 345548 386148 345604 386158
rect 345324 237794 345380 237804
rect 345436 358820 345492 358830
rect 345436 208348 345492 358764
rect 345548 336084 345604 386092
rect 345660 367108 345716 410088
rect 350476 403396 350532 403406
rect 347228 396900 347284 396910
rect 345660 367042 345716 367052
rect 346444 379764 346500 379774
rect 345548 229460 345604 336028
rect 345548 229394 345604 229404
rect 345660 342692 345716 342702
rect 345436 208292 345604 208348
rect 345212 198034 345268 198044
rect 345100 197820 345268 197876
rect 345212 196952 345268 197820
rect 345548 196644 345604 208292
rect 345548 196578 345604 196588
rect 344988 196532 345044 196542
rect 344988 196438 345044 196476
rect 344764 196354 344820 196364
rect 345660 196420 345716 342636
rect 345996 272132 346052 272142
rect 345772 252532 345828 252542
rect 345772 208348 345828 252476
rect 345772 208292 345940 208348
rect 345660 196354 345716 196364
rect 345884 196420 345940 208292
rect 345996 198212 346052 272076
rect 346108 263844 346164 263854
rect 346108 240548 346164 263788
rect 346108 240482 346164 240492
rect 346220 253092 346276 253102
rect 346220 240436 346276 253036
rect 346220 240370 346276 240380
rect 345996 198146 346052 198156
rect 345884 196354 345940 196364
rect 311276 160692 311332 160702
rect 313404 160692 313460 160702
rect 311276 160690 311864 160692
rect 311276 160638 311278 160690
rect 311330 160638 311864 160690
rect 311276 160636 311864 160638
rect 311276 160626 311332 160636
rect 313404 160626 313460 160636
rect 314972 160132 315028 160142
rect 317436 160132 317492 160142
rect 316568 160076 317436 160132
rect 329084 160132 329140 160142
rect 314972 160066 315028 160076
rect 317436 160066 317492 160076
rect 318108 156996 318164 160104
rect 319676 157668 319732 160104
rect 319676 157602 319732 157612
rect 321244 157668 321300 160104
rect 321244 157602 321300 157612
rect 318108 156930 318164 156940
rect 322812 156884 322868 160104
rect 324380 157892 324436 160104
rect 324380 157826 324436 157836
rect 325948 157556 326004 160104
rect 327516 157780 327572 160104
rect 344764 160132 344820 160142
rect 329084 160066 329140 160076
rect 330652 157892 330708 160104
rect 330652 157826 330708 157836
rect 332220 157892 332276 160104
rect 332220 157826 332276 157836
rect 327516 157714 327572 157724
rect 325948 157490 326004 157500
rect 333788 157332 333844 160104
rect 335356 157892 335412 160104
rect 335356 157826 335412 157836
rect 336924 157556 336980 160104
rect 338492 158676 338548 160104
rect 340060 159572 340116 160104
rect 340060 159506 340116 159516
rect 338492 158610 338548 158620
rect 341628 157780 341684 160104
rect 343196 159796 343252 160104
rect 344764 160066 344820 160076
rect 343196 159730 343252 159740
rect 341628 157714 341684 157724
rect 346108 157892 346164 157902
rect 336924 157490 336980 157500
rect 346108 157444 346164 157836
rect 346444 157668 346500 379708
rect 346892 369572 346948 369582
rect 346556 196420 346612 196430
rect 346556 184828 346612 196364
rect 346556 184772 346836 184828
rect 346444 157602 346500 157612
rect 346108 157378 346164 157388
rect 346780 157444 346836 184772
rect 346892 167860 346948 369516
rect 347004 361508 347060 361518
rect 347004 171108 347060 361452
rect 347116 351652 347172 351662
rect 347116 172452 347172 351596
rect 347228 236180 347284 396844
rect 348572 370468 348628 370478
rect 347788 309540 347844 309550
rect 347676 296548 347732 296558
rect 347228 236114 347284 236124
rect 347564 284788 347620 284798
rect 347116 172386 347172 172396
rect 347004 171042 347060 171052
rect 347004 167860 347060 167870
rect 346892 167804 347004 167860
rect 347004 167794 347060 167804
rect 346780 157378 346836 157388
rect 333788 157266 333844 157276
rect 322812 156818 322868 156828
rect 345212 153860 345268 153870
rect 341852 147028 341908 147038
rect 341852 122612 341908 146972
rect 345212 126868 345268 153804
rect 345324 151844 345380 151854
rect 345324 140084 345380 151788
rect 345324 140018 345380 140028
rect 345212 126802 345268 126812
rect 341852 122546 341908 122556
rect 311164 96338 311220 96348
rect 307468 50372 307524 50382
rect 315308 50372 315364 50382
rect 307524 50316 307944 50372
rect 315112 50316 315308 50372
rect 307468 50306 307524 50316
rect 315308 50306 315364 50316
rect 293580 48692 293636 50120
rect 293580 48626 293636 48636
rect 290220 48514 290276 48524
rect 300748 48580 300804 50120
rect 300748 48514 300804 48524
rect 322252 48580 322308 50120
rect 322252 48514 322308 48524
rect 347564 48580 347620 284732
rect 347676 50372 347732 296492
rect 347788 238644 347844 309484
rect 347788 238578 347844 238588
rect 347900 198100 347956 198110
rect 347788 196532 347844 196542
rect 347788 157556 347844 196476
rect 347900 160020 347956 198044
rect 348572 171332 348628 370412
rect 350252 365092 350308 365102
rect 348572 171266 348628 171276
rect 348684 362404 348740 362414
rect 348684 169428 348740 362348
rect 348796 354340 348852 354350
rect 348796 172676 348852 354284
rect 348796 172610 348852 172620
rect 348908 352548 348964 352558
rect 348684 169362 348740 169372
rect 348908 168756 348964 352492
rect 349020 349860 349076 349870
rect 349020 174244 349076 349804
rect 349132 283892 349188 283902
rect 349132 242004 349188 283836
rect 349356 283780 349412 283790
rect 349132 241938 349188 241948
rect 349244 248612 349300 248622
rect 349020 174178 349076 174188
rect 348908 168690 348964 168700
rect 347900 159954 347956 159964
rect 347788 157490 347844 157500
rect 349244 150612 349300 248556
rect 349244 150546 349300 150556
rect 349356 148932 349412 283724
rect 349580 271908 349636 271918
rect 349468 257572 349524 257582
rect 349468 226100 349524 257516
rect 349580 240884 349636 271852
rect 349580 240818 349636 240828
rect 349468 226034 349524 226044
rect 349580 196308 349636 196318
rect 349580 160132 349636 196252
rect 350252 169540 350308 365036
rect 350364 356132 350420 356142
rect 350364 172788 350420 356076
rect 350476 237972 350532 403340
rect 350700 394100 350756 394110
rect 350476 237906 350532 237916
rect 350588 296548 350644 296558
rect 350364 172722 350420 172732
rect 350476 189812 350532 189822
rect 350252 169474 350308 169484
rect 349580 160066 349636 160076
rect 350476 153076 350532 189756
rect 350476 149548 350532 153020
rect 349356 148866 349412 148876
rect 350252 149492 350532 149548
rect 350588 162372 350644 296492
rect 350700 238196 350756 394044
rect 350924 392532 350980 392542
rect 350700 238130 350756 238140
rect 350812 305732 350868 305742
rect 350700 197428 350756 197438
rect 350700 164276 350756 197372
rect 350812 189812 350868 305676
rect 350924 237636 350980 392476
rect 351036 372260 351092 410088
rect 353612 408100 353668 408110
rect 351932 407876 351988 407886
rect 351932 385700 351988 407820
rect 352156 407764 352212 407774
rect 352156 397460 352212 407708
rect 352156 397394 352212 397404
rect 352268 401828 352324 401838
rect 351932 385634 351988 385644
rect 351036 372194 351092 372204
rect 351148 379876 351204 379886
rect 350924 237570 350980 237580
rect 351036 209972 351092 209982
rect 350812 189746 350868 189756
rect 350924 193284 350980 193294
rect 350700 164210 350756 164220
rect 350812 188132 350868 188142
rect 350812 186564 350868 188076
rect 350588 153524 350644 162316
rect 350700 160132 350756 160142
rect 350700 157220 350756 160076
rect 350700 157154 350756 157164
rect 350588 149548 350644 153468
rect 350588 149492 350756 149548
rect 350252 143780 350308 149492
rect 350700 145348 350756 149492
rect 350700 145282 350756 145292
rect 350252 143714 350308 143724
rect 350812 126028 350868 186508
rect 350252 125972 350868 126028
rect 350252 119364 350308 125972
rect 350252 101668 350308 119308
rect 350252 101602 350308 101612
rect 347676 50306 347732 50316
rect 347564 48514 347620 48524
rect 350924 48468 350980 193228
rect 351036 50260 351092 209916
rect 351148 156996 351204 379820
rect 351932 367780 351988 367790
rect 351260 313348 351316 313358
rect 351260 231364 351316 313292
rect 351372 268324 351428 268334
rect 351372 240772 351428 268268
rect 351372 240706 351428 240716
rect 351260 231298 351316 231308
rect 351820 236852 351876 236862
rect 351260 197316 351316 197326
rect 351260 184828 351316 197260
rect 351820 188132 351876 236796
rect 351820 188066 351876 188076
rect 351260 184772 351540 184828
rect 351484 157332 351540 184772
rect 351932 169652 351988 367724
rect 352044 359716 352100 359726
rect 352044 170996 352100 359660
rect 352156 348964 352212 348974
rect 352156 173684 352212 348908
rect 352268 238084 352324 401772
rect 352268 238018 352324 238028
rect 352380 397460 352436 397470
rect 352380 236292 352436 397404
rect 353612 385588 353668 408044
rect 355404 407316 355460 407326
rect 355180 407204 355236 407214
rect 353612 385522 353668 385532
rect 354172 405076 354228 405086
rect 352604 383124 352660 383134
rect 352380 236226 352436 236236
rect 352492 380660 352548 380670
rect 352492 331044 352548 380604
rect 352492 232708 352548 330988
rect 352604 305732 352660 383068
rect 352604 305666 352660 305676
rect 352828 379428 352884 379438
rect 352492 232642 352548 232652
rect 352156 173618 352212 173628
rect 352268 197204 352324 197214
rect 352044 170930 352100 170940
rect 351932 169586 351988 169596
rect 352268 164164 352324 197148
rect 352716 191716 352772 191726
rect 352268 164098 352324 164108
rect 352604 191604 352660 191614
rect 352492 159572 352548 159582
rect 352492 157668 352548 159516
rect 352492 157602 352548 157612
rect 351484 157266 351540 157276
rect 351148 156930 351204 156940
rect 352604 120260 352660 191548
rect 352604 120194 352660 120204
rect 351036 50194 351092 50204
rect 350924 48402 350980 48412
rect 352716 48356 352772 191660
rect 352828 156884 352884 379372
rect 353612 365988 353668 365998
rect 352828 156818 352884 156828
rect 352940 247828 352996 247838
rect 352940 151172 352996 247772
rect 353612 167636 353668 365932
rect 353724 357028 353780 357038
rect 353724 170884 353780 356972
rect 354060 346276 354116 346286
rect 353724 170818 353780 170828
rect 353836 294868 353892 294878
rect 353612 167570 353668 167580
rect 352940 151106 352996 151116
rect 353836 122052 353892 294812
rect 353836 121986 353892 121996
rect 353948 291508 354004 291518
rect 353948 120372 354004 291452
rect 354060 175252 354116 346220
rect 354172 238308 354228 405020
rect 355180 397348 355236 407148
rect 355180 397282 355236 397292
rect 355292 402612 355348 402622
rect 355292 382228 355348 402556
rect 355404 390740 355460 407260
rect 355404 390674 355460 390684
rect 355516 397012 355572 397022
rect 355292 382162 355348 382172
rect 355292 366884 355348 366894
rect 354172 238242 354228 238252
rect 354396 282212 354452 282222
rect 354060 175186 354116 175196
rect 354172 195972 354228 195982
rect 354172 174356 354228 195916
rect 354172 174290 354228 174300
rect 353948 120306 354004 120316
rect 352716 48290 352772 48300
rect 354396 48244 354452 282156
rect 354620 265636 354676 265646
rect 354620 227668 354676 265580
rect 354620 227602 354676 227612
rect 354508 195860 354564 195870
rect 354508 157780 354564 195804
rect 355292 167748 355348 366828
rect 355404 357924 355460 357934
rect 355404 172900 355460 357868
rect 355516 236404 355572 396956
rect 355740 389620 355796 389630
rect 355516 236338 355572 236348
rect 355628 348068 355684 348078
rect 355404 172834 355460 172844
rect 355516 210868 355572 210878
rect 355516 169092 355572 210812
rect 355628 172340 355684 348012
rect 355740 296548 355796 389564
rect 356412 378084 356468 410088
rect 359884 407988 359940 407998
rect 358764 407652 358820 407662
rect 357196 407428 357252 407438
rect 357084 394996 357140 395006
rect 356412 378018 356468 378028
rect 356748 394212 356804 394222
rect 355740 296482 355796 296492
rect 355964 280532 356020 280542
rect 355852 205044 355908 205054
rect 355852 173012 355908 204988
rect 355852 172946 355908 172956
rect 355628 172274 355684 172284
rect 355516 169026 355572 169036
rect 355292 167682 355348 167692
rect 354508 157714 354564 157724
rect 355964 122164 356020 280476
rect 355964 122098 356020 122108
rect 356076 280420 356132 280430
rect 356076 49924 356132 280364
rect 356188 251188 356244 251198
rect 356188 205044 356244 251132
rect 356636 245252 356692 245262
rect 356636 244132 356692 245196
rect 356636 236852 356692 244076
rect 356748 238420 356804 394156
rect 356972 372260 357028 372270
rect 356748 238354 356804 238364
rect 356860 284900 356916 284910
rect 356636 236786 356692 236796
rect 356188 204978 356244 204988
rect 356748 204148 356804 204158
rect 356748 203364 356804 204092
rect 356188 196084 356244 196094
rect 356188 185892 356244 196028
rect 356188 185826 356244 185836
rect 356748 167412 356804 203308
rect 356748 167346 356804 167356
rect 356860 166292 356916 284844
rect 356860 166226 356916 166236
rect 356972 154420 357028 372204
rect 357084 228452 357140 394940
rect 357196 245252 357252 407372
rect 357756 406756 357812 406766
rect 357420 406644 357476 406654
rect 357196 245186 357252 245196
rect 357308 397236 357364 397246
rect 357308 236516 357364 397180
rect 357420 249844 357476 406588
rect 357644 406644 357700 406654
rect 357532 399700 357588 399710
rect 357532 389620 357588 399644
rect 357532 389554 357588 389564
rect 357644 383796 357700 406588
rect 357644 383124 357700 383740
rect 357644 383058 357700 383068
rect 357420 249778 357476 249788
rect 357644 378084 357700 378094
rect 357308 236450 357364 236460
rect 357084 228386 357140 228396
rect 357196 232372 357252 232382
rect 356972 154354 357028 154364
rect 357084 226548 357140 226558
rect 357084 178500 357140 226492
rect 357196 181188 357252 232316
rect 357196 181122 357252 181132
rect 357308 214900 357364 214910
rect 356188 153412 356244 153422
rect 356188 151844 356244 153356
rect 357084 151956 357140 178444
rect 357308 173124 357364 214844
rect 357308 173058 357364 173068
rect 357420 209188 357476 209198
rect 357420 170436 357476 209132
rect 357420 170370 357476 170380
rect 357084 151890 357140 151900
rect 357532 166292 357588 166302
rect 357532 164724 357588 166236
rect 356188 151778 356244 151788
rect 356972 108276 357028 108286
rect 356972 93492 357028 108220
rect 357532 108276 357588 164668
rect 357644 153412 357700 378028
rect 357756 268772 357812 406700
rect 358652 397124 358708 397134
rect 357868 296436 357924 296446
rect 357868 295764 357924 296380
rect 357868 295698 357924 295708
rect 357756 268706 357812 268716
rect 358428 240324 358484 240334
rect 357868 195748 357924 195758
rect 357644 153346 357700 153356
rect 357756 179956 357812 179966
rect 357532 108210 357588 108220
rect 356972 93426 357028 93436
rect 357756 61684 357812 179900
rect 357868 158676 357924 195692
rect 358428 174692 358484 240268
rect 358652 236740 358708 397068
rect 358764 390852 358820 407596
rect 359548 398356 359604 398366
rect 359212 397572 359268 397582
rect 358764 390786 358820 390796
rect 358988 397348 359044 397358
rect 358876 290724 358932 290734
rect 358764 278964 358820 278974
rect 358764 273028 358820 278908
rect 358764 272962 358820 272972
rect 358652 236674 358708 236684
rect 358764 249508 358820 249518
rect 358764 239988 358820 249452
rect 358428 174626 358484 174636
rect 358540 235172 358596 235182
rect 358540 165732 358596 235116
rect 358540 165666 358596 165676
rect 358652 183876 358708 183886
rect 358652 162932 358708 183820
rect 358764 169204 358820 239932
rect 358876 170660 358932 290668
rect 358988 240100 359044 397292
rect 358988 240034 359044 240044
rect 359100 302148 359156 302158
rect 359100 174132 359156 302092
rect 359212 241332 359268 397516
rect 359548 389284 359604 398300
rect 359884 392308 359940 407932
rect 361788 406644 361844 410088
rect 361788 406578 361844 406588
rect 367164 399700 367220 410088
rect 372540 407540 372596 410088
rect 372540 407474 372596 407484
rect 367164 399634 367220 399644
rect 375228 397348 375284 397358
rect 362908 395108 362964 395118
rect 362908 394996 362964 395052
rect 362908 394940 363160 394996
rect 369170 394940 369180 394996
rect 369236 394940 369246 394996
rect 375228 394968 375284 397292
rect 377916 394548 377972 410088
rect 383292 407988 383348 410088
rect 383292 407922 383348 407932
rect 388668 407204 388724 410088
rect 391356 408660 391412 408670
rect 391356 408212 391412 408604
rect 391356 408146 391412 408156
rect 388668 407138 388724 407148
rect 393148 407540 393204 407550
rect 393148 402948 393204 407484
rect 394044 407316 394100 410088
rect 394044 407250 394100 407260
rect 393148 402882 393204 402892
rect 399420 401380 399476 410088
rect 404796 408100 404852 410088
rect 404796 408034 404852 408044
rect 405692 410004 405748 410014
rect 405692 407988 405748 409948
rect 405692 407922 405748 407932
rect 410172 407652 410228 410088
rect 415548 407876 415604 410088
rect 417452 408548 417508 408558
rect 417452 408100 417508 408492
rect 417452 408034 417508 408044
rect 415548 407810 415604 407820
rect 420924 407876 420980 410088
rect 426300 407988 426356 410088
rect 426300 407922 426356 407932
rect 420924 407810 420980 407820
rect 421596 407764 421652 407774
rect 410172 407586 410228 407596
rect 412412 407652 412468 407662
rect 399420 401314 399476 401324
rect 381276 397460 381332 397470
rect 381276 394968 381332 397404
rect 387324 397236 387380 397246
rect 387324 394968 387380 397180
rect 393372 397124 393428 397134
rect 393372 394968 393428 397068
rect 399420 397012 399476 397022
rect 399420 394968 399476 396956
rect 411516 396900 411572 396910
rect 411516 394968 411572 396844
rect 412412 394660 412468 407596
rect 421596 406420 421652 407708
rect 421596 406354 421652 406364
rect 423612 398356 423668 398366
rect 417564 396788 417620 396798
rect 417564 394968 417620 396732
rect 423612 394968 423668 398300
rect 429660 394968 429716 410060
rect 431676 402836 431732 410088
rect 437052 404628 437108 410088
rect 442428 408212 442484 410088
rect 442428 408146 442484 408156
rect 441868 407876 441924 407886
rect 441868 406308 441924 407820
rect 441868 406242 441924 406252
rect 437052 404562 437108 404572
rect 447804 404516 447860 410088
rect 447804 404450 447860 404460
rect 431676 402770 431732 402780
rect 435708 403508 435764 403518
rect 435708 394968 435764 403452
rect 453180 399588 453236 410088
rect 458556 408100 458612 410088
rect 458556 408034 458612 408044
rect 453628 407988 453684 407998
rect 453628 402724 453684 407932
rect 463932 407988 463988 410088
rect 463932 407922 463988 407932
rect 453628 402658 453684 402668
rect 459900 405076 459956 405086
rect 453180 399522 453236 399532
rect 459900 394968 459956 405020
rect 469308 404292 469364 410088
rect 469308 404226 469364 404236
rect 471996 408324 472052 408334
rect 471884 400036 471940 400046
rect 471884 397460 471940 399980
rect 471884 397394 471940 397404
rect 471996 394968 472052 408268
rect 474684 407764 474740 410088
rect 480060 407876 480116 410088
rect 480060 407810 480116 407820
rect 484092 408436 484148 408446
rect 474684 407698 474740 407708
rect 479612 407764 479668 407774
rect 478044 403396 478100 403406
rect 478044 394968 478100 403340
rect 479612 396340 479668 407708
rect 479612 396274 479668 396284
rect 484092 394968 484148 408380
rect 485436 407652 485492 410088
rect 490812 407764 490868 410088
rect 490812 407698 490868 407708
rect 485436 407586 485492 407596
rect 486332 407652 486388 407662
rect 453852 394884 453908 394894
rect 453852 394818 453908 394828
rect 412412 394594 412468 394604
rect 377916 394482 377972 394492
rect 405468 394548 405524 394558
rect 405468 394482 405524 394492
rect 441756 394548 441812 394558
rect 441756 394482 441812 394492
rect 486332 394436 486388 407596
rect 491372 406644 491428 406654
rect 490140 401828 490196 401838
rect 490140 394968 490196 401772
rect 491372 396228 491428 406588
rect 496188 406644 496244 410088
rect 496188 406578 496244 406588
rect 491372 396162 491428 396172
rect 496188 399924 496244 399934
rect 496188 394968 496244 399868
rect 501564 396116 501620 410088
rect 501564 396050 501620 396060
rect 502236 404964 502292 404974
rect 502236 394968 502292 404908
rect 506940 396004 506996 410088
rect 506940 395938 506996 395948
rect 508284 396676 508340 396686
rect 508284 394968 508340 396620
rect 512316 395892 512372 410088
rect 517692 407652 517748 410088
rect 517692 407586 517748 407596
rect 520380 398132 520436 398142
rect 512316 395826 512372 395836
rect 514332 397572 514388 397582
rect 514332 394968 514388 397516
rect 520380 394968 520436 398076
rect 523068 395780 523124 410088
rect 528444 407428 528500 410088
rect 533820 407652 533876 410088
rect 533820 407586 533876 407596
rect 539196 407652 539252 410088
rect 539196 407586 539252 407596
rect 544572 407540 544628 410088
rect 549388 409108 549444 423388
rect 549388 409042 549444 409052
rect 544572 407474 544628 407484
rect 528444 407362 528500 407372
rect 544572 401716 544628 401726
rect 523068 395714 523124 395724
rect 526428 396900 526484 396910
rect 526428 394968 526484 396844
rect 532476 396788 532532 396798
rect 532476 394968 532532 396732
rect 544572 394968 544628 401660
rect 549500 399476 549556 484428
rect 549500 399410 549556 399420
rect 549612 475524 549668 475534
rect 549612 399252 549668 475468
rect 549612 399186 549668 399196
rect 549724 465780 549780 465790
rect 549724 399028 549780 465724
rect 549836 428484 549892 428494
rect 549836 405860 549892 428428
rect 549836 405794 549892 405804
rect 549948 401268 550004 507836
rect 551068 409556 551124 541548
rect 551068 409490 551124 409500
rect 551180 532196 551236 532206
rect 551180 409332 551236 532140
rect 551180 409266 551236 409276
rect 551292 513380 551348 513390
rect 549948 401202 550004 401212
rect 551292 401156 551348 513324
rect 551292 401090 551348 401100
rect 551404 480452 551460 480462
rect 551404 399364 551460 480396
rect 551404 399298 551460 399308
rect 551516 471044 551572 471054
rect 551516 399140 551572 470988
rect 551628 419300 551684 419310
rect 551628 400708 551684 419244
rect 552748 402612 552804 560364
rect 554428 546308 554484 546318
rect 552748 402546 552804 402556
rect 552860 452228 552916 452238
rect 551628 400642 551684 400652
rect 551516 399074 551572 399084
rect 549724 398962 549780 398972
rect 550620 396564 550676 396574
rect 550620 394968 550676 396508
rect 552860 395668 552916 452172
rect 552972 447524 553028 447534
rect 552972 406196 553028 447468
rect 552972 406130 553028 406140
rect 553084 442820 553140 442830
rect 553084 406084 553140 442764
rect 553084 406018 553140 406028
rect 553196 438116 553252 438126
rect 553196 405972 553252 438060
rect 553196 405906 553252 405916
rect 553308 433412 553364 433422
rect 553308 405748 553364 433356
rect 554428 409444 554484 546252
rect 554428 409378 554484 409388
rect 554540 518084 554596 518094
rect 553308 405682 553364 405692
rect 554540 404180 554596 518028
rect 554540 404114 554596 404124
rect 554652 503972 554708 503982
rect 554652 401044 554708 503916
rect 554652 400978 554708 400988
rect 554764 499268 554820 499278
rect 554764 400932 554820 499212
rect 563612 496132 563668 496142
rect 554988 461636 555044 461646
rect 554764 400866 554820 400876
rect 554876 456932 554932 456942
rect 554876 400820 554932 456876
rect 554988 409220 555044 461580
rect 554988 409154 555044 409164
rect 554876 400754 554932 400764
rect 558908 407428 558964 407438
rect 552860 395602 552916 395612
rect 556668 396676 556724 396686
rect 556668 394968 556724 396620
rect 538524 394884 538580 394894
rect 538524 394818 538580 394828
rect 486332 394370 486388 394380
rect 447804 394324 447860 394334
rect 447804 394258 447860 394268
rect 465948 394324 466004 394334
rect 465948 394258 466004 394268
rect 359884 392242 359940 392252
rect 359884 389956 359940 389966
rect 359884 389396 359940 389900
rect 359884 389330 359940 389340
rect 359548 389218 359604 389228
rect 359772 354732 359828 354742
rect 359772 349468 359828 354676
rect 359772 349412 359940 349468
rect 359436 337204 359492 337214
rect 359436 336084 359492 337148
rect 359212 241266 359268 241276
rect 359324 296436 359380 296446
rect 359100 174066 359156 174076
rect 358876 170594 358932 170604
rect 358764 169138 358820 169148
rect 358652 162866 358708 162876
rect 359324 162372 359380 296380
rect 359436 173908 359492 336028
rect 359884 236628 359940 349412
rect 359884 236562 359940 236572
rect 359884 209300 359940 209310
rect 359884 205828 359940 209244
rect 359884 205762 359940 205772
rect 359436 173842 359492 173852
rect 359884 198100 359940 198110
rect 359884 172564 359940 198044
rect 359884 172498 359940 172508
rect 361228 175364 361284 175374
rect 361228 167524 361284 175308
rect 369180 175252 369236 175262
rect 369180 175186 369236 175196
rect 375228 175252 375284 175262
rect 375228 175186 375284 175196
rect 399420 175140 399476 175150
rect 361228 167458 361284 167468
rect 361340 173124 361396 173134
rect 361340 165844 361396 173068
rect 363132 173012 363188 175112
rect 363132 172946 363188 172956
rect 381276 172340 381332 175112
rect 387324 173684 387380 175112
rect 393372 174244 393428 175112
rect 399420 175074 399476 175084
rect 393372 174178 393428 174188
rect 387324 173618 387380 173628
rect 405468 172452 405524 175112
rect 405468 172386 405524 172396
rect 381276 172274 381332 172284
rect 411516 168756 411572 175112
rect 417564 174692 417620 175112
rect 417564 174626 417620 174636
rect 423612 172676 423668 175112
rect 423612 172610 423668 172620
rect 429660 172564 429716 175112
rect 435708 172788 435764 175112
rect 435708 172722 435764 172732
rect 429660 172498 429716 172508
rect 441756 170884 441812 175112
rect 447804 172900 447860 175112
rect 453852 174356 453908 175112
rect 453852 174290 453908 174300
rect 447804 172834 447860 172844
rect 459900 170996 459956 175112
rect 465948 174468 466004 175112
rect 465948 174402 466004 174412
rect 459900 170930 459956 170940
rect 469532 172340 469588 172350
rect 441756 170818 441812 170828
rect 411516 168690 411572 168700
rect 420812 170436 420868 170446
rect 361340 165778 361396 165788
rect 359324 162306 359380 162316
rect 357868 157892 357924 158620
rect 357868 157826 357924 157836
rect 420812 154980 420868 170380
rect 467852 169316 467908 169326
rect 423164 167524 423220 167534
rect 420924 167412 420980 167422
rect 420924 156436 420980 167356
rect 422940 165844 422996 165854
rect 421596 163268 421652 163278
rect 421596 162932 421652 163212
rect 421652 162876 421876 162932
rect 421596 162866 421652 162876
rect 420924 156370 420980 156380
rect 421708 162596 421764 162606
rect 421708 156324 421764 162540
rect 421708 156258 421764 156268
rect 420812 154914 420868 154924
rect 421708 151956 421764 151966
rect 417116 143668 417172 143678
rect 405020 133924 405076 133934
rect 378812 130452 378868 130462
rect 376796 127428 376852 127438
rect 362684 124292 362740 124302
rect 362684 119896 362740 124236
rect 370748 124180 370804 124190
rect 368732 124068 368788 124078
rect 364700 123956 364756 123966
rect 364700 119896 364756 123900
rect 366716 123396 366772 123406
rect 366716 119896 366772 123340
rect 368732 119896 368788 124012
rect 370748 119896 370804 124124
rect 374780 123732 374836 123742
rect 372764 123620 372820 123630
rect 372764 119896 372820 123564
rect 374780 119896 374836 123676
rect 376796 119896 376852 127372
rect 378812 119896 378868 130396
rect 400988 130340 401044 130350
rect 392924 127316 392980 127326
rect 382844 123844 382900 123854
rect 380828 123508 380884 123518
rect 380828 119896 380884 123452
rect 382844 119896 382900 123788
rect 384860 122724 384916 122734
rect 384860 119896 384916 122668
rect 386876 122724 386932 122734
rect 386876 119896 386932 122668
rect 388892 122724 388948 122734
rect 388892 119896 388948 122668
rect 390908 122724 390964 122734
rect 390908 119896 390964 122668
rect 392924 119896 392980 127260
rect 396956 127204 397012 127214
rect 394940 122724 394996 122734
rect 394940 119896 394996 122668
rect 396956 119896 397012 127148
rect 398972 127092 399028 127102
rect 398972 119896 399028 127036
rect 400988 119896 401044 130284
rect 403004 130228 403060 130238
rect 403004 119896 403060 130172
rect 405020 119896 405076 133868
rect 407036 133812 407092 133822
rect 407036 119896 407092 133756
rect 409052 133700 409108 133710
rect 409052 119896 409108 133644
rect 411068 133588 411124 133598
rect 411068 119896 411124 133532
rect 413084 122724 413140 122734
rect 413084 119896 413140 122668
rect 414988 122724 415044 122734
rect 414988 119924 415044 122668
rect 414988 119868 415128 119924
rect 417116 119896 417172 143612
rect 420140 95284 420196 95294
rect 420140 90748 420196 95228
rect 356076 49858 356132 49868
rect 356188 51940 356244 51950
rect 356188 48692 356244 51884
rect 357756 51940 357812 61628
rect 420028 90692 420196 90748
rect 357756 51874 357812 51884
rect 419244 53060 419300 53070
rect 419244 50708 419300 53004
rect 420028 52836 420084 90692
rect 420028 52770 420084 52780
rect 420140 88340 420196 88350
rect 419244 50642 419300 50652
rect 420140 50596 420196 88284
rect 421708 81396 421764 151900
rect 421820 95284 421876 162876
rect 422492 156436 422548 156446
rect 422492 154196 422548 156380
rect 421932 119364 421988 119374
rect 421932 102452 421988 119308
rect 421932 102386 421988 102396
rect 421820 95218 421876 95228
rect 421708 78988 421764 81340
rect 421708 78932 422100 78988
rect 420140 50530 420196 50540
rect 420252 74452 420308 74462
rect 420252 49700 420308 74396
rect 421820 68852 421876 68862
rect 421820 67508 421876 68796
rect 421820 49812 421876 67452
rect 421932 60564 421988 60574
rect 421932 50484 421988 60508
rect 421932 50418 421988 50428
rect 421820 49746 421876 49756
rect 420252 49634 420308 49644
rect 422044 49588 422100 78932
rect 422492 53620 422548 154140
rect 422604 156324 422660 156334
rect 422604 88340 422660 156268
rect 422604 88274 422660 88284
rect 422716 154980 422772 154990
rect 422716 154084 422772 154924
rect 422716 60564 422772 154028
rect 422940 153972 422996 165788
rect 422940 68852 422996 153916
rect 423164 153860 423220 167468
rect 423164 74452 423220 153804
rect 466284 162484 466340 162494
rect 466284 154196 466340 162428
rect 423276 153300 423332 153310
rect 423276 151956 423332 153244
rect 423276 151890 423332 151900
rect 459452 151284 459508 151294
rect 457996 122164 458052 122174
rect 457884 120372 457940 120382
rect 457772 117012 457828 117022
rect 457772 92708 457828 116956
rect 457884 101444 457940 120316
rect 457996 107268 458052 122108
rect 458220 122052 458276 122062
rect 458108 120260 458164 120270
rect 458108 113092 458164 120204
rect 458108 113026 458164 113036
rect 458220 110180 458276 121996
rect 458220 110114 458276 110124
rect 458556 117572 458612 117582
rect 457996 107202 458052 107212
rect 458556 104356 458612 117516
rect 458556 104290 458612 104300
rect 459452 102452 459508 151228
rect 466284 149912 466340 154140
rect 467852 154084 467908 169260
rect 467852 149940 467908 154028
rect 467656 149884 467908 149940
rect 468972 164388 469028 164398
rect 468972 153972 469028 164332
rect 468972 149912 469028 153916
rect 469532 153860 469588 172284
rect 471996 171108 472052 175112
rect 471996 171042 472052 171052
rect 478044 169428 478100 175112
rect 484092 171220 484148 175112
rect 484092 171154 484148 171164
rect 489132 174132 489188 174142
rect 478044 169362 478100 169372
rect 486444 170660 486500 170670
rect 483756 169204 483812 169214
rect 482412 165732 482468 165742
rect 477036 164948 477092 164958
rect 474348 163268 474404 163278
rect 473004 156324 473060 156334
rect 473004 154532 473060 156268
rect 469532 149940 469588 153804
rect 471660 153860 471716 153870
rect 471660 153300 471716 153804
rect 469532 149884 470344 149940
rect 471660 149912 471716 153244
rect 473004 149912 473060 154476
rect 474348 154420 474404 163212
rect 474348 149912 474404 154364
rect 475692 151284 475748 151294
rect 475692 149912 475748 151228
rect 477036 149912 477092 164892
rect 478380 164836 478436 164846
rect 478380 149912 478436 164780
rect 479724 163156 479780 163166
rect 479724 149912 479780 163100
rect 482412 149912 482468 165676
rect 483756 149912 483812 169148
rect 485100 164724 485156 164734
rect 485100 149912 485156 164668
rect 486444 149912 486500 170604
rect 487788 162372 487844 162382
rect 487788 149912 487844 162316
rect 489132 149912 489188 174076
rect 490140 172116 490196 175112
rect 490140 172050 490196 172060
rect 495852 174020 495908 174030
rect 494508 170548 494564 170558
rect 491820 154308 491876 154318
rect 490476 154084 490532 154094
rect 490476 149912 490532 154028
rect 491820 149912 491876 154252
rect 493164 153300 493220 153310
rect 493164 149912 493220 153244
rect 494508 149912 494564 170492
rect 495852 149912 495908 173964
rect 496188 169540 496244 175112
rect 496188 169474 496244 169484
rect 497196 173908 497252 173918
rect 497196 149912 497252 173852
rect 502236 167636 502292 175112
rect 508284 167748 508340 175112
rect 514332 169652 514388 175112
rect 520380 174580 520436 175112
rect 520380 174514 520436 174524
rect 514332 169586 514388 169596
rect 508284 167682 508340 167692
rect 516012 169092 516068 169102
rect 502236 167570 502292 167580
rect 498540 166404 498596 166414
rect 498540 149912 498596 166348
rect 510636 164276 510692 164286
rect 499884 163044 499940 163054
rect 499884 149912 499940 162988
rect 503916 155988 503972 155998
rect 503916 153972 503972 155932
rect 503916 153906 503972 153916
rect 505260 153748 505316 153758
rect 503916 153300 503972 153310
rect 502572 152964 502628 152974
rect 502572 149912 502628 152908
rect 503132 152964 503188 152974
rect 481068 149828 481124 149838
rect 503132 149828 503188 152908
rect 503916 150948 503972 153244
rect 503916 150882 503972 150892
rect 505260 149912 505316 153692
rect 509292 153636 509348 153646
rect 506604 153412 506660 153422
rect 505596 153188 505652 153198
rect 505596 152852 505652 153132
rect 505596 152786 505652 152796
rect 506604 149912 506660 153356
rect 506828 153412 506884 153422
rect 506828 150276 506884 153356
rect 506828 150210 506884 150220
rect 507948 153076 508004 153086
rect 507948 149912 508004 153020
rect 508172 153076 508228 153086
rect 508172 150836 508228 153020
rect 508172 150770 508228 150780
rect 509292 149912 509348 153580
rect 510636 149912 510692 164220
rect 511980 161812 512036 161822
rect 511980 149912 512036 161756
rect 513324 159348 513380 159358
rect 513324 149912 513380 159292
rect 514668 152292 514724 152302
rect 514668 149912 514724 152236
rect 516012 149912 516068 169036
rect 526428 167860 526484 175112
rect 532476 171332 532532 175112
rect 538524 173012 538580 175112
rect 538524 172946 538580 172956
rect 544572 172900 544628 175112
rect 550620 173012 550676 175112
rect 550620 172946 550676 172956
rect 544572 172834 544628 172844
rect 556668 172900 556724 175112
rect 556668 172834 556724 172844
rect 532476 171266 532532 171276
rect 526428 167794 526484 167804
rect 524076 164164 524132 164174
rect 521388 160692 521444 160702
rect 520044 160356 520100 160366
rect 518700 160244 518756 160254
rect 517356 159908 517412 159918
rect 517356 149912 517412 159852
rect 518700 149912 518756 160188
rect 520044 149912 520100 160300
rect 521388 149912 521444 160636
rect 522732 160580 522788 160590
rect 522732 149912 522788 160524
rect 524076 149912 524132 164108
rect 546588 161924 546644 161934
rect 524188 159460 524244 159470
rect 524188 153748 524244 159404
rect 540876 159124 540932 159134
rect 524188 153682 524244 153692
rect 526764 156212 526820 156222
rect 525420 153300 525476 153310
rect 525420 149912 525476 153244
rect 526764 149912 526820 156156
rect 530796 156100 530852 156110
rect 528108 155876 528164 155886
rect 528108 149912 528164 155820
rect 529452 155764 529508 155774
rect 529452 149912 529508 155708
rect 530796 149912 530852 156044
rect 537516 155540 537572 155550
rect 532140 153972 532196 153982
rect 532140 149912 532196 153916
rect 534828 153188 534884 153198
rect 532588 152964 532644 152974
rect 532588 151060 532644 152908
rect 532588 150994 532644 151004
rect 533484 152404 533540 152414
rect 533484 149912 533540 152348
rect 534828 149912 534884 153132
rect 537516 149912 537572 155484
rect 540876 154084 540932 159068
rect 544348 159012 544404 159022
rect 540876 154018 540932 154028
rect 544236 155652 544292 155662
rect 542892 153412 542948 153422
rect 540204 153076 540260 153086
rect 538860 152180 538916 152190
rect 538860 149912 538916 152124
rect 540204 149912 540260 153020
rect 541548 152964 541604 152974
rect 541548 149912 541604 152908
rect 542892 149912 542948 153356
rect 544236 149912 544292 155596
rect 544348 154308 544404 158956
rect 544348 154242 544404 154252
rect 546588 154196 546644 161868
rect 549612 159236 549668 159246
rect 546588 154130 546644 154140
rect 548268 158900 548324 158910
rect 546924 154084 546980 154094
rect 545580 153748 545636 153758
rect 545580 149912 545636 153692
rect 546924 149912 546980 154028
rect 548268 149912 548324 158844
rect 549612 149912 549668 159180
rect 558908 154420 558964 407372
rect 559468 403284 559524 403294
rect 559020 392420 559076 392430
rect 559020 391524 559076 392364
rect 559020 172340 559076 391468
rect 559020 172274 559076 172284
rect 559468 154532 559524 403228
rect 563612 402500 563668 496076
rect 587132 443268 587188 443278
rect 583772 416836 583828 416846
rect 583772 404068 583828 416780
rect 587132 407428 587188 443212
rect 587132 407362 587188 407372
rect 583772 404002 583828 404012
rect 563612 402434 563668 402444
rect 559468 154466 559524 154476
rect 559580 397460 559636 397470
rect 559580 396564 559636 397404
rect 558908 154354 558964 154364
rect 550956 154308 551012 154318
rect 550956 149912 551012 154252
rect 552300 154196 552356 154206
rect 552300 149912 552356 154140
rect 559580 153860 559636 396508
rect 590604 396564 590660 396574
rect 566972 394772 567028 394782
rect 562828 393428 562884 393438
rect 559692 393316 559748 393326
rect 559692 172788 559748 393260
rect 559692 172722 559748 172732
rect 560252 205380 560308 205390
rect 560252 162484 560308 205324
rect 562828 173012 562884 393372
rect 566972 337540 567028 394716
rect 566972 337474 567028 337484
rect 578732 393204 578788 393214
rect 578732 297892 578788 393148
rect 578732 297826 578788 297836
rect 590492 392644 590548 392654
rect 562828 172946 562884 172956
rect 565292 284676 565348 284686
rect 565292 164388 565348 284620
rect 590492 258468 590548 392588
rect 590604 364196 590660 396508
rect 590940 392308 590996 392318
rect 590604 364130 590660 364140
rect 590716 391524 590772 391534
rect 590716 324548 590772 391468
rect 590940 350980 590996 392252
rect 590940 350914 590996 350924
rect 590716 324482 590772 324492
rect 590492 258402 590548 258412
rect 587132 245028 587188 245038
rect 587132 169316 587188 244972
rect 587132 169250 587188 169260
rect 565292 164322 565348 164332
rect 560252 162418 560308 162428
rect 560364 162148 560420 162158
rect 560140 157892 560196 157902
rect 559916 157556 559972 157566
rect 559804 157444 559860 157454
rect 559580 153794 559636 153804
rect 559692 157220 559748 157230
rect 552636 150724 552692 150734
rect 552692 150668 552916 150724
rect 552636 150658 552692 150668
rect 552860 149940 552916 150668
rect 552860 149884 553672 149940
rect 503132 149772 503944 149828
rect 481068 149762 481124 149772
rect 536172 149604 536228 149614
rect 536172 149538 536228 149548
rect 501228 149268 501284 149278
rect 501228 149202 501284 149212
rect 559468 149268 559524 149278
rect 559468 118468 559524 149212
rect 559580 148708 559636 148718
rect 559580 124404 559636 148652
rect 559692 142100 559748 157164
rect 559692 142034 559748 142044
rect 559804 132580 559860 157388
rect 559916 134372 559972 157500
rect 560028 157108 560084 157118
rect 560028 140644 560084 157052
rect 560028 140578 560084 140588
rect 560140 135156 560196 157836
rect 560252 157668 560308 157678
rect 560252 136724 560308 157612
rect 560252 136658 560308 136668
rect 560140 135090 560196 135100
rect 559916 134306 559972 134316
rect 559804 132514 559860 132524
rect 559580 124338 559636 124348
rect 559468 118402 559524 118412
rect 560364 111636 560420 162092
rect 564508 162036 564564 162046
rect 561372 158788 561428 158798
rect 561148 157780 561204 157790
rect 561148 138292 561204 157724
rect 561260 149492 561316 149502
rect 561260 142996 561316 149436
rect 561260 142930 561316 142940
rect 561148 138226 561204 138236
rect 561372 127316 561428 158732
rect 561596 152068 561652 152078
rect 561372 127250 561428 127260
rect 561484 150388 561540 150398
rect 560364 111570 560420 111580
rect 561484 108500 561540 150332
rect 561596 114772 561652 152012
rect 563164 150612 563220 150622
rect 561596 114706 561652 114716
rect 562828 149716 562884 149726
rect 561484 108434 561540 108444
rect 459452 102386 459508 102396
rect 457884 101378 457940 101388
rect 457772 92642 457828 92652
rect 423164 74386 423220 74396
rect 562828 70868 562884 149660
rect 562940 148932 562996 148942
rect 562940 80276 562996 148876
rect 563052 148820 563108 148830
rect 563052 86548 563108 148764
rect 563164 88116 563220 150556
rect 564508 122612 564564 161980
rect 566188 160468 566244 160478
rect 564732 157332 564788 157342
rect 564508 122546 564564 122556
rect 564620 155428 564676 155438
rect 564620 119476 564676 155372
rect 564732 130452 564788 157276
rect 564732 130386 564788 130396
rect 566188 128884 566244 160412
rect 566188 128818 566244 128828
rect 564620 119410 564676 119420
rect 563164 88050 563220 88060
rect 563052 86482 563108 86492
rect 562940 80210 562996 80220
rect 563500 81844 563556 81854
rect 562828 70802 562884 70812
rect 563388 72436 563444 72446
rect 422940 68786 422996 68796
rect 422716 60498 422772 60508
rect 563164 67732 563220 67742
rect 562940 59892 562996 59902
rect 422492 53554 422548 53564
rect 562828 58324 562884 58334
rect 562828 49924 562884 58268
rect 562828 49858 562884 49868
rect 422044 49522 422100 49532
rect 356188 48626 356244 48636
rect 562940 48356 562996 59836
rect 562940 48290 562996 48300
rect 354396 48178 354452 48188
rect 563164 48244 563220 67676
rect 563276 63028 563332 63038
rect 563276 50372 563332 62972
rect 563276 50306 563332 50316
rect 563388 48580 563444 72380
rect 563388 48514 563444 48524
rect 563164 48178 563220 48188
rect 563500 45332 563556 81788
rect 563724 69300 563780 69310
rect 563612 61460 563668 61470
rect 563612 48020 563668 61404
rect 563724 48468 563780 69244
rect 563724 48402 563780 48412
rect 563612 47954 563668 47964
rect 563500 45266 563556 45276
rect 289996 24322 290052 24332
rect 289772 4610 289828 4620
rect 277340 4050 277396 4060
rect 580636 4228 580692 4238
rect 580636 480 580692 4172
rect 582540 4228 582596 4238
rect 582540 480 582596 4172
rect 584444 4228 584500 4238
rect 584444 480 584500 4172
rect 207452 392 207704 480
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 392 209636 480
rect 211288 392 211540 480
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 213192 -960 213416 480
rect 215096 -960 215320 480
rect 217000 -960 217224 480
rect 218904 -960 219128 480
rect 220808 -960 221032 480
rect 222712 -960 222936 480
rect 224616 -960 224840 480
rect 226520 -960 226744 480
rect 228424 -960 228648 480
rect 230328 -960 230552 480
rect 232232 -960 232456 480
rect 234136 -960 234360 480
rect 236040 -960 236264 480
rect 237944 -960 238168 480
rect 239848 -960 240072 480
rect 241752 -960 241976 480
rect 243656 -960 243880 480
rect 245560 -960 245784 480
rect 247464 -960 247688 480
rect 249368 -960 249592 480
rect 251272 -960 251496 480
rect 253176 -960 253400 480
rect 255080 -960 255304 480
rect 256984 -960 257208 480
rect 258888 -960 259112 480
rect 260792 -960 261016 480
rect 262696 -960 262920 480
rect 264600 -960 264824 480
rect 266504 -960 266728 480
rect 268408 -960 268632 480
rect 270312 -960 270536 480
rect 272216 -960 272440 480
rect 274120 -960 274344 480
rect 276024 -960 276248 480
rect 277928 -960 278152 480
rect 279832 -960 280056 480
rect 281736 -960 281960 480
rect 283640 -960 283864 480
rect 285544 -960 285768 480
rect 287448 -960 287672 480
rect 289352 -960 289576 480
rect 291256 -960 291480 480
rect 293160 -960 293384 480
rect 295064 -960 295288 480
rect 296968 -960 297192 480
rect 298872 -960 299096 480
rect 300776 -960 301000 480
rect 302680 -960 302904 480
rect 304584 -960 304808 480
rect 306488 -960 306712 480
rect 308392 -960 308616 480
rect 310296 -960 310520 480
rect 312200 -960 312424 480
rect 314104 -960 314328 480
rect 316008 -960 316232 480
rect 317912 -960 318136 480
rect 319816 -960 320040 480
rect 321720 -960 321944 480
rect 323624 -960 323848 480
rect 325528 -960 325752 480
rect 327432 -960 327656 480
rect 329336 -960 329560 480
rect 331240 -960 331464 480
rect 333144 -960 333368 480
rect 335048 -960 335272 480
rect 336952 -960 337176 480
rect 338856 -960 339080 480
rect 340760 -960 340984 480
rect 342664 -960 342888 480
rect 344568 -960 344792 480
rect 346472 -960 346696 480
rect 348376 -960 348600 480
rect 350280 -960 350504 480
rect 352184 -960 352408 480
rect 354088 -960 354312 480
rect 355992 -960 356216 480
rect 357896 -960 358120 480
rect 359800 -960 360024 480
rect 361704 -960 361928 480
rect 363608 -960 363832 480
rect 365512 -960 365736 480
rect 367416 -960 367640 480
rect 369320 -960 369544 480
rect 371224 -960 371448 480
rect 373128 -960 373352 480
rect 375032 -960 375256 480
rect 376936 -960 377160 480
rect 378840 -960 379064 480
rect 380744 -960 380968 480
rect 382648 -960 382872 480
rect 384552 -960 384776 480
rect 386456 -960 386680 480
rect 388360 -960 388584 480
rect 390264 -960 390488 480
rect 392168 -960 392392 480
rect 394072 -960 394296 480
rect 395976 -960 396200 480
rect 397880 -960 398104 480
rect 399784 -960 400008 480
rect 401688 -960 401912 480
rect 403592 -960 403816 480
rect 405496 -960 405720 480
rect 407400 -960 407624 480
rect 409304 -960 409528 480
rect 411208 -960 411432 480
rect 413112 -960 413336 480
rect 415016 -960 415240 480
rect 416920 -960 417144 480
rect 418824 -960 419048 480
rect 420728 -960 420952 480
rect 422632 -960 422856 480
rect 424536 -960 424760 480
rect 426440 -960 426664 480
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432152 -960 432376 480
rect 434056 -960 434280 480
rect 435960 -960 436184 480
rect 437864 -960 438088 480
rect 439768 -960 439992 480
rect 441672 -960 441896 480
rect 443576 -960 443800 480
rect 445480 -960 445704 480
rect 447384 -960 447608 480
rect 449288 -960 449512 480
rect 451192 -960 451416 480
rect 453096 -960 453320 480
rect 455000 -960 455224 480
rect 456904 -960 457128 480
rect 458808 -960 459032 480
rect 460712 -960 460936 480
rect 462616 -960 462840 480
rect 464520 -960 464744 480
rect 466424 -960 466648 480
rect 468328 -960 468552 480
rect 470232 -960 470456 480
rect 472136 -960 472360 480
rect 474040 -960 474264 480
rect 475944 -960 476168 480
rect 477848 -960 478072 480
rect 479752 -960 479976 480
rect 481656 -960 481880 480
rect 483560 -960 483784 480
rect 485464 -960 485688 480
rect 487368 -960 487592 480
rect 489272 -960 489496 480
rect 491176 -960 491400 480
rect 493080 -960 493304 480
rect 494984 -960 495208 480
rect 496888 -960 497112 480
rect 498792 -960 499016 480
rect 500696 -960 500920 480
rect 502600 -960 502824 480
rect 504504 -960 504728 480
rect 506408 -960 506632 480
rect 508312 -960 508536 480
rect 510216 -960 510440 480
rect 512120 -960 512344 480
rect 514024 -960 514248 480
rect 515928 -960 516152 480
rect 517832 -960 518056 480
rect 519736 -960 519960 480
rect 521640 -960 521864 480
rect 523544 -960 523768 480
rect 525448 -960 525672 480
rect 527352 -960 527576 480
rect 529256 -960 529480 480
rect 531160 -960 531384 480
rect 533064 -960 533288 480
rect 534968 -960 535192 480
rect 536872 -960 537096 480
rect 538776 -960 539000 480
rect 540680 -960 540904 480
rect 542584 -960 542808 480
rect 544488 -960 544712 480
rect 546392 -960 546616 480
rect 548296 -960 548520 480
rect 550200 -960 550424 480
rect 552104 -960 552328 480
rect 554008 -960 554232 480
rect 555912 -960 556136 480
rect 557816 -960 558040 480
rect 559720 -960 559944 480
rect 561624 -960 561848 480
rect 563528 -960 563752 480
rect 565432 -960 565656 480
rect 567336 -960 567560 480
rect 569240 -960 569464 480
rect 571144 -960 571368 480
rect 573048 -960 573272 480
rect 574952 -960 575176 480
rect 576856 -960 577080 480
rect 578760 -960 578984 480
rect 580636 392 580888 480
rect 582540 392 582792 480
rect 584444 392 584696 480
rect 580664 -960 580888 392
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 4172 388108 4228 388164
rect 4172 333340 4228 333396
rect 12572 573020 12628 573076
rect 14252 530684 14308 530740
rect 14252 397292 14308 397348
rect 15932 488348 15988 488404
rect 12572 395612 12628 395668
rect 15932 393932 15988 393988
rect 99484 590492 99540 590548
rect 77308 572012 77364 572068
rect 121324 570332 121380 570388
rect 141932 590492 141988 590548
rect 57932 544796 57988 544852
rect 56252 502460 56308 502516
rect 56252 409836 56308 409892
rect 57932 409724 57988 409780
rect 55132 409164 55188 409220
rect 33068 392252 33124 392308
rect 103404 407372 103460 407428
rect 99932 386652 99988 386708
rect 38556 386540 38612 386596
rect 38444 386428 38500 386484
rect 11004 301532 11060 301588
rect 12572 383068 12628 383124
rect 4172 290780 4228 290836
rect 32732 380156 32788 380212
rect 29372 380044 29428 380100
rect 27692 379932 27748 379988
rect 20972 379820 21028 379876
rect 12572 276668 12628 276724
rect 14252 379260 14308 379316
rect 4172 239372 4228 239428
rect 13244 229404 13300 229460
rect 4172 208684 4228 208740
rect 4172 121660 4228 121716
rect 11340 47852 11396 47908
rect 14252 191996 14308 192052
rect 20860 229292 20916 229348
rect 14252 79100 14308 79156
rect 14252 50316 14308 50372
rect 15372 4172 15428 4228
rect 17276 4172 17332 4228
rect 19180 4172 19236 4228
rect 20972 64988 21028 65044
rect 22764 232652 22820 232708
rect 26572 222572 26628 222628
rect 25116 4172 25172 4228
rect 29372 107324 29428 107380
rect 30380 227612 30436 227668
rect 27692 22652 27748 22708
rect 32284 214172 32340 214228
rect 38332 379484 38388 379540
rect 40908 383964 40964 384020
rect 40684 379372 40740 379428
rect 38556 238476 38612 238532
rect 40236 378588 40292 378644
rect 40236 238364 40292 238420
rect 38444 238252 38500 238308
rect 38332 238140 38388 238196
rect 41132 380716 41188 380772
rect 62412 303996 62468 304052
rect 47404 302428 47460 302484
rect 77420 303996 77476 304052
rect 92428 303996 92484 304052
rect 60844 240716 60900 240772
rect 74956 240716 75012 240772
rect 64876 240492 64932 240548
rect 62860 240380 62916 240436
rect 66892 240268 66948 240324
rect 68908 240156 68964 240212
rect 46732 238476 46788 238532
rect 52780 238364 52836 238420
rect 50764 238252 50820 238308
rect 48748 238140 48804 238196
rect 40684 237916 40740 237972
rect 56812 240044 56868 240100
rect 58828 239820 58884 239876
rect 54796 237916 54852 237972
rect 72940 238476 72996 238532
rect 76972 238476 77028 238532
rect 81004 239708 81060 239764
rect 78988 237916 79044 237972
rect 87052 238140 87108 238196
rect 85036 238028 85092 238084
rect 83020 237804 83076 237860
rect 91084 238476 91140 238532
rect 95116 238476 95172 238532
rect 103292 385084 103348 385140
rect 100380 384972 100436 385028
rect 99932 238476 99988 238532
rect 100156 384748 100212 384804
rect 97132 238364 97188 238420
rect 93100 238252 93156 238308
rect 89068 237692 89124 237748
rect 96572 238140 96628 238196
rect 143388 410732 143444 410788
rect 186396 590492 186452 590548
rect 179004 587132 179060 587188
rect 175532 572012 175588 572068
rect 172172 570332 172228 570388
rect 172172 408044 172228 408100
rect 173852 446012 173908 446068
rect 173852 398972 173908 399028
rect 165452 392364 165508 392420
rect 141932 390684 141988 390740
rect 111692 386764 111748 386820
rect 103404 284396 103460 284452
rect 103516 384860 103572 384916
rect 106652 383292 106708 383348
rect 104972 379036 105028 379092
rect 103628 286524 103684 286580
rect 103628 272748 103684 272804
rect 103516 238140 103572 238196
rect 103292 237916 103348 237972
rect 100380 237804 100436 237860
rect 100156 237692 100212 237748
rect 96572 237580 96628 237636
rect 106652 238364 106708 238420
rect 118412 383516 118468 383572
rect 115052 382060 115108 382116
rect 113372 321804 113428 321860
rect 113372 278572 113428 278628
rect 115164 320124 115220 320180
rect 115164 261100 115220 261156
rect 115052 239820 115108 239876
rect 111692 238252 111748 238308
rect 126812 381724 126868 381780
rect 120092 381612 120148 381668
rect 120092 239932 120148 239988
rect 125132 381500 125188 381556
rect 125244 378924 125300 378980
rect 125244 319004 125300 319060
rect 126812 241052 126868 241108
rect 130172 380268 130228 380324
rect 125132 239708 125188 239764
rect 118412 238028 118468 238084
rect 104972 237580 105028 237636
rect 70924 235116 70980 235172
rect 130284 378700 130340 378756
rect 130284 361340 130340 361396
rect 140252 322028 140308 322084
rect 168028 322028 168084 322084
rect 152796 321916 152852 321972
rect 143612 321692 143668 321748
rect 143612 302428 143668 302484
rect 143612 288988 143668 289044
rect 151116 288876 151172 288932
rect 168028 321580 168084 321636
rect 173964 301532 174020 301588
rect 161308 299852 161364 299908
rect 169148 289772 169204 289828
rect 168812 286636 168868 286692
rect 151228 285292 151284 285348
rect 165452 285292 165508 285348
rect 165452 278796 165508 278852
rect 169148 283948 169204 284004
rect 168812 277900 168868 277956
rect 174636 278796 174692 278852
rect 174636 275996 174692 276052
rect 173964 272972 174020 273028
rect 178892 414540 178948 414596
rect 177324 410732 177380 410788
rect 176316 360332 176372 360388
rect 175532 271628 175588 271684
rect 175980 337484 176036 337540
rect 140252 266924 140308 266980
rect 174636 268716 174692 268772
rect 174636 267148 174692 267204
rect 174636 239932 174692 239988
rect 130172 234332 130228 234388
rect 175980 232988 176036 233044
rect 176092 333452 176148 333508
rect 40236 229516 40292 229572
rect 38556 224364 38612 224420
rect 37996 222796 38052 222852
rect 32732 149660 32788 149716
rect 33516 210812 33572 210868
rect 33516 4396 33572 4452
rect 34412 4172 34468 4228
rect 38444 219212 38500 219268
rect 38332 214396 38388 214452
rect 38332 4172 38388 4228
rect 38556 4956 38612 5012
rect 39900 222684 39956 222740
rect 38444 4060 38500 4116
rect 176092 221004 176148 221060
rect 176204 329420 176260 329476
rect 176428 346220 176484 346276
rect 176428 286524 176484 286580
rect 177212 275996 177268 276052
rect 177996 357644 178052 357700
rect 177324 270284 177380 270340
rect 177884 338828 177940 338884
rect 177212 265468 177268 265524
rect 177884 234108 177940 234164
rect 178556 342860 178612 342916
rect 178332 336028 178388 336084
rect 178220 332780 178276 332836
rect 178220 249452 178276 249508
rect 178444 330092 178500 330148
rect 184716 578732 184772 578788
rect 179004 409276 179060 409332
rect 180460 577052 180516 577108
rect 179228 403676 179284 403732
rect 179004 390908 179060 390964
rect 179228 390796 179284 390852
rect 179676 362908 179732 362964
rect 179452 356188 179508 356244
rect 179004 342860 179060 342916
rect 179116 354396 179172 354452
rect 179116 336028 179172 336084
rect 178892 321692 178948 321748
rect 178556 321580 178612 321636
rect 178332 255276 178388 255332
rect 179004 249452 179060 249508
rect 178892 224700 178948 224756
rect 177996 224588 178052 224644
rect 179116 243628 179172 243684
rect 179452 232764 179508 232820
rect 179564 350924 179620 350980
rect 179116 231308 179172 231364
rect 183932 460124 183988 460180
rect 181468 417788 181524 417844
rect 181468 409500 181524 409556
rect 183932 409388 183988 409444
rect 182476 407596 182532 407652
rect 180908 397404 180964 397460
rect 180796 395724 180852 395780
rect 180684 385420 180740 385476
rect 180460 262220 180516 262276
rect 180572 380380 180628 380436
rect 182364 394156 182420 394212
rect 182252 379708 182308 379764
rect 182252 379484 182308 379540
rect 182252 369740 182308 369796
rect 181244 361676 181300 361732
rect 181132 352268 181188 352324
rect 180908 346220 180964 346276
rect 181020 349580 181076 349636
rect 180796 322700 180852 322756
rect 180908 344204 180964 344260
rect 180684 240716 180740 240772
rect 180572 235116 180628 235172
rect 179676 234668 179732 234724
rect 181020 234780 181076 234836
rect 180908 232876 180964 232932
rect 181132 229628 181188 229684
rect 184044 394044 184100 394100
rect 183932 385532 183988 385588
rect 182476 354396 182532 354452
rect 183820 368396 183876 368452
rect 183036 353612 183092 353668
rect 182812 348236 182868 348292
rect 182364 330204 182420 330260
rect 182588 334796 182644 334852
rect 182252 299852 182308 299908
rect 181356 272076 181412 272132
rect 181468 265468 181524 265524
rect 181468 255388 181524 255444
rect 181356 240604 181412 240660
rect 182588 239484 182644 239540
rect 182700 330764 182756 330820
rect 182700 229852 182756 229908
rect 182812 227836 182868 227892
rect 182924 341516 182980 341572
rect 181244 227724 181300 227780
rect 179564 223020 179620 223076
rect 179004 222908 179060 222964
rect 176316 220892 176372 220948
rect 176204 217756 176260 217812
rect 154924 217644 154980 217700
rect 40236 4620 40292 4676
rect 41132 215852 41188 215908
rect 183820 322252 183876 322308
rect 184044 332780 184100 332836
rect 184156 380492 184212 380548
rect 184604 365708 184660 365764
rect 184492 345548 184548 345604
rect 184380 332108 184436 332164
rect 184156 240492 184212 240548
rect 184268 328076 184324 328132
rect 183932 240268 183988 240324
rect 183036 219324 183092 219380
rect 184492 224812 184548 224868
rect 184380 219436 184436 219492
rect 184268 217868 184324 217924
rect 182924 217644 182980 217700
rect 186284 565068 186340 565124
rect 186172 550732 186228 550788
rect 186060 543564 186116 543620
rect 186060 388892 186116 388948
rect 187180 514892 187236 514948
rect 187180 408940 187236 408996
rect 187292 507724 187348 507780
rect 186396 404124 186452 404180
rect 186284 390572 186340 390628
rect 186172 387212 186228 387268
rect 186396 358988 186452 359044
rect 186284 346892 186340 346948
rect 186172 340172 186228 340228
rect 185612 283836 185668 283892
rect 184716 263564 184772 263620
rect 185724 273868 185780 273924
rect 185612 255388 185668 255444
rect 185612 243516 185668 243572
rect 185724 240492 185780 240548
rect 186284 231084 186340 231140
rect 186172 227948 186228 228004
rect 186508 296492 186564 296548
rect 189644 591276 189700 591332
rect 189196 590940 189252 590996
rect 189084 575372 189140 575428
rect 187852 557900 187908 557956
rect 187516 487228 187572 487284
rect 187740 536396 187796 536452
rect 187292 289772 187348 289828
rect 187404 471884 187460 471940
rect 186508 286636 186564 286692
rect 187180 285628 187236 285684
rect 187628 464716 187684 464772
rect 187404 283836 187460 283892
rect 187516 450380 187572 450436
rect 188076 493388 188132 493444
rect 187852 410396 187908 410452
rect 187964 443212 188020 443268
rect 187740 409612 187796 409668
rect 187852 295596 187908 295652
rect 187852 285740 187908 285796
rect 187628 283612 187684 283668
rect 188860 487228 188916 487284
rect 189084 407932 189140 407988
rect 188860 407820 188916 407876
rect 189196 407484 189252 407540
rect 189308 590716 189364 590772
rect 189532 572012 189588 572068
rect 189308 405692 189364 405748
rect 189420 570332 189476 570388
rect 189308 367052 189364 367108
rect 189196 354956 189252 355012
rect 189084 342860 189140 342916
rect 188860 336140 188916 336196
rect 188076 288428 188132 288484
rect 188748 326732 188804 326788
rect 187964 282156 188020 282212
rect 187516 281372 187572 281428
rect 187180 280476 187236 280532
rect 188188 243516 188244 243572
rect 188076 242060 188132 242116
rect 188188 238476 188244 238532
rect 188076 236236 188132 236292
rect 188748 233100 188804 233156
rect 188860 231196 188916 231252
rect 189196 230972 189252 231028
rect 189084 229740 189140 229796
rect 186396 223132 186452 223188
rect 209580 591276 209636 591332
rect 190652 591164 190708 591220
rect 189644 268940 189700 268996
rect 189756 588812 189812 588868
rect 189532 267596 189588 267652
rect 189420 266252 189476 266308
rect 231644 591164 231700 591220
rect 253708 591052 253764 591108
rect 297836 590940 297892 590996
rect 319900 590828 319956 590884
rect 275772 572012 275828 572068
rect 364028 590716 364084 590772
rect 386316 590716 386372 590772
rect 401436 590716 401492 590772
rect 430220 590604 430276 590660
rect 452508 590604 452564 590660
rect 408268 588812 408324 588868
rect 401436 587916 401492 587972
rect 407372 587916 407428 587972
rect 341964 570332 342020 570388
rect 496412 590492 496468 590548
rect 518476 590156 518532 590212
rect 474348 578732 474404 578788
rect 562604 591276 562660 591332
rect 584668 590156 584724 590212
rect 540540 577052 540596 577108
rect 407372 566972 407428 567028
rect 552748 560364 552804 560420
rect 551068 541548 551124 541604
rect 549948 507836 550004 507892
rect 549500 484428 549556 484484
rect 549388 423388 549444 423444
rect 341404 410396 341460 410452
rect 190652 399084 190708 399140
rect 195132 394156 195188 394212
rect 205884 407596 205940 407652
rect 208348 407932 208404 407988
rect 204764 404012 204820 404068
rect 200508 394044 200564 394100
rect 202860 394716 202916 394772
rect 201964 393148 202020 393204
rect 197372 382172 197428 382228
rect 196476 381948 196532 382004
rect 190652 380604 190708 380660
rect 189756 264908 189812 264964
rect 190092 292572 190148 292628
rect 189308 212604 189364 212660
rect 199164 382172 199220 382228
rect 198044 381948 198100 382004
rect 200844 382172 200900 382228
rect 199724 381948 199780 382004
rect 201404 381948 201460 382004
rect 206556 402444 206612 402500
rect 211036 405804 211092 405860
rect 210140 404124 210196 404180
rect 204316 381948 204372 382004
rect 206108 381948 206164 382004
rect 208236 382172 208292 382228
rect 210364 399756 210420 399812
rect 210364 398188 210420 398244
rect 209916 382172 209972 382228
rect 212828 407484 212884 407540
rect 211260 399756 211316 399812
rect 211932 405692 211988 405748
rect 213724 399084 213780 399140
rect 214508 392364 214564 392420
rect 216300 392252 216356 392308
rect 215404 390684 215460 390740
rect 232764 407372 232820 407428
rect 243516 407932 243572 407988
rect 254268 407932 254324 407988
rect 259644 407596 259700 407652
rect 248892 407484 248948 407540
rect 238140 407036 238196 407092
rect 227612 406588 227668 406644
rect 265020 406588 265076 406644
rect 270396 409052 270452 409108
rect 276332 407708 276388 407764
rect 270396 406588 270452 406644
rect 275548 407484 275604 407540
rect 222012 403228 222068 403284
rect 219996 398972 220052 399028
rect 218204 397292 218260 397348
rect 216636 391356 216692 391412
rect 217196 395612 217252 395668
rect 218988 393932 219044 393988
rect 222012 397404 222068 397460
rect 276332 406588 276388 406644
rect 280028 409052 280084 409108
rect 278236 400652 278292 400708
rect 220780 390796 220836 390852
rect 272188 386764 272244 386820
rect 252028 386540 252084 386596
rect 246764 385308 246820 385364
rect 240716 383628 240772 383684
rect 235116 383180 235172 383236
rect 223468 383068 223524 383124
rect 231644 382284 231700 382340
rect 230076 382172 230132 382228
rect 223692 380268 223748 380324
rect 225484 380156 225540 380212
rect 226828 380044 226884 380100
rect 231756 382172 231812 382228
rect 228956 379932 229012 379988
rect 232204 381948 232260 382004
rect 232652 381836 232708 381892
rect 240156 381836 240212 381892
rect 239484 381388 239540 381444
rect 245196 383628 245252 383684
rect 244972 383068 245028 383124
rect 246652 380156 246708 380212
rect 250572 383964 250628 384020
rect 250348 380716 250404 380772
rect 248556 380044 248612 380100
rect 248668 379932 248724 379988
rect 253708 386428 253764 386484
rect 260540 385532 260596 385588
rect 257068 382060 257124 382116
rect 256060 381612 256116 381668
rect 257740 381724 257796 381780
rect 258748 380604 258804 380660
rect 259532 380492 259588 380548
rect 264124 385420 264180 385476
rect 262108 383740 262164 383796
rect 263788 383404 263844 383460
rect 262332 380380 262388 380436
rect 265468 385196 265524 385252
rect 265916 385084 265972 385140
rect 267708 384972 267764 385028
rect 267260 381500 267316 381556
rect 271292 384860 271348 384916
rect 270732 384748 270788 384804
rect 268828 383516 268884 383572
rect 273084 386652 273140 386708
rect 273868 383292 273924 383348
rect 277228 394492 277284 394548
rect 277116 382060 277172 382116
rect 279020 392252 279076 392308
rect 285516 409164 285572 409220
rect 285516 408156 285572 408212
rect 281372 407820 281428 407876
rect 281372 406588 281428 406644
rect 286412 408044 286468 408100
rect 286412 406588 286468 406644
rect 291452 408156 291508 408212
rect 288988 406140 289044 406196
rect 288204 406028 288260 406084
rect 285404 405916 285460 405972
rect 281820 405804 281876 405860
rect 280924 397292 280980 397348
rect 283612 405692 283668 405748
rect 282604 390684 282660 390740
rect 284508 401324 284564 401380
rect 287980 390796 288036 390852
rect 286972 385532 287028 385588
rect 287196 382060 287252 382116
rect 288204 382060 288260 382116
rect 290668 395612 290724 395668
rect 290556 385644 290612 385700
rect 293468 409948 293524 410004
rect 292572 400764 292628 400820
rect 291676 397404 291732 397460
rect 302652 409724 302708 409780
rect 296492 409276 296548 409332
rect 294364 409164 294420 409220
rect 295260 402780 295316 402836
rect 296156 398972 296212 399028
rect 298844 408604 298900 408660
rect 296492 385756 296548 385812
rect 297052 404572 297108 404628
rect 297948 399084 298004 399140
rect 300636 404460 300692 404516
rect 299740 399196 299796 399252
rect 302428 399532 302484 399588
rect 301532 399308 301588 399364
rect 291452 380492 291508 380548
rect 308028 409836 308084 409892
rect 304220 408492 304276 408548
rect 303324 399420 303380 399476
rect 303212 385868 303268 385924
rect 307804 404236 307860 404292
rect 306012 402668 306068 402724
rect 313404 409388 313460 409444
rect 318332 409500 318388 409556
rect 309596 406364 309652 406420
rect 308252 385980 308308 386036
rect 308700 400876 308756 400932
rect 311388 406252 311444 406308
rect 310492 400988 310548 401044
rect 312284 401212 312340 401268
rect 313068 394604 313124 394660
rect 305676 382060 305732 382116
rect 307356 382060 307412 382116
rect 315756 407596 315812 407652
rect 315756 404348 315812 404404
rect 315868 404124 315924 404180
rect 314076 401100 314132 401156
rect 313292 380604 313348 380660
rect 314860 396284 314916 396340
rect 316652 396172 316708 396228
rect 318780 409500 318836 409556
rect 321244 409276 321300 409332
rect 318332 386092 318388 386148
rect 318444 396060 318500 396116
rect 318332 382060 318388 382116
rect 320236 395948 320292 396004
rect 320124 382060 320180 382116
rect 324156 406588 324212 406644
rect 324828 409500 324884 409556
rect 322028 395836 322084 395892
rect 323820 394380 323876 394436
rect 323596 382060 323652 382116
rect 326620 409388 326676 409444
rect 325612 395724 325668 395780
rect 329420 392588 329476 392644
rect 327404 392364 327460 392420
rect 329196 382060 329252 382116
rect 334908 406588 334964 406644
rect 340172 408268 340228 408324
rect 332892 402892 332948 402948
rect 329532 388108 329588 388164
rect 330988 390908 331044 390964
rect 330876 382060 330932 382116
rect 340060 388780 340116 388836
rect 332556 382172 332612 382228
rect 339500 383628 339556 383684
rect 334236 382060 334292 382116
rect 335468 381500 335524 381556
rect 228060 379820 228116 379876
rect 240604 379820 240660 379876
rect 210364 379708 210420 379764
rect 236124 379708 236180 379764
rect 242396 379708 242452 379764
rect 253148 379484 253204 379540
rect 254940 379484 254996 379540
rect 195468 379372 195524 379428
rect 221788 379372 221844 379428
rect 222684 379372 222740 379428
rect 225372 379372 225428 379428
rect 235228 379372 235284 379428
rect 237020 379372 237076 379428
rect 238476 379372 238532 379428
rect 243292 379372 243348 379428
rect 249900 379372 249956 379428
rect 255836 379372 255892 379428
rect 270172 379372 270228 379428
rect 339388 354508 339444 354564
rect 339276 261436 339332 261492
rect 339276 259980 339332 260036
rect 190652 245420 190708 245476
rect 190652 241052 190708 241108
rect 339276 243516 339332 243572
rect 190540 240380 190596 240436
rect 315644 240604 315700 240660
rect 317884 240604 317940 240660
rect 318556 240604 318612 240660
rect 322588 240604 322644 240660
rect 323260 240604 323316 240660
rect 337148 240604 337204 240660
rect 315644 240380 315700 240436
rect 336028 240268 336084 240324
rect 317212 240156 317268 240212
rect 320572 240156 320628 240212
rect 206332 238476 206388 238532
rect 206332 234332 206388 234388
rect 207676 232652 207732 232708
rect 207004 229404 207060 229460
rect 208348 227612 208404 227668
rect 210364 236124 210420 236180
rect 209692 224364 209748 224420
rect 209020 222796 209076 222852
rect 211036 219212 211092 219268
rect 190092 211260 190148 211316
rect 212380 229516 212436 229572
rect 214396 240044 214452 240100
rect 215068 234556 215124 234612
rect 215740 234444 215796 234500
rect 218428 237020 218484 237076
rect 218316 236908 218372 236964
rect 217084 234556 217140 234612
rect 216412 234444 216468 234500
rect 219772 231644 219828 231700
rect 220444 231532 220500 231588
rect 219100 231420 219156 231476
rect 221116 228060 221172 228116
rect 222460 228172 222516 228228
rect 221788 227612 221844 227668
rect 213724 224476 213780 224532
rect 223804 235004 223860 235060
rect 225148 235116 225204 235172
rect 225820 234220 225876 234276
rect 227836 236460 227892 236516
rect 227164 231756 227220 231812
rect 226492 230860 226548 230916
rect 229180 236908 229236 236964
rect 228508 228284 228564 228340
rect 224476 224924 224532 224980
rect 223132 224364 223188 224420
rect 213052 217532 213108 217588
rect 230524 222684 230580 222740
rect 231196 214396 231252 214452
rect 231868 214284 231924 214340
rect 229852 214172 229908 214228
rect 233212 237244 233268 237300
rect 235900 237244 235956 237300
rect 236796 236908 236852 236964
rect 237244 228396 237300 228452
rect 237916 227500 237972 227556
rect 235228 224252 235284 224308
rect 234556 215964 234612 216020
rect 233884 215852 233940 215908
rect 232540 212492 232596 212548
rect 211708 210812 211764 210868
rect 239260 225036 239316 225092
rect 240604 232652 240660 232708
rect 241948 238476 242004 238532
rect 242620 238476 242676 238532
rect 243292 238364 243348 238420
rect 244636 238252 244692 238308
rect 243964 237804 244020 237860
rect 245980 237916 246036 237972
rect 245308 237692 245364 237748
rect 241276 224252 241332 224308
rect 239932 224140 239988 224196
rect 247324 238476 247380 238532
rect 249340 238140 249396 238196
rect 248668 238028 248724 238084
rect 247996 237468 248052 237524
rect 246652 213276 246708 213332
rect 251356 236348 251412 236404
rect 250684 236124 250740 236180
rect 253372 223244 253428 223300
rect 252700 215964 252756 216020
rect 252028 214172 252084 214228
rect 256060 221340 256116 221396
rect 255388 221228 255444 221284
rect 254716 214956 254772 215012
rect 258076 229404 258132 229460
rect 257404 224476 257460 224532
rect 256732 212492 256788 212548
rect 254044 211596 254100 211652
rect 260092 236572 260148 236628
rect 259420 226492 259476 226548
rect 264796 218204 264852 218260
rect 264124 217532 264180 217588
rect 263452 214844 263508 214900
rect 262780 214396 262836 214452
rect 262108 214284 262164 214340
rect 261436 214060 261492 214116
rect 266140 218316 266196 218372
rect 267484 237020 267540 237076
rect 268604 236908 268660 236964
rect 266812 217420 266868 217476
rect 265468 213052 265524 213108
rect 260764 211484 260820 211540
rect 258748 211372 258804 211428
rect 250012 210700 250068 210756
rect 238588 209916 238644 209972
rect 184604 209468 184660 209524
rect 269500 237020 269556 237076
rect 269724 238252 269780 238308
rect 269276 143612 269332 143668
rect 269388 236460 269444 236516
rect 53228 49532 53284 49588
rect 41132 4508 41188 4564
rect 41804 42812 41860 42868
rect 45612 4956 45668 5012
rect 49420 4284 49476 4340
rect 47516 4172 47572 4228
rect 95116 49532 95172 49588
rect 87500 48188 87556 48244
rect 85708 37884 85764 37940
rect 57148 37772 57204 37828
rect 55132 3388 55188 3444
rect 62748 27692 62804 27748
rect 58940 4060 58996 4116
rect 60844 3388 60900 3444
rect 79884 24556 79940 24612
rect 68460 24444 68516 24500
rect 66556 4844 66612 4900
rect 64652 4396 64708 4452
rect 74172 24332 74228 24388
rect 70364 4620 70420 4676
rect 72268 4508 72324 4564
rect 76076 4956 76132 5012
rect 77980 4732 78036 4788
rect 83692 4284 83748 4340
rect 81788 4172 81844 4228
rect 93212 48076 93268 48132
rect 89404 41132 89460 41188
rect 91532 3388 91588 3444
rect 197932 49756 197988 49812
rect 97356 48636 97412 48692
rect 123676 49644 123732 49700
rect 116060 48076 116116 48132
rect 97356 47852 97412 47908
rect 98924 47964 98980 48020
rect 97020 34412 97076 34468
rect 110348 47964 110404 48020
rect 104636 47852 104692 47908
rect 100828 41244 100884 41300
rect 102732 34524 102788 34580
rect 106540 37996 106596 38052
rect 108444 34636 108500 34692
rect 114380 4620 114436 4676
rect 112476 4172 112532 4228
rect 121772 44492 121828 44548
rect 117964 38108 118020 38164
rect 119868 31052 119924 31108
rect 190316 48412 190372 48468
rect 186508 48300 186564 48356
rect 138908 48188 138964 48244
rect 133196 44716 133252 44772
rect 127484 44604 127540 44660
rect 125580 34748 125636 34804
rect 129388 41356 129444 41412
rect 131292 31164 131348 31220
rect 135100 38332 135156 38388
rect 137004 38220 137060 38276
rect 184604 45276 184660 45332
rect 178892 45164 178948 45220
rect 167468 45052 167524 45108
rect 144620 44940 144676 44996
rect 140812 26012 140868 26068
rect 142940 3388 142996 3444
rect 148428 44828 148484 44884
rect 146748 7532 146804 7588
rect 161756 41692 161812 41748
rect 156044 41580 156100 41636
rect 150332 41468 150388 41524
rect 152236 17612 152292 17668
rect 154364 4284 154420 4340
rect 159852 31276 159908 31332
rect 158172 5852 158228 5908
rect 163660 12572 163716 12628
rect 165788 4396 165844 4452
rect 175084 42924 175140 42980
rect 173180 41804 173236 41860
rect 169372 29372 169428 29428
rect 171500 4060 171556 4116
rect 176988 38444 177044 38500
rect 181020 4844 181076 4900
rect 182924 4508 182980 4564
rect 188412 31388 188468 31444
rect 196028 41020 196084 41076
rect 192220 24668 192276 24724
rect 194348 4732 194404 4788
rect 201740 48524 201796 48580
rect 199948 41916 200004 41972
rect 207452 47740 207508 47796
rect 203644 44380 203700 44436
rect 205772 4956 205828 5012
rect 269612 231756 269668 231812
rect 269388 48524 269444 48580
rect 269500 211260 269556 211316
rect 212268 47628 212324 47684
rect 269500 47628 269556 47684
rect 269612 41020 269668 41076
rect 269836 237468 269892 237524
rect 270396 236908 270452 236964
rect 270732 238476 270788 238532
rect 270620 232652 270676 232708
rect 269836 24668 269892 24724
rect 270508 213276 270564 213332
rect 269724 12572 269780 12628
rect 271068 234444 271124 234500
rect 270844 159292 270900 159348
rect 270956 225036 271012 225092
rect 270732 48300 270788 48356
rect 270620 41356 270676 41412
rect 271068 47852 271124 47908
rect 271180 231420 271236 231476
rect 271292 228284 271348 228340
rect 272412 211260 272468 211316
rect 272188 210812 272244 210868
rect 272300 210924 272356 210980
rect 271516 152236 271572 152292
rect 272188 209916 272244 209972
rect 271292 47740 271348 47796
rect 271180 44604 271236 44660
rect 270956 38108 271012 38164
rect 270508 4844 270564 4900
rect 211484 4620 211540 4676
rect 209580 4060 209636 4116
rect 272860 210924 272916 210980
rect 272972 231420 273028 231476
rect 272636 209916 272692 209972
rect 272524 209132 272580 209188
rect 272748 209804 272804 209860
rect 272748 180796 272804 180852
rect 272636 177884 272692 177940
rect 272524 174972 272580 175028
rect 272412 172060 272468 172116
rect 272300 160412 272356 160468
rect 272524 153580 272580 153636
rect 272300 145292 272356 145348
rect 272412 142940 272468 142996
rect 272524 131292 272580 131348
rect 273868 238140 273924 238196
rect 273532 211036 273588 211092
rect 273756 236012 273812 236068
rect 273756 235116 273812 235172
rect 273084 205884 273140 205940
rect 273420 154476 273476 154532
rect 273196 154252 273252 154308
rect 273196 134204 273252 134260
rect 273308 145404 273364 145460
rect 273756 153580 273812 153636
rect 273532 143724 273588 143780
rect 273532 142940 273588 142996
rect 273420 137116 273476 137172
rect 273308 128380 273364 128436
rect 273756 126812 273812 126868
rect 273756 125468 273812 125524
rect 273084 102172 273140 102228
rect 272972 99260 273028 99316
rect 273308 101612 273364 101668
rect 273308 73052 273364 73108
rect 273084 70140 273140 70196
rect 272972 67228 273028 67284
rect 273084 52780 273140 52836
rect 273196 61404 273252 61460
rect 272972 50540 273028 50596
rect 272412 50316 272468 50372
rect 273196 49644 273252 49700
rect 273980 238028 274036 238084
rect 273980 49756 274036 49812
rect 274092 228172 274148 228228
rect 273868 44380 273924 44436
rect 274428 231532 274484 231588
rect 274204 160300 274260 160356
rect 274316 224924 274372 224980
rect 274428 48188 274484 48244
rect 274540 228060 274596 228116
rect 274652 210028 274708 210084
rect 274876 160636 274932 160692
rect 275772 227612 275828 227668
rect 275548 160524 275604 160580
rect 275660 224252 275716 224308
rect 274652 154364 274708 154420
rect 274652 141932 274708 141988
rect 274652 81788 274708 81844
rect 275436 58492 275492 58548
rect 275548 52668 275604 52724
rect 275548 50652 275604 50708
rect 275436 49756 275492 49812
rect 274540 44940 274596 44996
rect 274316 41804 274372 41860
rect 274092 41580 274148 41636
rect 275884 224364 275940 224420
rect 276220 197148 276276 197204
rect 276332 224364 276388 224420
rect 275884 41692 275940 41748
rect 275772 41468 275828 41524
rect 275660 38332 275716 38388
rect 272300 36764 272356 36820
rect 276444 219212 276500 219268
rect 276892 150892 276948 150948
rect 277228 237804 277284 237860
rect 276556 138572 276612 138628
rect 276556 75964 276612 76020
rect 276556 64316 276612 64372
rect 276556 49532 276612 49588
rect 276444 38444 276500 38500
rect 276332 24444 276388 24500
rect 278908 238140 278964 238196
rect 278236 238028 278292 238084
rect 277564 237804 277620 237860
rect 279020 237916 279076 237972
rect 278908 237692 278964 237748
rect 278124 224252 278180 224308
rect 278012 219660 278068 219716
rect 277228 5852 277284 5908
rect 277340 210700 277396 210756
rect 272188 4172 272244 4228
rect 278236 131964 278292 132020
rect 278236 78876 278292 78932
rect 278124 41916 278180 41972
rect 278012 31388 278068 31444
rect 279580 237692 279636 237748
rect 279020 42924 279076 42980
rect 279692 236236 279748 236292
rect 279692 33628 279748 33684
rect 279804 227612 279860 227668
rect 279916 222796 279972 222852
rect 280028 219772 280084 219828
rect 280924 238252 280980 238308
rect 280252 155932 280308 155988
rect 280364 219884 280420 219940
rect 282268 237916 282324 237972
rect 283164 226156 283220 226212
rect 282940 155484 282996 155540
rect 283052 222684 283108 222740
rect 281596 152796 281652 152852
rect 280364 44828 280420 44884
rect 280028 42812 280084 42868
rect 279916 38220 279972 38276
rect 279804 31276 279860 31332
rect 283612 152124 283668 152180
rect 284956 151004 285012 151060
rect 284284 150780 284340 150836
rect 286300 238476 286356 238532
rect 286636 226268 286692 226324
rect 285628 149100 285684 149156
rect 286412 226044 286468 226100
rect 283164 34748 283220 34804
rect 286412 34636 286468 34692
rect 286860 225932 286916 225988
rect 286972 159404 287028 159460
rect 287644 159068 287700 159124
rect 288204 239260 288260 239316
rect 286860 34524 286916 34580
rect 286636 34412 286692 34468
rect 283052 31164 283108 31220
rect 278908 29372 278964 29428
rect 288988 238364 289044 238420
rect 289660 158956 289716 159012
rect 289772 234332 289828 234388
rect 288316 158844 288372 158900
rect 288988 55580 289044 55636
rect 288988 50428 289044 50484
rect 288204 4956 288260 5012
rect 289884 226380 289940 226436
rect 289884 31052 289940 31108
rect 289996 216412 290052 216468
rect 290220 216300 290276 216356
rect 290332 161868 290388 161924
rect 291004 150668 291060 150724
rect 292348 237020 292404 237076
rect 293244 238252 293300 238308
rect 293020 162092 293076 162148
rect 293132 211596 293188 211652
rect 291676 150332 291732 150388
rect 293804 236908 293860 236964
rect 293244 152348 293300 152404
rect 294812 238476 294868 238532
rect 295596 236908 295652 236964
rect 294812 155596 294868 155652
rect 294364 152012 294420 152068
rect 295708 149436 295764 149492
rect 296380 149212 296436 149268
rect 296492 214956 296548 215012
rect 297724 236908 297780 236964
rect 297052 155372 297108 155428
rect 298172 236348 298228 236404
rect 298396 161980 298452 162036
rect 299740 236908 299796 236964
rect 299964 238364 300020 238420
rect 299068 148652 299124 148708
rect 299852 212492 299908 212548
rect 298172 123900 298228 123956
rect 296492 123676 296548 123732
rect 293132 123564 293188 123620
rect 299964 159180 300020 159236
rect 301644 238140 301700 238196
rect 301084 160412 301140 160468
rect 301532 236124 301588 236180
rect 300412 158732 300468 158788
rect 301756 233436 301812 233492
rect 303100 240044 303156 240100
rect 302428 228396 302484 228452
rect 303548 237916 303604 237972
rect 303436 221340 303492 221396
rect 303212 221228 303268 221284
rect 301644 155708 301700 155764
rect 303100 213052 303156 213108
rect 303100 133756 303156 133812
rect 303212 127372 303268 127428
rect 303324 215964 303380 216020
rect 301532 124236 301588 124292
rect 303772 236236 303828 236292
rect 303996 238028 304052 238084
rect 303548 149548 303604 149604
rect 303660 218316 303716 218372
rect 303660 133644 303716 133700
rect 303884 217420 303940 217476
rect 304444 236460 304500 236516
rect 304892 239372 304948 239428
rect 303996 155820 304052 155876
rect 305004 237804 305060 237860
rect 305116 236684 305172 236740
rect 306460 237580 306516 237636
rect 305788 236348 305844 236404
rect 307132 236124 307188 236180
rect 307356 239260 307412 239316
rect 307356 236572 307412 236628
rect 307356 236012 307412 236068
rect 308476 237468 308532 237524
rect 308700 237692 308756 237748
rect 307804 236012 307860 236068
rect 305116 231308 305172 231364
rect 305116 204092 305172 204148
rect 306572 223244 306628 223300
rect 305004 156156 305060 156212
rect 304892 152460 304948 152516
rect 303884 133532 303940 133588
rect 303436 130396 303492 130452
rect 307020 218204 307076 218260
rect 306796 217532 306852 217588
rect 306684 214396 306740 214452
rect 306796 130172 306852 130228
rect 306908 214284 306964 214340
rect 307020 133868 307076 133924
rect 307132 214844 307188 214900
rect 308252 214172 308308 214228
rect 307132 130284 307188 130340
rect 307244 211484 307300 211540
rect 307244 127260 307300 127316
rect 306908 127148 306964 127204
rect 306684 127036 306740 127092
rect 306572 124124 306628 124180
rect 303324 124012 303380 124068
rect 299852 123452 299908 123508
rect 311164 238140 311220 238196
rect 313180 238364 313236 238420
rect 312508 238252 312564 238308
rect 311836 237804 311892 237860
rect 310492 237692 310548 237748
rect 312508 237468 312564 237524
rect 314524 237916 314580 237972
rect 313852 237468 313908 237524
rect 312508 235004 312564 235060
rect 315868 238028 315924 238084
rect 316540 236796 316596 236852
rect 318332 239484 318388 239540
rect 315196 234892 315252 234948
rect 311164 234556 311220 234612
rect 309820 230860 309876 230916
rect 309932 232652 309988 232708
rect 309148 230076 309204 230132
rect 308700 156044 308756 156100
rect 308252 123340 308308 123396
rect 311052 230188 311108 230244
rect 310156 229404 310212 229460
rect 310044 224476 310100 224532
rect 310044 123788 310100 123844
rect 310268 219548 310324 219604
rect 310940 214620 310996 214676
rect 310380 211036 310436 211092
rect 310380 160188 310436 160244
rect 310604 210924 310660 210980
rect 310604 159852 310660 159908
rect 310268 157612 310324 157668
rect 310156 119644 310212 119700
rect 309932 116732 309988 116788
rect 311052 105084 311108 105140
rect 311612 233100 311668 233156
rect 314972 229852 315028 229908
rect 312732 217868 312788 217924
rect 313852 217756 313908 217812
rect 317212 221004 317268 221060
rect 316092 219436 316148 219492
rect 319900 240044 319956 240100
rect 319228 239484 319284 239540
rect 321244 238476 321300 238532
rect 325836 240044 325892 240100
rect 325836 239372 325892 239428
rect 321916 238476 321972 238532
rect 330652 234780 330708 234836
rect 321692 234108 321748 234164
rect 320572 232988 320628 233044
rect 319452 231196 319508 231252
rect 326172 232876 326228 232932
rect 325052 229740 325108 229796
rect 322812 227948 322868 228004
rect 321804 224700 321860 224756
rect 321804 214172 321860 214228
rect 323932 217644 323988 217700
rect 328412 231084 328468 231140
rect 327292 224812 327348 224868
rect 329532 227836 329588 227892
rect 336028 231084 336084 231140
rect 336252 232764 336308 232820
rect 335132 230972 335188 231028
rect 332892 229628 332948 229684
rect 331772 223020 331828 223076
rect 331996 222908 332052 222964
rect 331996 209132 332052 209188
rect 334012 219324 334068 219380
rect 337148 219884 337204 219940
rect 337372 224588 337428 224644
rect 338492 223132 338548 223188
rect 339276 216412 339332 216468
rect 339388 198156 339444 198212
rect 339612 381388 339668 381444
rect 339948 281148 340004 281204
rect 339948 280588 340004 280644
rect 339612 239372 339668 239428
rect 341292 409612 341348 409668
rect 340284 360444 340340 360500
rect 340284 359548 340340 359604
rect 340396 396732 340452 396788
rect 340172 237468 340228 237524
rect 340060 236796 340116 236852
rect 340732 389340 340788 389396
rect 340396 236012 340452 236068
rect 340508 389116 340564 389172
rect 340956 389228 341012 389284
rect 341180 381836 341236 381892
rect 341068 252140 341124 252196
rect 341068 243516 341124 243572
rect 345324 394828 345380 394884
rect 343756 393372 343812 393428
rect 343532 393260 343588 393316
rect 341852 392700 341908 392756
rect 341628 381500 341684 381556
rect 341404 294812 341460 294868
rect 341404 294252 341460 294308
rect 341516 380156 341572 380212
rect 341292 291564 341348 291620
rect 341292 282604 341348 282660
rect 341292 240604 341348 240660
rect 341404 261100 341460 261156
rect 341180 239036 341236 239092
rect 340956 235004 341012 235060
rect 340732 234892 340788 234948
rect 340508 230076 340564 230132
rect 340732 227724 340788 227780
rect 339500 197820 339556 197876
rect 339612 220892 339668 220948
rect 341404 222684 341460 222740
rect 341516 197708 341572 197764
rect 341740 234668 341796 234724
rect 342972 390572 343028 390628
rect 341852 233436 341908 233492
rect 341964 389452 342020 389508
rect 342860 388892 342916 388948
rect 342076 385868 342132 385924
rect 342076 319788 342132 319844
rect 342972 295148 343028 295204
rect 343084 387212 343140 387268
rect 343756 373996 343812 374052
rect 345212 385308 345268 385364
rect 343532 371308 343588 371364
rect 344764 364140 344820 364196
rect 343532 345324 343588 345380
rect 343084 293132 343140 293188
rect 343196 340844 343252 340900
rect 342748 292460 342804 292516
rect 342076 290668 342132 290724
rect 342860 273644 342916 273700
rect 342748 262892 342804 262948
rect 342748 241612 342804 241668
rect 342076 234556 342132 234612
rect 342188 240716 342244 240772
rect 341964 230860 342020 230916
rect 342972 272748 343028 272804
rect 342972 241164 343028 241220
rect 343084 266476 343140 266532
rect 343084 240940 343140 240996
rect 342860 234332 342916 234388
rect 342188 219212 342244 219268
rect 342972 201516 343028 201572
rect 341628 196476 341684 196532
rect 343308 264684 343364 264740
rect 344092 339052 344148 339108
rect 343532 251132 343588 251188
rect 343644 338156 343700 338212
rect 343308 241836 343364 241892
rect 343420 249452 343476 249508
rect 343420 231196 343476 231252
rect 343532 240380 343588 240436
rect 343532 215852 343588 215908
rect 343756 240828 343812 240884
rect 343756 224252 343812 224308
rect 343980 209468 344036 209524
rect 344316 278796 344372 278852
rect 344316 264572 344372 264628
rect 343196 196364 343252 196420
rect 344316 196364 344372 196420
rect 345100 252028 345156 252084
rect 345100 240268 345156 240324
rect 345100 212604 345156 212660
rect 345548 386092 345604 386148
rect 345324 237804 345380 237860
rect 345436 358764 345492 358820
rect 350476 403340 350532 403396
rect 347228 396844 347284 396900
rect 345660 367052 345716 367108
rect 346444 379708 346500 379764
rect 345548 336028 345604 336084
rect 345548 229404 345604 229460
rect 345660 342636 345716 342692
rect 345212 198044 345268 198100
rect 345548 196588 345604 196644
rect 344988 196530 345044 196532
rect 344988 196478 344990 196530
rect 344990 196478 345042 196530
rect 345042 196478 345044 196530
rect 344988 196476 345044 196478
rect 344764 196364 344820 196420
rect 345996 272076 346052 272132
rect 345772 252476 345828 252532
rect 345660 196364 345716 196420
rect 346108 263788 346164 263844
rect 346108 240492 346164 240548
rect 346220 253036 346276 253092
rect 346220 240380 346276 240436
rect 345996 198156 346052 198212
rect 345884 196364 345940 196420
rect 313404 160636 313460 160692
rect 314972 160076 315028 160132
rect 317436 160076 317492 160132
rect 319676 157612 319732 157668
rect 321244 157612 321300 157668
rect 318108 156940 318164 156996
rect 324380 157836 324436 157892
rect 329084 160076 329140 160132
rect 330652 157836 330708 157892
rect 332220 157836 332276 157892
rect 327516 157724 327572 157780
rect 325948 157500 326004 157556
rect 335356 157836 335412 157892
rect 340060 159516 340116 159572
rect 338492 158620 338548 158676
rect 344764 160076 344820 160132
rect 343196 159740 343252 159796
rect 341628 157724 341684 157780
rect 346108 157836 346164 157892
rect 336924 157500 336980 157556
rect 346892 369516 346948 369572
rect 346556 196364 346612 196420
rect 346444 157612 346500 157668
rect 346108 157388 346164 157444
rect 347004 361452 347060 361508
rect 347116 351596 347172 351652
rect 348572 370412 348628 370468
rect 347788 309484 347844 309540
rect 347676 296492 347732 296548
rect 347228 236124 347284 236180
rect 347564 284732 347620 284788
rect 347116 172396 347172 172452
rect 347004 171052 347060 171108
rect 347004 167804 347060 167860
rect 346780 157388 346836 157444
rect 333788 157276 333844 157332
rect 322812 156828 322868 156884
rect 345212 153804 345268 153860
rect 341852 146972 341908 147028
rect 345324 151788 345380 151844
rect 345324 140028 345380 140084
rect 345212 126812 345268 126868
rect 341852 122556 341908 122612
rect 311164 96348 311220 96404
rect 307468 50316 307524 50372
rect 315308 50316 315364 50372
rect 293580 48636 293636 48692
rect 290220 48524 290276 48580
rect 300748 48524 300804 48580
rect 322252 48524 322308 48580
rect 347788 238588 347844 238644
rect 347900 198044 347956 198100
rect 347788 196476 347844 196532
rect 350252 365036 350308 365092
rect 348572 171276 348628 171332
rect 348684 362348 348740 362404
rect 348796 354284 348852 354340
rect 348796 172620 348852 172676
rect 348908 352492 348964 352548
rect 348684 169372 348740 169428
rect 349020 349804 349076 349860
rect 349132 283836 349188 283892
rect 349356 283724 349412 283780
rect 349132 241948 349188 242004
rect 349244 248556 349300 248612
rect 349020 174188 349076 174244
rect 348908 168700 348964 168756
rect 347900 159964 347956 160020
rect 347788 157500 347844 157556
rect 349244 150556 349300 150612
rect 349580 271852 349636 271908
rect 349468 257516 349524 257572
rect 349580 240828 349636 240884
rect 349468 226044 349524 226100
rect 349580 196252 349636 196308
rect 350364 356076 350420 356132
rect 350700 394044 350756 394100
rect 350476 237916 350532 237972
rect 350588 296492 350644 296548
rect 350364 172732 350420 172788
rect 350476 189756 350532 189812
rect 350252 169484 350308 169540
rect 349580 160076 349636 160132
rect 350476 153020 350532 153076
rect 349356 148876 349412 148932
rect 350924 392476 350980 392532
rect 350700 238140 350756 238196
rect 350812 305676 350868 305732
rect 350700 197372 350756 197428
rect 353612 408044 353668 408100
rect 351932 407820 351988 407876
rect 352156 407708 352212 407764
rect 352156 397404 352212 397460
rect 352268 401772 352324 401828
rect 351932 385644 351988 385700
rect 351036 372204 351092 372260
rect 351148 379820 351204 379876
rect 350924 237580 350980 237636
rect 351036 209916 351092 209972
rect 350812 189756 350868 189812
rect 350924 193228 350980 193284
rect 350700 164220 350756 164276
rect 350812 188076 350868 188132
rect 350812 186508 350868 186564
rect 350588 162316 350644 162372
rect 350700 160076 350756 160132
rect 350700 157164 350756 157220
rect 350588 153468 350644 153524
rect 350700 145292 350756 145348
rect 350252 143724 350308 143780
rect 350252 119308 350308 119364
rect 350252 101612 350308 101668
rect 347676 50316 347732 50372
rect 347564 48524 347620 48580
rect 351932 367724 351988 367780
rect 351260 313292 351316 313348
rect 351372 268268 351428 268324
rect 351372 240716 351428 240772
rect 351260 231308 351316 231364
rect 351820 236796 351876 236852
rect 351260 197260 351316 197316
rect 351820 188076 351876 188132
rect 352044 359660 352100 359716
rect 352156 348908 352212 348964
rect 352268 238028 352324 238084
rect 352380 397404 352436 397460
rect 355404 407260 355460 407316
rect 355180 407148 355236 407204
rect 353612 385532 353668 385588
rect 354172 405020 354228 405076
rect 352604 383068 352660 383124
rect 352380 236236 352436 236292
rect 352492 380604 352548 380660
rect 352492 330988 352548 331044
rect 352604 305676 352660 305732
rect 352828 379372 352884 379428
rect 352492 232652 352548 232708
rect 352156 173628 352212 173684
rect 352268 197148 352324 197204
rect 352044 170940 352100 170996
rect 351932 169596 351988 169652
rect 352716 191660 352772 191716
rect 352268 164108 352324 164164
rect 352604 191548 352660 191604
rect 352492 159516 352548 159572
rect 352492 157612 352548 157668
rect 351484 157276 351540 157332
rect 351148 156940 351204 156996
rect 352604 120204 352660 120260
rect 351036 50204 351092 50260
rect 350924 48412 350980 48468
rect 353612 365932 353668 365988
rect 352828 156828 352884 156884
rect 352940 247772 352996 247828
rect 353724 356972 353780 357028
rect 354060 346220 354116 346276
rect 353724 170828 353780 170884
rect 353836 294812 353892 294868
rect 353612 167580 353668 167636
rect 352940 151116 352996 151172
rect 353836 121996 353892 122052
rect 353948 291452 354004 291508
rect 355180 397292 355236 397348
rect 355292 402556 355348 402612
rect 355404 390684 355460 390740
rect 355516 396956 355572 397012
rect 355292 382172 355348 382228
rect 355292 366828 355348 366884
rect 354172 238252 354228 238308
rect 354396 282156 354452 282212
rect 354060 175196 354116 175252
rect 354172 195916 354228 195972
rect 354172 174300 354228 174356
rect 353948 120316 354004 120372
rect 352716 48300 352772 48356
rect 354620 265580 354676 265636
rect 354620 227612 354676 227668
rect 354508 195804 354564 195860
rect 355404 357868 355460 357924
rect 355740 389564 355796 389620
rect 355516 236348 355572 236404
rect 355628 348012 355684 348068
rect 355404 172844 355460 172900
rect 355516 210812 355572 210868
rect 359884 407932 359940 407988
rect 358764 407596 358820 407652
rect 357196 407372 357252 407428
rect 357084 394940 357140 394996
rect 356412 378028 356468 378084
rect 356748 394156 356804 394212
rect 355740 296492 355796 296548
rect 355964 280476 356020 280532
rect 355852 204988 355908 205044
rect 355852 172956 355908 173012
rect 355628 172284 355684 172340
rect 355516 169036 355572 169092
rect 355292 167692 355348 167748
rect 354508 157724 354564 157780
rect 355964 122108 356020 122164
rect 356076 280364 356132 280420
rect 356188 251132 356244 251188
rect 356636 245196 356692 245252
rect 356636 244076 356692 244132
rect 356972 372204 357028 372260
rect 356748 238364 356804 238420
rect 356860 284844 356916 284900
rect 356636 236796 356692 236852
rect 356188 204988 356244 205044
rect 356748 204092 356804 204148
rect 356748 203308 356804 203364
rect 356188 196028 356244 196084
rect 356188 185836 356244 185892
rect 356748 167356 356804 167412
rect 356860 166236 356916 166292
rect 357756 406700 357812 406756
rect 357420 406588 357476 406644
rect 357196 245196 357252 245252
rect 357308 397180 357364 397236
rect 357644 406588 357700 406644
rect 357532 399644 357588 399700
rect 357532 389564 357588 389620
rect 357644 383740 357700 383796
rect 357644 383068 357700 383124
rect 357420 249788 357476 249844
rect 357644 378028 357700 378084
rect 357308 236460 357364 236516
rect 357084 228396 357140 228452
rect 357196 232316 357252 232372
rect 356972 154364 357028 154420
rect 357084 226492 357140 226548
rect 357196 181132 357252 181188
rect 357308 214844 357364 214900
rect 357084 178444 357140 178500
rect 356188 153356 356244 153412
rect 357308 173068 357364 173124
rect 357420 209132 357476 209188
rect 357420 170380 357476 170436
rect 357084 151900 357140 151956
rect 357532 166236 357588 166292
rect 357532 164668 357588 164724
rect 356188 151788 356244 151844
rect 356972 108220 357028 108276
rect 358652 397068 358708 397124
rect 357868 296380 357924 296436
rect 357868 295708 357924 295764
rect 357756 268716 357812 268772
rect 358428 240268 358484 240324
rect 357868 195692 357924 195748
rect 357644 153356 357700 153412
rect 357756 179900 357812 179956
rect 357532 108220 357588 108276
rect 356972 93436 357028 93492
rect 359548 398300 359604 398356
rect 359212 397516 359268 397572
rect 358764 390796 358820 390852
rect 358988 397292 359044 397348
rect 358876 290668 358932 290724
rect 358764 278908 358820 278964
rect 358764 272972 358820 273028
rect 358652 236684 358708 236740
rect 358764 249452 358820 249508
rect 358764 239932 358820 239988
rect 358428 174636 358484 174692
rect 358540 235116 358596 235172
rect 358540 165676 358596 165732
rect 358652 183820 358708 183876
rect 358988 240044 359044 240100
rect 359100 302092 359156 302148
rect 361788 406588 361844 406644
rect 372540 407484 372596 407540
rect 367164 399644 367220 399700
rect 375228 397292 375284 397348
rect 362908 395052 362964 395108
rect 369180 394940 369236 394996
rect 383292 407932 383348 407988
rect 391356 408604 391412 408660
rect 391356 408156 391412 408212
rect 388668 407148 388724 407204
rect 393148 407484 393204 407540
rect 394044 407260 394100 407316
rect 393148 402892 393204 402948
rect 404796 408044 404852 408100
rect 405692 409948 405748 410004
rect 405692 407932 405748 407988
rect 417452 408492 417508 408548
rect 417452 408044 417508 408100
rect 415548 407820 415604 407876
rect 426300 407932 426356 407988
rect 429660 410060 429716 410116
rect 420924 407820 420980 407876
rect 421596 407708 421652 407764
rect 410172 407596 410228 407652
rect 412412 407596 412468 407652
rect 399420 401324 399476 401380
rect 381276 397404 381332 397460
rect 387324 397180 387380 397236
rect 393372 397068 393428 397124
rect 399420 396956 399476 397012
rect 411516 396844 411572 396900
rect 421596 406364 421652 406420
rect 423612 398300 423668 398356
rect 417564 396732 417620 396788
rect 442428 408156 442484 408212
rect 441868 407820 441924 407876
rect 441868 406252 441924 406308
rect 437052 404572 437108 404628
rect 447804 404460 447860 404516
rect 431676 402780 431732 402836
rect 435708 403452 435764 403508
rect 458556 408044 458612 408100
rect 453628 407932 453684 407988
rect 463932 407932 463988 407988
rect 453628 402668 453684 402724
rect 459900 405020 459956 405076
rect 453180 399532 453236 399588
rect 469308 404236 469364 404292
rect 471996 408268 472052 408324
rect 471884 399980 471940 400036
rect 471884 397404 471940 397460
rect 480060 407820 480116 407876
rect 484092 408380 484148 408436
rect 474684 407708 474740 407764
rect 479612 407708 479668 407764
rect 478044 403340 478100 403396
rect 479612 396284 479668 396340
rect 490812 407708 490868 407764
rect 485436 407596 485492 407652
rect 486332 407596 486388 407652
rect 453852 394828 453908 394884
rect 412412 394604 412468 394660
rect 377916 394492 377972 394548
rect 405468 394492 405524 394548
rect 441756 394492 441812 394548
rect 491372 406588 491428 406644
rect 490140 401772 490196 401828
rect 496188 406588 496244 406644
rect 491372 396172 491428 396228
rect 496188 399868 496244 399924
rect 501564 396060 501620 396116
rect 502236 404908 502292 404964
rect 506940 395948 506996 396004
rect 508284 396620 508340 396676
rect 517692 407596 517748 407652
rect 520380 398076 520436 398132
rect 512316 395836 512372 395892
rect 514332 397516 514388 397572
rect 533820 407596 533876 407652
rect 539196 407596 539252 407652
rect 549388 409052 549444 409108
rect 544572 407484 544628 407540
rect 528444 407372 528500 407428
rect 544572 401660 544628 401716
rect 523068 395724 523124 395780
rect 526428 396844 526484 396900
rect 532476 396732 532532 396788
rect 549500 399420 549556 399476
rect 549612 475468 549668 475524
rect 549612 399196 549668 399252
rect 549724 465724 549780 465780
rect 549836 428428 549892 428484
rect 549836 405804 549892 405860
rect 551068 409500 551124 409556
rect 551180 532140 551236 532196
rect 551180 409276 551236 409332
rect 551292 513324 551348 513380
rect 549948 401212 550004 401268
rect 551292 401100 551348 401156
rect 551404 480396 551460 480452
rect 551404 399308 551460 399364
rect 551516 470988 551572 471044
rect 551628 419244 551684 419300
rect 554428 546252 554484 546308
rect 552748 402556 552804 402612
rect 552860 452172 552916 452228
rect 551628 400652 551684 400708
rect 551516 399084 551572 399140
rect 549724 398972 549780 399028
rect 550620 396508 550676 396564
rect 552972 447468 553028 447524
rect 552972 406140 553028 406196
rect 553084 442764 553140 442820
rect 553084 406028 553140 406084
rect 553196 438060 553252 438116
rect 553196 405916 553252 405972
rect 553308 433356 553364 433412
rect 554428 409388 554484 409444
rect 554540 518028 554596 518084
rect 553308 405692 553364 405748
rect 554540 404124 554596 404180
rect 554652 503916 554708 503972
rect 554652 400988 554708 401044
rect 554764 499212 554820 499268
rect 563612 496076 563668 496132
rect 554988 461580 555044 461636
rect 554764 400876 554820 400932
rect 554876 456876 554932 456932
rect 554988 409164 555044 409220
rect 554876 400764 554932 400820
rect 558908 407372 558964 407428
rect 552860 395612 552916 395668
rect 556668 396620 556724 396676
rect 538524 394828 538580 394884
rect 486332 394380 486388 394436
rect 447804 394268 447860 394324
rect 465948 394268 466004 394324
rect 359884 392252 359940 392308
rect 359884 389900 359940 389956
rect 359884 389340 359940 389396
rect 359548 389228 359604 389284
rect 359772 354676 359828 354732
rect 359436 337148 359492 337204
rect 359436 336028 359492 336084
rect 359212 241276 359268 241332
rect 359324 296380 359380 296436
rect 359100 174076 359156 174132
rect 358876 170604 358932 170660
rect 358764 169148 358820 169204
rect 358652 162876 358708 162932
rect 359884 236572 359940 236628
rect 359884 209244 359940 209300
rect 359884 205772 359940 205828
rect 359436 173852 359492 173908
rect 359884 198044 359940 198100
rect 359884 172508 359940 172564
rect 361228 175308 361284 175364
rect 369180 175196 369236 175252
rect 375228 175196 375284 175252
rect 361228 167468 361284 167524
rect 361340 173068 361396 173124
rect 363132 172956 363188 173012
rect 399420 175084 399476 175140
rect 393372 174188 393428 174244
rect 387324 173628 387380 173684
rect 405468 172396 405524 172452
rect 381276 172284 381332 172340
rect 417564 174636 417620 174692
rect 423612 172620 423668 172676
rect 435708 172732 435764 172788
rect 429660 172508 429716 172564
rect 453852 174300 453908 174356
rect 447804 172844 447860 172900
rect 465948 174412 466004 174468
rect 459900 170940 459956 170996
rect 469532 172284 469588 172340
rect 441756 170828 441812 170884
rect 411516 168700 411572 168756
rect 420812 170380 420868 170436
rect 361340 165788 361396 165844
rect 359324 162316 359380 162372
rect 357868 158620 357924 158676
rect 357868 157836 357924 157892
rect 467852 169260 467908 169316
rect 423164 167468 423220 167524
rect 420924 167356 420980 167412
rect 422940 165788 422996 165844
rect 421596 163212 421652 163268
rect 421596 162876 421652 162932
rect 420924 156380 420980 156436
rect 421708 162540 421764 162596
rect 421708 156268 421764 156324
rect 420812 154924 420868 154980
rect 421708 151900 421764 151956
rect 417116 143612 417172 143668
rect 405020 133868 405076 133924
rect 378812 130396 378868 130452
rect 376796 127372 376852 127428
rect 362684 124236 362740 124292
rect 370748 124124 370804 124180
rect 368732 124012 368788 124068
rect 364700 123900 364756 123956
rect 366716 123340 366772 123396
rect 374780 123676 374836 123732
rect 372764 123564 372820 123620
rect 400988 130284 401044 130340
rect 392924 127260 392980 127316
rect 382844 123788 382900 123844
rect 380828 123452 380884 123508
rect 384860 122668 384916 122724
rect 386876 122668 386932 122724
rect 388892 122668 388948 122724
rect 390908 122668 390964 122724
rect 396956 127148 397012 127204
rect 394940 122668 394996 122724
rect 398972 127036 399028 127092
rect 403004 130172 403060 130228
rect 407036 133756 407092 133812
rect 409052 133644 409108 133700
rect 411068 133532 411124 133588
rect 413084 122668 413140 122724
rect 414988 122668 415044 122724
rect 420140 95228 420196 95284
rect 357756 61628 357812 61684
rect 356076 49868 356132 49924
rect 356188 51884 356244 51940
rect 357756 51884 357812 51940
rect 419244 53004 419300 53060
rect 420028 52780 420084 52836
rect 420140 88284 420196 88340
rect 419244 50652 419300 50708
rect 422492 156380 422548 156436
rect 422492 154140 422548 154196
rect 421932 119308 421988 119364
rect 421932 102396 421988 102452
rect 421820 95228 421876 95284
rect 421708 81340 421764 81396
rect 420140 50540 420196 50596
rect 420252 74396 420308 74452
rect 421820 68796 421876 68852
rect 421820 67452 421876 67508
rect 421932 60508 421988 60564
rect 421932 50428 421988 50484
rect 421820 49756 421876 49812
rect 420252 49644 420308 49700
rect 422604 156268 422660 156324
rect 422604 88284 422660 88340
rect 422716 154924 422772 154980
rect 422716 154028 422772 154084
rect 422940 153916 422996 153972
rect 423164 153804 423220 153860
rect 466284 162428 466340 162484
rect 466284 154140 466340 154196
rect 423276 153244 423332 153300
rect 423276 151900 423332 151956
rect 459452 151228 459508 151284
rect 457996 122108 458052 122164
rect 457884 120316 457940 120372
rect 457772 116956 457828 117012
rect 458220 121996 458276 122052
rect 458108 120204 458164 120260
rect 458108 113036 458164 113092
rect 458220 110124 458276 110180
rect 458556 117516 458612 117572
rect 457996 107212 458052 107268
rect 458556 104300 458612 104356
rect 467852 154028 467908 154084
rect 468972 164332 469028 164388
rect 468972 153916 469028 153972
rect 471996 171052 472052 171108
rect 484092 171164 484148 171220
rect 489132 174076 489188 174132
rect 478044 169372 478100 169428
rect 486444 170604 486500 170660
rect 483756 169148 483812 169204
rect 482412 165676 482468 165732
rect 477036 164892 477092 164948
rect 474348 163212 474404 163268
rect 473004 156268 473060 156324
rect 473004 154476 473060 154532
rect 469532 153804 469588 153860
rect 471660 153804 471716 153860
rect 471660 153244 471716 153300
rect 474348 154364 474404 154420
rect 475692 151228 475748 151284
rect 478380 164780 478436 164836
rect 479724 163100 479780 163156
rect 485100 164668 485156 164724
rect 487788 162316 487844 162372
rect 490140 172060 490196 172116
rect 495852 173964 495908 174020
rect 494508 170492 494564 170548
rect 491820 154252 491876 154308
rect 490476 154028 490532 154084
rect 493164 153244 493220 153300
rect 496188 169484 496244 169540
rect 497196 173852 497252 173908
rect 520380 174524 520436 174580
rect 514332 169596 514388 169652
rect 508284 167692 508340 167748
rect 516012 169036 516068 169092
rect 502236 167580 502292 167636
rect 498540 166348 498596 166404
rect 510636 164220 510692 164276
rect 499884 162988 499940 163044
rect 503916 155932 503972 155988
rect 503916 153916 503972 153972
rect 505260 153692 505316 153748
rect 503916 153244 503972 153300
rect 502572 152908 502628 152964
rect 503132 152908 503188 152964
rect 481068 149772 481124 149828
rect 503916 150892 503972 150948
rect 509292 153580 509348 153636
rect 506604 153356 506660 153412
rect 505596 153132 505652 153188
rect 505596 152796 505652 152852
rect 506828 153356 506884 153412
rect 506828 150220 506884 150276
rect 507948 153020 508004 153076
rect 508172 153020 508228 153076
rect 508172 150780 508228 150836
rect 511980 161756 512036 161812
rect 513324 159292 513380 159348
rect 514668 152236 514724 152292
rect 538524 172956 538580 173012
rect 550620 172956 550676 173012
rect 544572 172844 544628 172900
rect 556668 172844 556724 172900
rect 532476 171276 532532 171332
rect 526428 167804 526484 167860
rect 524076 164108 524132 164164
rect 521388 160636 521444 160692
rect 520044 160300 520100 160356
rect 518700 160188 518756 160244
rect 517356 159852 517412 159908
rect 522732 160524 522788 160580
rect 546588 161868 546644 161924
rect 524188 159404 524244 159460
rect 540876 159068 540932 159124
rect 524188 153692 524244 153748
rect 526764 156156 526820 156212
rect 525420 153244 525476 153300
rect 530796 156044 530852 156100
rect 528108 155820 528164 155876
rect 529452 155708 529508 155764
rect 537516 155484 537572 155540
rect 532140 153916 532196 153972
rect 534828 153132 534884 153188
rect 532588 152908 532644 152964
rect 532588 151004 532644 151060
rect 533484 152348 533540 152404
rect 544348 158956 544404 159012
rect 540876 154028 540932 154084
rect 544236 155596 544292 155652
rect 542892 153356 542948 153412
rect 540204 153020 540260 153076
rect 538860 152124 538916 152180
rect 541548 152908 541604 152964
rect 544348 154252 544404 154308
rect 549612 159180 549668 159236
rect 546588 154140 546644 154196
rect 548268 158844 548324 158900
rect 546924 154028 546980 154084
rect 545580 153692 545636 153748
rect 559468 403228 559524 403284
rect 559020 392364 559076 392420
rect 559020 391468 559076 391524
rect 559020 172284 559076 172340
rect 587132 443212 587188 443268
rect 583772 416780 583828 416836
rect 587132 407372 587188 407428
rect 583772 404012 583828 404068
rect 563612 402444 563668 402500
rect 559468 154476 559524 154532
rect 559580 397404 559636 397460
rect 559580 396508 559636 396564
rect 558908 154364 558964 154420
rect 550956 154252 551012 154308
rect 552300 154140 552356 154196
rect 590604 396508 590660 396564
rect 566972 394716 567028 394772
rect 562828 393372 562884 393428
rect 559692 393260 559748 393316
rect 559692 172732 559748 172788
rect 560252 205324 560308 205380
rect 566972 337484 567028 337540
rect 578732 393148 578788 393204
rect 578732 297836 578788 297892
rect 590492 392588 590548 392644
rect 562828 172956 562884 173012
rect 565292 284620 565348 284676
rect 590940 392252 590996 392308
rect 590604 364140 590660 364196
rect 590716 391468 590772 391524
rect 590940 350924 590996 350980
rect 590716 324492 590772 324548
rect 590492 258412 590548 258468
rect 587132 244972 587188 245028
rect 587132 169260 587188 169316
rect 565292 164332 565348 164388
rect 560252 162428 560308 162484
rect 560364 162092 560420 162148
rect 560140 157836 560196 157892
rect 559916 157500 559972 157556
rect 559804 157388 559860 157444
rect 559580 153804 559636 153860
rect 559692 157164 559748 157220
rect 552636 150668 552692 150724
rect 536172 149548 536228 149604
rect 501228 149212 501284 149268
rect 559468 149212 559524 149268
rect 559580 148652 559636 148708
rect 559692 142044 559748 142100
rect 560028 157052 560084 157108
rect 560028 140588 560084 140644
rect 560252 157612 560308 157668
rect 560252 136668 560308 136724
rect 560140 135100 560196 135156
rect 559916 134316 559972 134372
rect 559804 132524 559860 132580
rect 559580 124348 559636 124404
rect 559468 118412 559524 118468
rect 564508 161980 564564 162036
rect 561372 158732 561428 158788
rect 561148 157724 561204 157780
rect 561260 149436 561316 149492
rect 561260 142940 561316 142996
rect 561148 138236 561204 138292
rect 561596 152012 561652 152068
rect 561372 127260 561428 127316
rect 561484 150332 561540 150388
rect 560364 111580 560420 111636
rect 563164 150556 563220 150612
rect 561596 114716 561652 114772
rect 562828 149660 562884 149716
rect 561484 108444 561540 108500
rect 459452 102396 459508 102452
rect 457884 101388 457940 101444
rect 457772 92652 457828 92708
rect 423164 74396 423220 74452
rect 562940 148876 562996 148932
rect 563052 148764 563108 148820
rect 566188 160412 566244 160468
rect 564732 157276 564788 157332
rect 564508 122556 564564 122612
rect 564620 155372 564676 155428
rect 564732 130396 564788 130452
rect 566188 128828 566244 128884
rect 564620 119420 564676 119476
rect 563164 88060 563220 88116
rect 563052 86492 563108 86548
rect 562940 80220 562996 80276
rect 563500 81788 563556 81844
rect 562828 70812 562884 70868
rect 563388 72380 563444 72436
rect 422940 68796 422996 68852
rect 422716 60508 422772 60564
rect 563164 67676 563220 67732
rect 562940 59836 562996 59892
rect 422492 53564 422548 53620
rect 562828 58268 562884 58324
rect 562828 49868 562884 49924
rect 422044 49532 422100 49588
rect 356188 48636 356244 48692
rect 562940 48300 562996 48356
rect 354396 48188 354452 48244
rect 563276 62972 563332 63028
rect 563276 50316 563332 50372
rect 563388 48524 563444 48580
rect 563164 48188 563220 48244
rect 563724 69244 563780 69300
rect 563612 61404 563668 61460
rect 563724 48412 563780 48468
rect 563612 47964 563668 48020
rect 563500 45276 563556 45332
rect 289996 24332 290052 24388
rect 289772 4620 289828 4676
rect 277340 4060 277396 4116
rect 580636 4172 580692 4228
rect 582540 4172 582596 4228
rect 584444 4172 584500 4228
<< metal3 >>
rect 189634 591276 189644 591332
rect 189700 591276 209580 591332
rect 209636 591276 209646 591332
rect 560242 591276 560252 591332
rect 560308 591276 562604 591332
rect 562660 591276 562670 591332
rect 190642 591164 190652 591220
rect 190708 591164 231644 591220
rect 231700 591164 231710 591220
rect 193106 591052 193116 591108
rect 193172 591052 253708 591108
rect 253764 591052 253774 591108
rect 189186 590940 189196 590996
rect 189252 590940 297836 590996
rect 297892 590940 297902 590996
rect 193330 590828 193340 590884
rect 193396 590828 319900 590884
rect 319956 590828 319966 590884
rect 189298 590716 189308 590772
rect 189364 590716 364028 590772
rect 364084 590716 364094 590772
rect 386306 590716 386316 590772
rect 386372 590716 401436 590772
rect 401492 590716 401502 590772
rect 194226 590604 194236 590660
rect 194292 590604 430220 590660
rect 430276 590604 430286 590660
rect 452498 590604 452508 590660
rect 452564 590604 511308 590660
rect 511364 590604 511374 590660
rect 99474 590492 99484 590548
rect 99540 590492 141932 590548
rect 141988 590492 141998 590548
rect 186386 590492 186396 590548
rect 186452 590492 496412 590548
rect 496468 590492 496478 590548
rect 514882 590156 514892 590212
rect 514948 590156 518476 590212
rect 518532 590156 518542 590212
rect 584658 590156 584668 590212
rect 584724 590156 584762 590212
rect 189746 588812 189756 588868
rect 189812 588812 408268 588868
rect 408324 588812 408334 588868
rect 595560 588644 597000 588840
rect 590482 588588 590492 588644
rect 590548 588616 597000 588644
rect 590548 588588 595672 588616
rect 401426 587916 401436 587972
rect 401492 587916 407372 587972
rect 407428 587916 407438 587972
rect -960 587188 480 587384
rect -960 587160 179004 587188
rect 392 587132 179004 587160
rect 179060 587132 179070 587188
rect 184706 578732 184716 578788
rect 184772 578732 474348 578788
rect 474404 578732 474414 578788
rect 180450 577052 180460 577108
rect 180516 577052 540540 577108
rect 540596 577052 540606 577108
rect 183026 575484 183036 575540
rect 183092 575484 590492 575540
rect 590548 575484 590558 575540
rect 595560 575428 597000 575624
rect 189074 575372 189084 575428
rect 189140 575400 597000 575428
rect 189140 575372 595672 575400
rect -960 573076 480 573272
rect -960 573048 12572 573076
rect 392 573020 12572 573048
rect 12628 573020 12638 573076
rect 77298 572012 77308 572068
rect 77364 572012 175532 572068
rect 175588 572012 175598 572068
rect 189522 572012 189532 572068
rect 189588 572012 275772 572068
rect 275828 572012 275838 572068
rect 121314 570332 121324 570388
rect 121380 570332 172172 570388
rect 172228 570332 172238 570388
rect 189410 570332 189420 570388
rect 189476 570332 341964 570388
rect 342020 570332 342030 570388
rect 184706 567868 184716 567924
rect 184772 567868 590492 567924
rect 590548 567868 590558 567924
rect 407362 566972 407372 567028
rect 407428 566972 511420 567028
rect 511476 566972 511486 567028
rect 186274 565068 186284 565124
rect 186340 565068 190120 565124
rect 549864 565068 556108 565124
rect 556164 565068 556174 565124
rect 595560 562212 597000 562408
rect 585442 562156 585452 562212
rect 585508 562184 597000 562212
rect 585508 562156 595672 562184
rect 549864 560364 552748 560420
rect 552804 560364 552814 560420
rect -960 558964 480 559160
rect -960 558936 4172 558964
rect 392 558908 4172 558936
rect 4228 558908 4238 558964
rect 187842 557900 187852 557956
rect 187908 557900 190120 557956
rect 549864 555660 552748 555716
rect 552804 555660 552814 555716
rect 549864 550956 556220 551012
rect 556276 550956 556286 551012
rect 186162 550732 186172 550788
rect 186228 550732 190120 550788
rect 590482 549164 590492 549220
rect 590548 549192 595672 549220
rect 590548 549164 597000 549192
rect 595560 548968 597000 549164
rect 549864 546252 554428 546308
rect 554484 546252 554494 546308
rect -960 544852 480 545048
rect -960 544824 57932 544852
rect 392 544796 57932 544824
rect 57988 544796 57998 544852
rect 186050 543564 186060 543620
rect 186116 543564 190120 543620
rect 549864 541548 551068 541604
rect 551124 541548 551134 541604
rect 549864 536844 556444 536900
rect 556500 536844 556510 536900
rect 187730 536396 187740 536452
rect 187796 536396 190120 536452
rect 595560 535780 597000 535976
rect 565282 535724 565292 535780
rect 565348 535752 597000 535780
rect 565348 535724 595672 535752
rect 549864 532140 551180 532196
rect 551236 532140 551246 532196
rect -960 530740 480 530936
rect -960 530712 14252 530740
rect 392 530684 14252 530712
rect 14308 530684 14318 530740
rect 186386 529228 186396 529284
rect 186452 529228 190120 529284
rect 549864 527436 556332 527492
rect 556388 527436 556398 527492
rect 549378 522732 549388 522788
rect 549444 522732 549454 522788
rect 595560 522564 597000 522760
rect 568642 522508 568652 522564
rect 568708 522536 597000 522564
rect 568708 522508 595672 522536
rect 184482 522060 184492 522116
rect 184548 522060 190120 522116
rect 549864 518028 554540 518084
rect 554596 518028 554606 518084
rect -960 516628 480 516824
rect -960 516600 4284 516628
rect 392 516572 4284 516600
rect 4340 516572 4350 516628
rect 187170 514892 187180 514948
rect 187236 514892 190120 514948
rect 549864 513324 551292 513380
rect 551348 513324 551358 513380
rect 595560 509348 597000 509544
rect 590482 509292 590492 509348
rect 590548 509320 597000 509348
rect 590548 509292 595672 509320
rect 549836 508004 549892 508648
rect 549836 507948 550004 508004
rect 549948 507892 550004 507948
rect 549938 507836 549948 507892
rect 550004 507836 550014 507892
rect 187282 507724 187292 507780
rect 187348 507724 190120 507780
rect 549864 503916 554652 503972
rect 554708 503916 554718 503972
rect -960 502516 480 502712
rect -960 502488 56252 502516
rect 392 502460 56252 502488
rect 56308 502460 56318 502516
rect 183922 500556 183932 500612
rect 183988 500556 190120 500612
rect 549864 499212 554764 499268
rect 554820 499212 554830 499268
rect 595560 496132 597000 496328
rect 563602 496076 563612 496132
rect 563668 496104 597000 496132
rect 563668 496076 595672 496104
rect 549864 494508 551068 494564
rect 551124 494508 551134 494564
rect 188066 493388 188076 493444
rect 188132 493388 190120 493444
rect 549490 489804 549500 489860
rect 549556 489804 549566 489860
rect -960 488404 480 488600
rect -960 488376 15932 488404
rect 392 488348 15932 488376
rect 15988 488348 15998 488404
rect 187506 487228 187516 487284
rect 187572 487228 188860 487284
rect 188916 487228 188926 487284
rect 187506 486220 187516 486276
rect 187572 486220 190120 486276
rect 549500 484484 549556 485128
rect 549490 484428 549500 484484
rect 549556 484428 549566 484484
rect 595560 482916 597000 483112
rect 566962 482860 566972 482916
rect 567028 482888 597000 482916
rect 567028 482860 595672 482888
rect 549864 480396 551404 480452
rect 551460 480396 551470 480452
rect 187954 479052 187964 479108
rect 188020 479052 190120 479108
rect 549612 475524 549668 475720
rect 549602 475468 549612 475524
rect 549668 475468 549678 475524
rect -960 474292 480 474488
rect -960 474264 4396 474292
rect 392 474236 4396 474264
rect 4452 474236 4462 474292
rect 187394 471884 187404 471940
rect 187460 471884 190120 471940
rect 549864 470988 551516 471044
rect 551572 470988 551582 471044
rect 595560 469700 597000 469896
rect 590594 469644 590604 469700
rect 590660 469672 597000 469700
rect 590660 469644 595672 469672
rect 4162 469532 4172 469588
rect 4228 469532 177212 469588
rect 177268 469532 177278 469588
rect 4274 467852 4284 467908
rect 4340 467852 180572 467908
rect 180628 467852 180638 467908
rect 4386 466172 4396 466228
rect 4452 466172 175532 466228
rect 175588 466172 175598 466228
rect 549724 465780 549780 466312
rect 549714 465724 549724 465780
rect 549780 465724 549790 465780
rect 187618 464716 187628 464772
rect 187684 464716 190120 464772
rect 549864 461580 554988 461636
rect 555044 461580 555054 461636
rect -960 460180 480 460376
rect -960 460152 183932 460180
rect 392 460124 183932 460152
rect 183988 460124 183998 460180
rect 187842 457548 187852 457604
rect 187908 457548 190120 457604
rect 549864 456876 554876 456932
rect 554932 456876 554942 456932
rect 595560 456484 597000 456680
rect 570322 456428 570332 456484
rect 570388 456456 597000 456484
rect 570388 456428 595672 456456
rect 549864 452172 552860 452228
rect 552916 452172 552926 452228
rect 187506 450380 187516 450436
rect 187572 450380 190120 450436
rect 549864 447468 552972 447524
rect 553028 447468 553038 447524
rect -960 446068 480 446264
rect -960 446040 173852 446068
rect 392 446012 173852 446040
rect 173908 446012 173918 446068
rect 595560 443268 597000 443464
rect 187954 443212 187964 443268
rect 188020 443212 190120 443268
rect 587122 443212 587132 443268
rect 587188 443240 597000 443268
rect 587188 443212 595672 443240
rect 549864 442764 553084 442820
rect 553140 442764 553150 442820
rect 549864 438060 553196 438116
rect 553252 438060 553262 438116
rect 187282 436044 187292 436100
rect 187348 436044 190120 436100
rect 549864 433356 553308 433412
rect 553364 433356 553374 433412
rect -960 431956 480 432152
rect -960 431928 177324 431956
rect 392 431900 177324 431928
rect 177380 431900 177390 431956
rect 595560 430164 597000 430248
rect 590706 430108 590716 430164
rect 590772 430108 597000 430164
rect 595560 430024 597000 430108
rect 185378 428876 185388 428932
rect 185444 428876 190120 428932
rect 549836 428484 549892 428680
rect 549826 428428 549836 428484
rect 549892 428428 549902 428484
rect 549388 423444 549444 423976
rect 549378 423388 549388 423444
rect 549444 423388 549454 423444
rect 190642 421820 190652 421876
rect 190708 421820 190718 421876
rect 190652 421736 190708 421820
rect 549864 419244 551628 419300
rect 551684 419244 551694 419300
rect -960 417844 480 418040
rect -960 417816 181468 417844
rect 392 417788 181468 417816
rect 181524 417788 181534 417844
rect 595560 416836 597000 417032
rect 583762 416780 583772 416836
rect 583828 416808 597000 416836
rect 583828 416780 595672 416808
rect 178882 414540 178892 414596
rect 178948 414540 190120 414596
rect 549864 414540 551180 414596
rect 551236 414540 551246 414596
rect 143378 410732 143388 410788
rect 143444 410732 177324 410788
rect 177380 410732 177390 410788
rect 187842 410396 187852 410452
rect 187908 410396 341404 410452
rect 341460 410396 341470 410452
rect 359874 410060 359884 410116
rect 359940 410060 429660 410116
rect 429716 410060 429726 410116
rect 293458 409948 293468 410004
rect 293524 409948 405692 410004
rect 405748 409948 405758 410004
rect 56242 409836 56252 409892
rect 56308 409836 308028 409892
rect 308084 409836 308094 409892
rect 57922 409724 57932 409780
rect 57988 409724 302652 409780
rect 302708 409724 302718 409780
rect 187730 409612 187740 409668
rect 187796 409612 341292 409668
rect 341348 409612 341358 409668
rect 181458 409500 181468 409556
rect 181524 409500 318332 409556
rect 318388 409500 318780 409556
rect 318836 409500 318846 409556
rect 324818 409500 324828 409556
rect 324884 409500 551068 409556
rect 551124 409500 551134 409556
rect 183922 409388 183932 409444
rect 183988 409388 313404 409444
rect 313460 409388 313470 409444
rect 326610 409388 326620 409444
rect 326676 409388 554428 409444
rect 554484 409388 554494 409444
rect 178994 409276 179004 409332
rect 179060 409276 296492 409332
rect 296548 409276 296558 409332
rect 321234 409276 321244 409332
rect 321300 409276 551180 409332
rect 551236 409276 551246 409332
rect 55122 409164 55132 409220
rect 55188 409164 285516 409220
rect 285572 409164 285582 409220
rect 294354 409164 294364 409220
rect 294420 409164 554988 409220
rect 555044 409164 555054 409220
rect 193330 409052 193340 409108
rect 193396 409052 270396 409108
rect 270452 409052 270462 409108
rect 280018 409052 280028 409108
rect 280084 409052 549388 409108
rect 549444 409052 549454 409108
rect 187170 408940 187180 408996
rect 187236 408940 339276 408996
rect 339332 408940 339342 408996
rect 298834 408604 298844 408660
rect 298900 408604 391356 408660
rect 391412 408604 391422 408660
rect 304210 408492 304220 408548
rect 304276 408492 417452 408548
rect 417508 408492 417518 408548
rect 359538 408380 359548 408436
rect 359604 408380 484092 408436
rect 484148 408380 484158 408436
rect 340162 408268 340172 408324
rect 340228 408268 471996 408324
rect 472052 408268 472062 408324
rect 285506 408156 285516 408212
rect 285572 408156 291452 408212
rect 291508 408156 291518 408212
rect 391346 408156 391356 408212
rect 391412 408156 442428 408212
rect 442484 408156 442494 408212
rect 172162 408044 172172 408100
rect 172228 408044 286412 408100
rect 286468 408044 286478 408100
rect 353602 408044 353612 408100
rect 353668 408044 404796 408100
rect 404852 408044 404862 408100
rect 417442 408044 417452 408100
rect 417508 408044 458556 408100
rect 458612 408044 458622 408100
rect 189074 407932 189084 407988
rect 189140 407932 208348 407988
rect 208404 407932 208414 407988
rect 243478 407932 243516 407988
rect 243572 407932 243582 407988
rect 254258 407932 254268 407988
rect 254324 407932 357308 407988
rect 357364 407932 357374 407988
rect 359874 407932 359884 407988
rect 359940 407932 383292 407988
rect 383348 407932 383358 407988
rect 405682 407932 405692 407988
rect 405748 407932 426300 407988
rect 426356 407932 426366 407988
rect 453618 407932 453628 407988
rect 453684 407932 463932 407988
rect 463988 407932 463998 407988
rect 188850 407820 188860 407876
rect 188916 407820 281372 407876
rect 281428 407820 281438 407876
rect 351922 407820 351932 407876
rect 351988 407820 415548 407876
rect 415604 407820 415614 407876
rect 419972 407820 420924 407876
rect 420980 407820 420990 407876
rect 441858 407820 441868 407876
rect 441924 407820 480060 407876
rect 480116 407820 480126 407876
rect 419972 407764 420028 407820
rect 193106 407708 193116 407764
rect 193172 407708 276332 407764
rect 276388 407708 276398 407764
rect 352146 407708 352156 407764
rect 352212 407708 420028 407764
rect 421586 407708 421596 407764
rect 421652 407708 474684 407764
rect 474740 407708 474750 407764
rect 479602 407708 479612 407764
rect 479668 407708 490812 407764
rect 490868 407708 490878 407764
rect 182466 407596 182476 407652
rect 182532 407596 205884 407652
rect 205940 407596 205950 407652
rect 259634 407596 259644 407652
rect 259700 407596 315756 407652
rect 315812 407596 315822 407652
rect 358754 407596 358764 407652
rect 358820 407596 410172 407652
rect 410228 407596 410238 407652
rect 412402 407596 412412 407652
rect 412468 407596 485436 407652
rect 485492 407596 485502 407652
rect 486322 407596 486332 407652
rect 486388 407596 517692 407652
rect 517748 407596 517758 407652
rect 533782 407596 533820 407652
rect 533876 407596 533886 407652
rect 539158 407596 539196 407652
rect 539252 407596 539262 407652
rect 189186 407484 189196 407540
rect 189252 407484 212828 407540
rect 212884 407484 212894 407540
rect 248854 407484 248892 407540
rect 248948 407484 248958 407540
rect 275538 407484 275548 407540
rect 275604 407484 372540 407540
rect 372596 407484 372606 407540
rect 393138 407484 393148 407540
rect 393204 407484 544572 407540
rect 544628 407484 544638 407540
rect 103394 407372 103404 407428
rect 103460 407372 232764 407428
rect 232820 407372 356188 407428
rect 356244 407372 357196 407428
rect 357252 407372 357262 407428
rect 362002 407372 362012 407428
rect 362068 407372 528444 407428
rect 528500 407372 528510 407428
rect 557778 407372 557788 407428
rect 557844 407372 558908 407428
rect 558964 407372 587132 407428
rect 587188 407372 587198 407428
rect 355394 407260 355404 407316
rect 355460 407260 394044 407316
rect 394100 407260 394110 407316
rect 355170 407148 355180 407204
rect 355236 407148 388668 407204
rect 388724 407148 388734 407204
rect 238130 407036 238140 407092
rect 238196 407036 357196 407092
rect 357252 407036 357262 407092
rect 357298 406700 357308 406756
rect 357364 406700 357756 406756
rect 357812 406700 357822 406756
rect 227574 406588 227612 406644
rect 227668 406588 227678 406644
rect 265010 406588 265020 406644
rect 265076 406588 266252 406644
rect 266308 406588 266318 406644
rect 270358 406588 270396 406644
rect 270452 406588 270462 406644
rect 276294 406588 276332 406644
rect 276388 406588 276398 406644
rect 281334 406588 281372 406644
rect 281428 406588 281438 406644
rect 286374 406588 286412 406644
rect 286468 406588 286478 406644
rect 323362 406588 323372 406644
rect 323428 406588 324156 406644
rect 324212 406588 324222 406644
rect 334898 406588 334908 406644
rect 334964 406588 335916 406644
rect 335972 406588 335982 406644
rect 357186 406588 357196 406644
rect 357252 406588 357420 406644
rect 357476 406588 357486 406644
rect 357634 406588 357644 406644
rect 357700 406588 361788 406644
rect 361844 406588 361854 406644
rect 491362 406588 491372 406644
rect 491428 406588 496188 406644
rect 496244 406588 496254 406644
rect 309586 406364 309596 406420
rect 309652 406364 421596 406420
rect 421652 406364 421662 406420
rect 311378 406252 311388 406308
rect 311444 406252 441868 406308
rect 441924 406252 441934 406308
rect 288978 406140 288988 406196
rect 289044 406140 552972 406196
rect 553028 406140 553038 406196
rect 288194 406028 288204 406084
rect 288260 406028 553084 406084
rect 553140 406028 553150 406084
rect 285394 405916 285404 405972
rect 285460 405916 553196 405972
rect 553252 405916 553262 405972
rect 194226 405804 194236 405860
rect 194292 405804 211036 405860
rect 211092 405804 211102 405860
rect 281810 405804 281820 405860
rect 281876 405804 549836 405860
rect 549892 405804 549902 405860
rect 189298 405692 189308 405748
rect 189364 405692 211932 405748
rect 211988 405692 211998 405748
rect 283602 405692 283612 405748
rect 283668 405692 553308 405748
rect 553364 405692 553374 405748
rect 354162 405020 354172 405076
rect 354228 405020 459900 405076
rect 459956 405020 459966 405076
rect 359762 404908 359772 404964
rect 359828 404908 502236 404964
rect 502292 404908 502302 404964
rect 297042 404572 297052 404628
rect 297108 404572 437052 404628
rect 437108 404572 437118 404628
rect 300626 404460 300636 404516
rect 300692 404460 447804 404516
rect 447860 404460 447870 404516
rect 315746 404348 315756 404404
rect 315812 404348 357196 404404
rect 357252 404348 511308 404404
rect 511364 404348 511374 404404
rect 307794 404236 307804 404292
rect 307860 404236 469308 404292
rect 469364 404236 469374 404292
rect 186386 404124 186396 404180
rect 186452 404124 210140 404180
rect 210196 404124 210206 404180
rect 315858 404124 315868 404180
rect 315924 404124 554540 404180
rect 554596 404124 554606 404180
rect 204754 404012 204764 404068
rect 204820 404012 583772 404068
rect 583828 404012 583838 404068
rect -960 403732 480 403928
rect -960 403704 179228 403732
rect 392 403676 179228 403704
rect 179284 403676 179294 403732
rect 595560 403620 597000 403816
rect 561092 403592 597000 403620
rect 561092 403564 595672 403592
rect 359986 403452 359996 403508
rect 360052 403452 435708 403508
rect 435764 403452 435774 403508
rect 350466 403340 350476 403396
rect 350532 403340 478044 403396
rect 478100 403340 478110 403396
rect 561092 403284 561148 403564
rect 222002 403228 222012 403284
rect 222068 403228 559468 403284
rect 559524 403228 561148 403284
rect 332882 402892 332892 402948
rect 332948 402892 393148 402948
rect 393204 402892 393214 402948
rect 295250 402780 295260 402836
rect 295316 402780 431676 402836
rect 431732 402780 431742 402836
rect 306002 402668 306012 402724
rect 306068 402668 453628 402724
rect 453684 402668 453694 402724
rect 355282 402556 355292 402612
rect 355348 402556 552748 402612
rect 552804 402556 552814 402612
rect 206546 402444 206556 402500
rect 206612 402444 563612 402500
rect 563668 402444 563678 402500
rect 186050 402332 186060 402388
rect 186116 402332 590716 402388
rect 590772 402332 590782 402388
rect 352258 401772 352268 401828
rect 352324 401772 490140 401828
rect 490196 401772 490206 401828
rect 348898 401660 348908 401716
rect 348964 401660 544572 401716
rect 544628 401660 544638 401716
rect 184594 401548 184604 401604
rect 184660 401548 590940 401604
rect 590996 401548 591006 401604
rect 284498 401324 284508 401380
rect 284564 401324 399420 401380
rect 399476 401324 399486 401380
rect 312274 401212 312284 401268
rect 312340 401212 549948 401268
rect 550004 401212 550014 401268
rect 314066 401100 314076 401156
rect 314132 401100 551292 401156
rect 551348 401100 551358 401156
rect 310482 400988 310492 401044
rect 310548 400988 554652 401044
rect 554708 400988 554718 401044
rect 308690 400876 308700 400932
rect 308756 400876 554764 400932
rect 554820 400876 554830 400932
rect 292562 400764 292572 400820
rect 292628 400764 554876 400820
rect 554932 400764 554942 400820
rect 278226 400652 278236 400708
rect 278292 400652 551628 400708
rect 551684 400652 551694 400708
rect 361890 399980 361900 400036
rect 361956 399980 471884 400036
rect 471940 399980 471950 400036
rect 360546 399868 360556 399924
rect 360612 399868 496188 399924
rect 496244 399868 496254 399924
rect 210354 399756 210364 399812
rect 210420 399756 211260 399812
rect 211316 399756 211326 399812
rect 357522 399644 357532 399700
rect 357588 399644 367164 399700
rect 367220 399644 367230 399700
rect 302418 399532 302428 399588
rect 302484 399532 453180 399588
rect 453236 399532 453246 399588
rect 303314 399420 303324 399476
rect 303380 399420 549500 399476
rect 549556 399420 549566 399476
rect 301522 399308 301532 399364
rect 301588 399308 551404 399364
rect 551460 399308 551470 399364
rect 299730 399196 299740 399252
rect 299796 399196 549612 399252
rect 549668 399196 549678 399252
rect 190642 399084 190652 399140
rect 190708 399084 213724 399140
rect 213780 399084 213790 399140
rect 297938 399084 297948 399140
rect 298004 399084 551516 399140
rect 551572 399084 551582 399140
rect 173842 398972 173852 399028
rect 173908 398972 219996 399028
rect 220052 398972 220062 399028
rect 296146 398972 296156 399028
rect 296212 398972 549724 399028
rect 549780 398972 549790 399028
rect 359538 398300 359548 398356
rect 359604 398300 423612 398356
rect 423668 398300 423678 398356
rect 210354 398188 210364 398244
rect 210420 398188 471996 398244
rect 472052 398188 472062 398244
rect 519138 398076 519148 398132
rect 519204 398076 520380 398132
rect 520436 398076 520446 398132
rect 359202 397516 359212 397572
rect 359268 397516 514332 397572
rect 514388 397516 514398 397572
rect 180898 397404 180908 397460
rect 180964 397404 222012 397460
rect 222068 397404 222078 397460
rect 291666 397404 291676 397460
rect 291732 397404 352156 397460
rect 352212 397404 352222 397460
rect 352370 397404 352380 397460
rect 352436 397404 381276 397460
rect 381332 397404 381342 397460
rect 471874 397404 471884 397460
rect 471940 397404 559580 397460
rect 559636 397404 559646 397460
rect 14242 397292 14252 397348
rect 14308 397292 218204 397348
rect 218260 397292 218270 397348
rect 280914 397292 280924 397348
rect 280980 397292 355180 397348
rect 355236 397292 355246 397348
rect 358978 397292 358988 397348
rect 359044 397292 375228 397348
rect 375284 397292 375294 397348
rect 375442 397292 375452 397348
rect 375508 397292 511420 397348
rect 511476 397292 511486 397348
rect 357298 397180 357308 397236
rect 357364 397180 387324 397236
rect 387380 397180 387390 397236
rect 358642 397068 358652 397124
rect 358708 397068 393372 397124
rect 393428 397068 393438 397124
rect 355506 396956 355516 397012
rect 355572 396956 399420 397012
rect 399476 396956 399486 397012
rect 347218 396844 347228 396900
rect 347284 396844 411516 396900
rect 411572 396844 411582 396900
rect 526390 396844 526428 396900
rect 526484 396844 526494 396900
rect 340386 396732 340396 396788
rect 340452 396732 417564 396788
rect 417620 396732 417630 396788
rect 532438 396732 532476 396788
rect 532532 396732 532542 396788
rect 359650 396620 359660 396676
rect 359716 396620 508284 396676
rect 508340 396620 508350 396676
rect 556630 396620 556668 396676
rect 556724 396620 556734 396676
rect 550582 396508 550620 396564
rect 550676 396508 550686 396564
rect 559570 396508 559580 396564
rect 559636 396508 590604 396564
rect 590660 396508 590670 396564
rect 314850 396284 314860 396340
rect 314916 396284 479612 396340
rect 479668 396284 479678 396340
rect 316642 396172 316652 396228
rect 316708 396172 491372 396228
rect 491428 396172 491438 396228
rect 318434 396060 318444 396116
rect 318500 396060 501564 396116
rect 501620 396060 501630 396116
rect 320226 395948 320236 396004
rect 320292 395948 506940 396004
rect 506996 395948 507006 396004
rect 322018 395836 322028 395892
rect 322084 395836 512316 395892
rect 512372 395836 512382 395892
rect 180786 395724 180796 395780
rect 180852 395724 227612 395780
rect 227668 395724 227678 395780
rect 325602 395724 325612 395780
rect 325668 395724 523068 395780
rect 523124 395724 523134 395780
rect 12562 395612 12572 395668
rect 12628 395612 217196 395668
rect 217252 395612 217262 395668
rect 290658 395612 290668 395668
rect 290724 395612 552860 395668
rect 552916 395612 552926 395668
rect 362870 395052 362908 395108
rect 362964 395052 362974 395108
rect 357074 394940 357084 394996
rect 357140 394940 369180 394996
rect 369236 394940 369246 394996
rect 345314 394828 345324 394884
rect 345380 394828 453852 394884
rect 453908 394828 453918 394884
rect 538486 394828 538524 394884
rect 538580 394828 538590 394884
rect 202850 394716 202860 394772
rect 202916 394716 566972 394772
rect 567028 394716 567038 394772
rect 313058 394604 313068 394660
rect 313124 394604 412412 394660
rect 412468 394604 412478 394660
rect 277218 394492 277228 394548
rect 277284 394492 377916 394548
rect 377972 394492 377982 394548
rect 405430 394492 405468 394548
rect 405524 394492 405534 394548
rect 441718 394492 441756 394548
rect 441812 394492 441822 394548
rect 323810 394380 323820 394436
rect 323876 394380 486332 394436
rect 486388 394380 486398 394436
rect 361172 394268 431788 394324
rect 361172 394212 361228 394268
rect 182354 394156 182364 394212
rect 182420 394156 195132 394212
rect 195188 394156 195198 394212
rect 356738 394156 356748 394212
rect 356804 394156 361228 394212
rect 431732 394212 431788 394268
rect 443100 394268 447804 394324
rect 447860 394268 447870 394324
rect 455252 394268 465948 394324
rect 466004 394268 466014 394324
rect 431732 394156 438508 394212
rect 438564 394156 438574 394212
rect 443100 394100 443156 394268
rect 455252 394100 455308 394268
rect 184034 394044 184044 394100
rect 184100 394044 200508 394100
rect 200564 394044 200574 394100
rect 350690 394044 350700 394100
rect 350756 394044 443156 394100
rect 450212 394044 455308 394100
rect 450212 393988 450268 394044
rect 15922 393932 15932 393988
rect 15988 393932 218988 393988
rect 219044 393932 219054 393988
rect 438498 393932 438508 393988
rect 438564 393932 450268 393988
rect 343746 393372 343756 393428
rect 343812 393372 562828 393428
rect 562884 393372 562894 393428
rect 343522 393260 343532 393316
rect 343588 393260 559692 393316
rect 559748 393260 559758 393316
rect 201954 393148 201964 393204
rect 202020 393148 578732 393204
rect 578788 393148 578798 393204
rect 341842 392700 341852 392756
rect 341908 392700 362908 392756
rect 362964 392700 362974 392756
rect 329410 392588 329420 392644
rect 329476 392588 360444 392644
rect 360500 392588 360510 392644
rect 361890 392588 361900 392644
rect 361956 392588 590492 392644
rect 590548 392588 590558 392644
rect 350914 392476 350924 392532
rect 350980 392476 405468 392532
rect 405524 392476 405534 392532
rect 165442 392364 165452 392420
rect 165508 392364 214508 392420
rect 214564 392364 214574 392420
rect 327394 392364 327404 392420
rect 327460 392364 361788 392420
rect 361844 392364 361854 392420
rect 471986 392364 471996 392420
rect 472052 392364 559020 392420
rect 559076 392364 559086 392420
rect 33058 392252 33068 392308
rect 33124 392252 216300 392308
rect 216356 392252 216366 392308
rect 279010 392252 279020 392308
rect 279076 392252 359884 392308
rect 359940 392252 359950 392308
rect 362114 392252 362124 392308
rect 362180 392252 590940 392308
rect 590996 392252 591006 392308
rect 559010 391468 559020 391524
rect 559076 391468 590716 391524
rect 590772 391468 590782 391524
rect 216598 391356 216636 391412
rect 216692 391356 216702 391412
rect 178994 390908 179004 390964
rect 179060 390908 215068 390964
rect 215124 390908 215134 390964
rect 330978 390908 330988 390964
rect 331044 390908 358988 390964
rect 359044 390908 359054 390964
rect 179218 390796 179228 390852
rect 179284 390796 220780 390852
rect 220836 390796 220846 390852
rect 287970 390796 287980 390852
rect 288036 390796 358764 390852
rect 358820 390796 358830 390852
rect 141922 390684 141932 390740
rect 141988 390684 215404 390740
rect 215460 390684 215470 390740
rect 282594 390684 282604 390740
rect 282660 390684 355404 390740
rect 355460 390684 355470 390740
rect 186274 390572 186284 390628
rect 186340 390572 342972 390628
rect 343028 390572 343038 390628
rect 590930 390572 590940 390628
rect 590996 390600 595672 390628
rect 590996 390572 597000 390600
rect 595560 390376 597000 390572
rect 359846 389900 359884 389956
rect 359940 389900 359950 389956
rect -960 389620 480 389816
rect 359436 389620 360136 389676
rect -960 389592 4396 389620
rect 392 389564 4396 389592
rect 4452 389564 4462 389620
rect 355730 389564 355740 389620
rect 355796 389564 357532 389620
rect 357588 389564 359492 389620
rect 341954 389452 341964 389508
rect 342020 389452 359884 389508
rect 359940 389452 359950 389508
rect 340722 389340 340732 389396
rect 340788 389340 359548 389396
rect 359604 389340 359614 389396
rect 359874 389340 359884 389396
rect 359940 389340 359950 389396
rect 340946 389228 340956 389284
rect 341012 389228 359548 389284
rect 359604 389228 359614 389284
rect 359884 389172 359940 389340
rect 340498 389116 340508 389172
rect 340564 389116 359940 389172
rect 186050 388892 186060 388948
rect 186116 388892 342860 388948
rect 342916 388892 342926 388948
rect 349412 388892 359884 388948
rect 359940 388892 359950 388948
rect 349412 388836 349468 388892
rect 340050 388780 340060 388836
rect 340116 388780 349468 388836
rect 4162 388108 4172 388164
rect 4228 388108 329084 388164
rect 329140 388108 329532 388164
rect 329588 388108 329598 388164
rect 186162 387212 186172 387268
rect 186228 387212 343084 387268
rect 343140 387212 343150 387268
rect 111682 386764 111692 386820
rect 111748 386764 272188 386820
rect 272244 386764 272254 386820
rect 99922 386652 99932 386708
rect 99988 386652 273084 386708
rect 273140 386652 273150 386708
rect 38546 386540 38556 386596
rect 38612 386540 252028 386596
rect 252084 386540 252094 386596
rect 38434 386428 38444 386484
rect 38500 386428 253708 386484
rect 253764 386428 253774 386484
rect 318322 386092 318332 386148
rect 318388 386092 345548 386148
rect 345604 386092 345614 386148
rect 308242 385980 308252 386036
rect 308308 385980 342300 386036
rect 342356 385980 342366 386036
rect 303202 385868 303212 385924
rect 303268 385868 342076 385924
rect 342132 385868 342142 385924
rect 296482 385756 296492 385812
rect 296548 385756 338492 385812
rect 338548 385756 338558 385812
rect 290546 385644 290556 385700
rect 290612 385644 351932 385700
rect 351988 385644 351998 385700
rect 183922 385532 183932 385588
rect 183988 385532 260540 385588
rect 260596 385532 260606 385588
rect 286962 385532 286972 385588
rect 287028 385532 353612 385588
rect 353668 385532 353678 385588
rect 180674 385420 180684 385476
rect 180740 385420 264124 385476
rect 264180 385420 264190 385476
rect 246754 385308 246764 385364
rect 246820 385308 345212 385364
rect 345268 385308 345278 385364
rect 110002 385196 110012 385252
rect 110068 385196 265468 385252
rect 265524 385196 265534 385252
rect 103282 385084 103292 385140
rect 103348 385084 265916 385140
rect 265972 385084 265982 385140
rect 100370 384972 100380 385028
rect 100436 384972 267708 385028
rect 267764 384972 267774 385028
rect 103506 384860 103516 384916
rect 103572 384860 271292 384916
rect 271348 384860 271358 384916
rect 100146 384748 100156 384804
rect 100212 384748 270732 384804
rect 270788 384748 270798 384804
rect 40898 383964 40908 384020
rect 40964 383964 250572 384020
rect 250628 383964 250638 384020
rect 186386 383852 186396 383908
rect 186452 383852 343084 383908
rect 343140 383852 343150 383908
rect 359436 383796 360136 383852
rect 197362 383740 197372 383796
rect 197428 383740 262108 383796
rect 262164 383740 262174 383796
rect 357634 383740 357644 383796
rect 357700 383740 359492 383796
rect 199490 383628 199500 383684
rect 199556 383628 240716 383684
rect 240772 383628 240782 383684
rect 245186 383628 245196 383684
rect 245252 383628 339500 383684
rect 339556 383628 339566 383684
rect 118402 383516 118412 383572
rect 118468 383516 268828 383572
rect 268884 383516 268894 383572
rect 99922 383404 99932 383460
rect 99988 383404 263788 383460
rect 263844 383404 263854 383460
rect 106642 383292 106652 383348
rect 106708 383292 273868 383348
rect 273924 383292 273934 383348
rect 235106 383180 235116 383236
rect 235172 383180 340060 383236
rect 340116 383180 340126 383236
rect 12562 383068 12572 383124
rect 12628 383068 223468 383124
rect 223524 383068 223534 383124
rect 244962 383068 244972 383124
rect 245028 383068 349468 383124
rect 349524 383068 349534 383124
rect 352594 383068 352604 383124
rect 352660 383068 357644 383124
rect 357700 383068 357710 383124
rect 231606 382284 231644 382340
rect 231700 382284 231710 382340
rect 197362 382172 197372 382228
rect 197428 382172 198156 382228
rect 198212 382172 198222 382228
rect 199154 382172 199164 382228
rect 199220 382172 199836 382228
rect 199892 382172 199902 382228
rect 200834 382172 200844 382228
rect 200900 382172 201516 382228
rect 201572 382172 201582 382228
rect 208198 382172 208236 382228
rect 208292 382172 208302 382228
rect 209878 382172 209916 382228
rect 209972 382172 209982 382228
rect 230038 382172 230076 382228
rect 230132 382172 230142 382228
rect 231718 382172 231756 382228
rect 231812 382172 231822 382228
rect 332546 382172 332556 382228
rect 332612 382172 355292 382228
rect 355348 382172 355358 382228
rect 115042 382060 115052 382116
rect 115108 382060 257068 382116
rect 257124 382060 257134 382116
rect 277078 382060 277116 382116
rect 277172 382060 277182 382116
rect 287186 382060 287196 382116
rect 287252 382060 288204 382116
rect 288260 382060 288270 382116
rect 305638 382060 305676 382116
rect 305732 382060 305742 382116
rect 307318 382060 307356 382116
rect 307412 382060 307422 382116
rect 318322 382060 318332 382116
rect 318388 382060 319116 382116
rect 319172 382060 319182 382116
rect 320114 382060 320124 382116
rect 320180 382060 320796 382116
rect 320852 382060 320862 382116
rect 323586 382060 323596 382116
rect 323652 382060 324156 382116
rect 324212 382060 324222 382116
rect 329158 382060 329196 382116
rect 329252 382060 329262 382116
rect 330838 382060 330876 382116
rect 330932 382060 330942 382116
rect 334198 382060 334236 382116
rect 334292 382060 334302 382116
rect 196438 381948 196476 382004
rect 196532 381948 196542 382004
rect 198006 381948 198044 382004
rect 198100 381948 198110 382004
rect 199686 381948 199724 382004
rect 199780 381948 199790 382004
rect 201366 381948 201404 382004
rect 201460 381948 201470 382004
rect 204306 381948 204316 382004
rect 204372 381948 204876 382004
rect 204932 381948 204942 382004
rect 206098 381948 206108 382004
rect 206164 381948 206556 382004
rect 206612 381948 206622 382004
rect 206770 381948 206780 382004
rect 206836 381948 232204 382004
rect 232260 381948 232270 382004
rect 199826 381836 199836 381892
rect 199892 381836 232652 381892
rect 232708 381836 232718 381892
rect 240146 381836 240156 381892
rect 240212 381836 341180 381892
rect 341236 381836 341246 381892
rect 126802 381724 126812 381780
rect 126868 381724 257740 381780
rect 257796 381724 257806 381780
rect 120082 381612 120092 381668
rect 120148 381612 256060 381668
rect 256116 381612 256126 381668
rect 125122 381500 125132 381556
rect 125188 381500 267260 381556
rect 267316 381500 267326 381556
rect 335458 381500 335468 381556
rect 335524 381500 341628 381556
rect 341684 381500 341694 381556
rect 199602 381388 199612 381444
rect 199668 381388 206780 381444
rect 206836 381388 206846 381444
rect 239474 381388 239484 381444
rect 239540 381388 339612 381444
rect 339668 381388 339678 381444
rect 41122 380716 41132 380772
rect 41188 380716 250348 380772
rect 250404 380716 250414 380772
rect 190642 380604 190652 380660
rect 190708 380604 258748 380660
rect 258804 380604 258814 380660
rect 313282 380604 313292 380660
rect 313348 380604 352492 380660
rect 352548 380604 352558 380660
rect 184146 380492 184156 380548
rect 184212 380492 259532 380548
rect 259588 380492 259598 380548
rect 291442 380492 291452 380548
rect 291508 380492 336924 380548
rect 336980 380492 336990 380548
rect 180562 380380 180572 380436
rect 180628 380380 262332 380436
rect 262388 380380 262398 380436
rect 130162 380268 130172 380324
rect 130228 380268 223692 380324
rect 223748 380268 223758 380324
rect 32722 380156 32732 380212
rect 32788 380156 225484 380212
rect 225540 380156 225550 380212
rect 246642 380156 246652 380212
rect 246708 380156 341516 380212
rect 341572 380156 341582 380212
rect 29362 380044 29372 380100
rect 29428 380044 226828 380100
rect 226884 380044 226894 380100
rect 248546 380044 248556 380100
rect 248612 380044 346108 380100
rect 346164 380044 346174 380100
rect 27682 379932 27692 379988
rect 27748 379932 228956 379988
rect 229012 379932 229022 379988
rect 248658 379932 248668 379988
rect 248724 379932 347788 379988
rect 347844 379932 347854 379988
rect 20962 379820 20972 379876
rect 21028 379820 228060 379876
rect 228116 379820 228126 379876
rect 240594 379820 240604 379876
rect 240660 379820 351148 379876
rect 351204 379820 351214 379876
rect 176372 379708 182252 379764
rect 182308 379708 182318 379764
rect 210326 379708 210364 379764
rect 210420 379708 210430 379764
rect 236086 379708 236124 379764
rect 236180 379708 236190 379764
rect 242386 379708 242396 379764
rect 242452 379708 346444 379764
rect 346500 379708 346510 379764
rect 176372 379540 176428 379708
rect 38322 379484 38332 379540
rect 38388 379484 176428 379540
rect 182028 379596 196364 379652
rect 196420 379596 196430 379652
rect 202402 379596 202412 379652
rect 202468 379596 342972 379652
rect 343028 379596 343038 379652
rect 182028 379428 182084 379596
rect 182242 379484 182252 379540
rect 182308 379484 253148 379540
rect 253204 379484 253214 379540
rect 253362 379484 253372 379540
rect 253428 379484 254940 379540
rect 254996 379484 255006 379540
rect 261212 379484 336812 379540
rect 336868 379484 336878 379540
rect 40674 379372 40684 379428
rect 40740 379372 182084 379428
rect 195458 379372 195468 379428
rect 195524 379372 196140 379428
rect 196196 379372 196206 379428
rect 196354 379372 196364 379428
rect 196420 379372 221564 379428
rect 221620 379372 221630 379428
rect 221750 379372 221788 379428
rect 221844 379372 221854 379428
rect 222646 379372 222684 379428
rect 222740 379372 222750 379428
rect 225362 379372 225372 379428
rect 225428 379372 225438 379428
rect 235190 379372 235228 379428
rect 235284 379372 235294 379428
rect 236982 379372 237020 379428
rect 237076 379372 237086 379428
rect 238438 379372 238476 379428
rect 238532 379372 238542 379428
rect 243282 379372 243292 379428
rect 243348 379372 249396 379428
rect 249890 379372 249900 379428
rect 249956 379372 249966 379428
rect 250114 379372 250124 379428
rect 250180 379372 255836 379428
rect 255892 379372 255902 379428
rect 225372 379316 225428 379372
rect 14242 379260 14252 379316
rect 14308 379260 220108 379316
rect 220052 379204 220108 379260
rect 221676 379260 225428 379316
rect 231812 379260 249116 379316
rect 249172 379260 249182 379316
rect 221676 379204 221732 379260
rect 231812 379204 231868 379260
rect 249340 379204 249396 379372
rect 249900 379316 249956 379372
rect 261212 379316 261268 379484
rect 264450 379372 264460 379428
rect 264516 379372 270172 379428
rect 270228 379372 270238 379428
rect 278852 379372 352828 379428
rect 352884 379372 352894 379428
rect 249900 379260 261268 379316
rect 192322 379148 192332 379204
rect 192388 379148 202412 379204
rect 202468 379148 202478 379204
rect 220052 379148 221732 379204
rect 221890 379148 221900 379204
rect 221956 379148 231868 379204
rect 249330 379148 249340 379204
rect 249396 379148 249406 379204
rect 250002 379148 250012 379204
rect 250068 379148 270508 379204
rect 270452 379092 270508 379148
rect 278852 379092 278908 379372
rect 104962 379036 104972 379092
rect 105028 379036 264460 379092
rect 264516 379036 264526 379092
rect 270452 379036 278908 379092
rect 125234 378924 125244 378980
rect 125300 378924 222684 378980
rect 222740 378924 222750 378980
rect 243572 378924 253372 378980
rect 253428 378924 253438 378980
rect 197586 378812 197596 378868
rect 197652 378812 210364 378868
rect 210420 378812 210430 378868
rect 220052 378812 221788 378868
rect 221844 378812 221854 378868
rect 220052 378756 220108 378812
rect 130274 378700 130284 378756
rect 130340 378700 220108 378756
rect 243572 378644 243628 378924
rect 40226 378588 40236 378644
rect 40292 378588 243628 378644
rect 356402 378028 356412 378084
rect 356468 378028 357644 378084
rect 357700 378028 359492 378084
rect 359436 377972 360136 378028
rect 182466 377804 182476 377860
rect 182532 377804 190120 377860
rect 590482 377356 590492 377412
rect 590548 377384 595672 377412
rect 590548 377356 597000 377384
rect 4386 377132 4396 377188
rect 4452 377132 182252 377188
rect 182308 377132 182318 377188
rect 595560 377160 597000 377356
rect 187394 376460 187404 376516
rect 187460 376460 190120 376516
rect 354274 376236 354284 376292
rect 354340 376236 357868 376292
rect 357924 376236 357934 376292
rect 392 375704 4172 375732
rect -960 375676 4172 375704
rect 4228 375676 4238 375732
rect -960 375480 480 375676
rect 184146 375116 184156 375172
rect 184212 375116 190120 375172
rect 339864 373996 343756 374052
rect 343812 373996 343822 374052
rect 180674 373772 180684 373828
rect 180740 373772 190120 373828
rect 339864 373100 344092 373156
rect 344148 373100 344158 373156
rect 184034 372428 184044 372484
rect 184100 372428 190120 372484
rect 339864 372204 344204 372260
rect 344260 372204 344270 372260
rect 351026 372204 351036 372260
rect 351092 372204 356972 372260
rect 357028 372204 359492 372260
rect 359436 372148 360136 372204
rect 339864 371308 343532 371364
rect 343588 371308 343598 371364
rect 185602 371084 185612 371140
rect 185668 371084 190120 371140
rect 339864 370412 348572 370468
rect 348628 370412 348638 370468
rect 182242 369740 182252 369796
rect 182308 369740 190120 369796
rect 339864 369516 346892 369572
rect 346948 369516 346958 369572
rect 183810 368396 183820 368452
rect 183876 368396 190120 368452
rect 339836 368004 339892 368648
rect 339836 367948 339948 368004
rect 340004 367948 340014 368004
rect 339864 367724 351932 367780
rect 351988 367724 351998 367780
rect 189298 367052 189308 367108
rect 189364 367052 190120 367108
rect 345650 367052 345660 367108
rect 345716 367052 357196 367108
rect 357252 367052 359940 367108
rect 339864 366828 355292 366884
rect 355348 366828 355358 366884
rect 359884 366380 359940 367052
rect 359884 366324 360136 366380
rect 339864 365932 353612 365988
rect 353668 365932 353678 365988
rect 184594 365708 184604 365764
rect 184660 365708 190120 365764
rect 339864 365036 350252 365092
rect 350308 365036 350318 365092
rect 185490 364364 185500 364420
rect 185556 364364 190120 364420
rect 339864 364140 344764 364196
rect 344820 364140 344830 364196
rect 590594 364140 590604 364196
rect 590660 364168 595672 364196
rect 590660 364140 597000 364168
rect 595560 363944 597000 364140
rect 339864 363244 345324 363300
rect 345380 363244 345390 363300
rect 175896 363020 182476 363076
rect 182532 363020 182542 363076
rect 184772 363020 190120 363076
rect 184772 362964 184828 363020
rect 179666 362908 179676 362964
rect 179732 362908 184828 362964
rect 339864 362348 348684 362404
rect 348740 362348 348750 362404
rect 181234 361676 181244 361732
rect 181300 361676 190120 361732
rect -960 361396 480 361592
rect 339864 361452 347004 361508
rect 347060 361452 347070 361508
rect -960 361368 130284 361396
rect 392 361340 130284 361368
rect 130340 361340 130350 361396
rect 339864 360556 345436 360612
rect 345492 360556 345502 360612
rect 359436 360500 360136 360556
rect 340274 360444 340284 360500
rect 340340 360444 359492 360500
rect 176306 360332 176316 360388
rect 176372 360332 190120 360388
rect 175896 359660 187404 359716
rect 187460 359660 187470 359716
rect 339864 359660 352044 359716
rect 352100 359660 352110 359716
rect 340162 359548 340172 359604
rect 340228 359548 340284 359604
rect 340340 359548 340350 359604
rect 186386 358988 186396 359044
rect 186452 358988 190120 359044
rect 339864 358764 345436 358820
rect 345492 358764 345502 358820
rect 178882 358652 178892 358708
rect 178948 358652 185612 358708
rect 185668 358652 185678 358708
rect 339864 357868 355404 357924
rect 355460 357868 355470 357924
rect 177986 357644 177996 357700
rect 178052 357644 190120 357700
rect 339864 356972 353724 357028
rect 353780 356972 353790 357028
rect 175896 356300 184156 356356
rect 184212 356300 184222 356356
rect 184772 356300 190120 356356
rect 184772 356244 184828 356300
rect 179442 356188 179452 356244
rect 179508 356188 184828 356244
rect 339864 356076 350364 356132
rect 350420 356076 350430 356132
rect 189186 354956 189196 355012
rect 189252 354956 190120 355012
rect 339388 354564 339444 355208
rect 356514 354732 356524 354788
rect 356580 354732 359492 354788
rect 359436 354676 359772 354732
rect 359828 354676 360136 354732
rect 339378 354508 339388 354564
rect 339444 354508 339454 354564
rect 179106 354396 179116 354452
rect 179172 354396 182476 354452
rect 182532 354396 182542 354452
rect 339864 354284 348796 354340
rect 348852 354284 348862 354340
rect 183026 353612 183036 353668
rect 183092 353612 190120 353668
rect 339864 353388 345212 353444
rect 345268 353388 345278 353444
rect 175896 352940 180684 352996
rect 180740 352940 180750 352996
rect 339864 352492 348908 352548
rect 348964 352492 348974 352548
rect 181122 352268 181132 352324
rect 181188 352268 190120 352324
rect 339864 351596 347116 351652
rect 347172 351596 347182 351652
rect 179554 350924 179564 350980
rect 179620 350924 190120 350980
rect 590930 350924 590940 350980
rect 590996 350952 595672 350980
rect 590996 350924 597000 350952
rect 339864 350700 341852 350756
rect 341908 350700 341918 350756
rect 595560 350728 597000 350924
rect 184034 350364 184044 350420
rect 184100 350364 184110 350420
rect 184044 350308 184100 350364
rect 175868 350252 184100 350308
rect 175868 349608 175924 350252
rect 339864 349804 349020 349860
rect 349076 349804 349086 349860
rect 181010 349580 181020 349636
rect 181076 349580 190120 349636
rect 339864 348908 352156 348964
rect 352212 348908 352222 348964
rect 359436 348852 360136 348908
rect 357074 348796 357084 348852
rect 357140 348796 359492 348852
rect 182802 348236 182812 348292
rect 182868 348236 190120 348292
rect 339864 348012 355628 348068
rect 355684 348012 355694 348068
rect 357074 347788 357084 347844
rect 357140 347788 357756 347844
rect 357812 347788 357822 347844
rect -960 347284 480 347480
rect -960 347256 4172 347284
rect 392 347228 4172 347256
rect 4228 347228 4238 347284
rect 339864 347116 345884 347172
rect 345940 347116 345950 347172
rect 186274 346892 186284 346948
rect 186340 346892 190120 346948
rect 175896 346220 176428 346276
rect 176484 346220 180908 346276
rect 180964 346220 180974 346276
rect 339864 346220 354060 346276
rect 354116 346220 354126 346276
rect 184482 345548 184492 345604
rect 184548 345548 190120 345604
rect 339864 345324 343532 345380
rect 343588 345324 343598 345380
rect 339864 344428 342972 344484
rect 343028 344428 343038 344484
rect 180898 344204 180908 344260
rect 180964 344204 190120 344260
rect 339864 343532 344428 343588
rect 344484 343532 344494 343588
rect 348562 343084 348572 343140
rect 348628 343084 357644 343140
rect 357700 343084 359492 343140
rect 359436 343028 360136 343084
rect 175896 342860 178556 342916
rect 178612 342860 179004 342916
rect 179060 342860 179070 342916
rect 189074 342860 189084 342916
rect 189140 342860 190120 342916
rect 339864 342636 345660 342692
rect 345716 342636 345726 342692
rect 339864 341740 344092 341796
rect 344148 341740 344158 341796
rect 182914 341516 182924 341572
rect 182980 341516 190120 341572
rect 339864 340844 343196 340900
rect 343252 340844 343262 340900
rect 186162 340172 186172 340228
rect 186228 340172 190120 340228
rect 339864 339948 344316 340004
rect 344372 339948 344382 340004
rect 175896 339500 178108 339556
rect 178164 339500 178174 339556
rect 339864 339052 344092 339108
rect 344148 339052 344158 339108
rect 177874 338828 177884 338884
rect 177940 338828 190120 338884
rect 339864 338156 343644 338212
rect 343700 338156 343710 338212
rect 595560 337540 597000 337736
rect 175970 337484 175980 337540
rect 176036 337484 190120 337540
rect 566962 337484 566972 337540
rect 567028 337512 597000 337540
rect 567028 337484 595672 337512
rect 339266 337260 339276 337316
rect 339332 337260 339342 337316
rect 359436 337204 360136 337260
rect 359426 337148 359436 337204
rect 359492 337148 359502 337204
rect 339378 336364 339388 336420
rect 339444 336364 339454 336420
rect 175896 336140 178388 336196
rect 188850 336140 188860 336196
rect 188916 336140 190120 336196
rect 178332 336084 178388 336140
rect 178322 336028 178332 336084
rect 178388 336028 179116 336084
rect 179172 336028 179182 336084
rect 345538 336028 345548 336084
rect 345604 336028 359436 336084
rect 359492 336028 359502 336084
rect 339864 335468 354060 335524
rect 354116 335468 354126 335524
rect 182578 334796 182588 334852
rect 182644 334796 190120 334852
rect 339864 334572 344428 334628
rect 344484 334572 344494 334628
rect 339864 333676 355628 333732
rect 355684 333676 355694 333732
rect 176082 333452 176092 333508
rect 176148 333452 190120 333508
rect 392 333368 4172 333396
rect -960 333340 4172 333368
rect 4228 333340 4238 333396
rect -960 333144 480 333340
rect 175896 332780 178220 332836
rect 178276 332780 184044 332836
rect 184100 332780 184110 332836
rect 339864 332780 350364 332836
rect 350420 332780 350430 332836
rect 184370 332108 184380 332164
rect 184436 332108 190120 332164
rect 339864 331884 352268 331940
rect 352324 331884 352334 331940
rect 359436 331380 360136 331436
rect 359436 331044 359492 331380
rect 339864 330988 348572 331044
rect 348628 330988 348638 331044
rect 352482 330988 352492 331044
rect 352548 330988 359436 331044
rect 359492 330988 359502 331044
rect 182690 330764 182700 330820
rect 182756 330764 190120 330820
rect 182354 330204 182364 330260
rect 182420 330204 182430 330260
rect 182364 330148 182420 330204
rect 175868 330092 178444 330148
rect 178500 330092 182420 330148
rect 339864 330092 346780 330148
rect 346836 330092 346846 330148
rect 175868 329448 175924 330092
rect 176194 329420 176204 329476
rect 176260 329420 190120 329476
rect 339864 329196 346668 329252
rect 346724 329196 346734 329252
rect 339864 328300 353948 328356
rect 354004 328300 354014 328356
rect 184258 328076 184268 328132
rect 184324 328076 190120 328132
rect 339864 327404 350476 327460
rect 350532 327404 350542 327460
rect 188738 326732 188748 326788
rect 188804 326732 190120 326788
rect 339864 326508 348684 326564
rect 348740 326508 348750 326564
rect 175896 326060 178892 326116
rect 178948 326060 178958 326116
rect 339864 325612 352380 325668
rect 352436 325612 352446 325668
rect 356178 325612 356188 325668
rect 356244 325612 357868 325668
rect 357924 325612 359492 325668
rect 359436 325556 360136 325612
rect 181346 325388 181356 325444
rect 181412 325388 190120 325444
rect 339864 324716 347900 324772
rect 347956 324716 347966 324772
rect 590706 324492 590716 324548
rect 590772 324520 595672 324548
rect 590772 324492 597000 324520
rect 595560 324296 597000 324492
rect 190652 323428 190708 324072
rect 339864 323820 348796 323876
rect 348852 323820 348862 323876
rect 190642 323372 190652 323428
rect 190708 323372 190718 323428
rect 339864 322924 350700 322980
rect 350756 322924 350766 322980
rect 175298 322700 175308 322756
rect 175364 322700 180796 322756
rect 180852 322700 180862 322756
rect 187394 322700 187404 322756
rect 187460 322700 190120 322756
rect 176372 322364 179788 322420
rect 140242 322028 140252 322084
rect 140308 322028 168028 322084
rect 168084 322028 168094 322084
rect 176372 321972 176428 322364
rect 179732 322196 179788 322364
rect 183810 322252 183820 322308
rect 183876 322252 183886 322308
rect 183820 322196 183876 322252
rect 179732 322140 183876 322196
rect 339864 322028 353612 322084
rect 353668 322028 353678 322084
rect 152786 321916 152796 321972
rect 152852 321916 176428 321972
rect 113362 321804 113372 321860
rect 113428 321804 175308 321860
rect 175364 321804 175374 321860
rect 143602 321692 143612 321748
rect 143668 321692 178892 321748
rect 178948 321692 178958 321748
rect 168018 321580 168028 321636
rect 168084 321580 178556 321636
rect 178612 321580 178622 321636
rect 174514 321356 174524 321412
rect 174580 321356 190120 321412
rect 339864 321132 348012 321188
rect 348068 321132 348078 321188
rect 339864 320236 348124 320292
rect 348180 320236 348190 320292
rect 115154 320124 115164 320180
rect 115220 320124 178108 320180
rect 178164 320124 178174 320180
rect 174626 320012 174636 320068
rect 174692 320012 190120 320068
rect 342066 319788 342076 319844
rect 342132 319788 359492 319844
rect 359436 319732 360108 319788
rect 360164 319732 360174 319788
rect 339864 319340 344540 319396
rect 344596 319340 344606 319396
rect -960 319060 480 319256
rect -960 319032 125244 319060
rect 392 319004 125244 319032
rect 125300 319004 125310 319060
rect 174402 318668 174412 318724
rect 174468 318668 190120 318724
rect 339266 318444 339276 318500
rect 339332 318444 339342 318500
rect 339864 317548 359884 317604
rect 359940 317548 359950 317604
rect 177874 317324 177884 317380
rect 177940 317324 190120 317380
rect 339864 316652 353724 316708
rect 353780 316652 353790 316708
rect 179666 315980 179676 316036
rect 179732 315980 190120 316036
rect 339864 315756 346220 315812
rect 346276 315756 346286 315812
rect 339864 314860 342188 314916
rect 342244 314860 342254 314916
rect 184370 314636 184380 314692
rect 184436 314636 190120 314692
rect 339864 313964 349580 314020
rect 349636 313964 349646 314020
rect 359436 313908 360136 313964
rect 359436 313348 359492 313908
rect 177986 313292 177996 313348
rect 178052 313292 190120 313348
rect 339378 313292 339388 313348
rect 339444 313292 351260 313348
rect 351316 313292 358988 313348
rect 359044 313292 359492 313348
rect 339864 313068 352828 313124
rect 352884 313068 352894 313124
rect 339864 312172 351932 312228
rect 351988 312172 351998 312228
rect 174290 311948 174300 312004
rect 174356 311948 190120 312004
rect 339864 311276 355292 311332
rect 355348 311276 355358 311332
rect 595560 311108 597000 311304
rect 590482 311052 590492 311108
rect 590548 311080 597000 311108
rect 590548 311052 595672 311080
rect 185826 310604 185836 310660
rect 185892 310604 190120 310660
rect 339864 310380 346332 310436
rect 346388 310380 346398 310436
rect 339266 309820 339276 309876
rect 339332 309820 339500 309876
rect 339556 309820 339566 309876
rect 339864 309484 347788 309540
rect 347844 309484 347854 309540
rect 190418 309260 190428 309316
rect 190484 309260 190494 309316
rect 339864 308588 351148 308644
rect 351204 308588 351214 308644
rect 359436 308084 360136 308140
rect 357298 308028 357308 308084
rect 357364 308028 359492 308084
rect 357980 307972 358036 308028
rect 185714 307916 185724 307972
rect 185780 307916 190120 307972
rect 357970 307916 357980 307972
rect 358036 307916 358046 307972
rect 339864 307692 354620 307748
rect 354676 307692 354686 307748
rect 339864 306796 349692 306852
rect 349748 306796 349758 306852
rect 4162 306572 4172 306628
rect 4228 306572 168812 306628
rect 168868 306572 168878 306628
rect 181234 306572 181244 306628
rect 181300 306572 190120 306628
rect 339864 305900 352492 305956
rect 352548 305900 352558 305956
rect 350802 305676 350812 305732
rect 350868 305676 352604 305732
rect 352660 305676 352670 305732
rect 184482 305228 184492 305284
rect 184548 305228 190120 305284
rect -960 304948 480 305144
rect 339266 305004 339276 305060
rect 339332 305004 339342 305060
rect -960 304920 167244 304948
rect 392 304892 167244 304920
rect 167300 304892 167310 304948
rect 339864 304108 354284 304164
rect 354340 304108 354350 304164
rect 62402 303996 62412 304052
rect 62468 303996 63756 304052
rect 63812 303996 63822 304052
rect 77410 303996 77420 304052
rect 77476 303996 78876 304052
rect 78932 303996 78942 304052
rect 92418 303996 92428 304052
rect 92484 303996 93996 304052
rect 94052 303996 94062 304052
rect 187730 303884 187740 303940
rect 187796 303884 190120 303940
rect 339602 303212 339612 303268
rect 339668 303212 339678 303268
rect 186946 302540 186956 302596
rect 187012 302540 190120 302596
rect 47394 302428 47404 302484
rect 47460 302428 143612 302484
rect 143668 302428 143678 302484
rect 339864 302316 354172 302372
rect 354228 302316 354238 302372
rect 359436 302260 360136 302316
rect 350578 302204 350588 302260
rect 350644 302204 350812 302260
rect 350868 302204 359492 302260
rect 359100 302148 359156 302204
rect 359090 302092 359100 302148
rect 359156 302092 359166 302148
rect 10994 301532 11004 301588
rect 11060 301532 173964 301588
rect 174020 301532 174030 301588
rect 339864 301420 352156 301476
rect 352212 301420 352222 301476
rect 186834 301196 186844 301252
rect 186900 301196 190120 301252
rect 339864 300524 355740 300580
rect 355796 300524 355806 300580
rect 161298 299852 161308 299908
rect 161364 299852 182252 299908
rect 182308 299852 182318 299908
rect 182914 299852 182924 299908
rect 182980 299852 190120 299908
rect 339864 299628 349468 299684
rect 349412 299572 349468 299628
rect 349412 299516 356524 299572
rect 356580 299516 356590 299572
rect 339864 298732 345660 298788
rect 345716 298732 345726 298788
rect 187058 298508 187068 298564
rect 187124 298508 190120 298564
rect 595560 297892 597000 298088
rect 339864 297836 342412 297892
rect 342468 297836 342478 297892
rect 578722 297836 578732 297892
rect 578788 297864 597000 297892
rect 578788 297836 595672 297864
rect 187618 297164 187628 297220
rect 187684 297164 190120 297220
rect 339864 296940 346892 296996
rect 346948 296940 346958 296996
rect 4162 296604 4172 296660
rect 4228 296604 172284 296660
rect 172340 296604 172350 296660
rect 186498 296492 186508 296548
rect 186564 296492 187516 296548
rect 187572 296492 187582 296548
rect 346322 296492 346332 296548
rect 346388 296492 347676 296548
rect 347732 296492 347742 296548
rect 350578 296492 350588 296548
rect 350644 296492 355740 296548
rect 355796 296492 355806 296548
rect 359436 296436 360136 296492
rect 357858 296380 357868 296436
rect 357924 296380 359324 296436
rect 359380 296380 359492 296436
rect 99960 296044 165452 296100
rect 165508 296044 165518 296100
rect 339864 296044 359884 296100
rect 359940 296044 359950 296100
rect 187394 295820 187404 295876
rect 187460 295820 190120 295876
rect 340274 295708 340284 295764
rect 340340 295708 357868 295764
rect 357924 295708 357934 295764
rect 187842 295596 187852 295652
rect 187908 295596 187964 295652
rect 188020 295596 188030 295652
rect 339864 295148 342972 295204
rect 343028 295148 351260 295204
rect 351316 295148 351326 295204
rect 341394 294812 341404 294868
rect 341460 294812 353836 294868
rect 353892 294812 353902 294868
rect 187506 294476 187516 294532
rect 187572 294476 190120 294532
rect 339864 294252 341404 294308
rect 341460 294252 341470 294308
rect 339836 293188 339892 293384
rect 190092 292628 190148 293160
rect 339836 293132 343084 293188
rect 343140 293132 354732 293188
rect 354788 293132 354798 293188
rect 190082 292572 190092 292628
rect 190148 292572 190158 292628
rect 339864 292460 342748 292516
rect 342804 292460 342814 292516
rect 121762 291788 121772 291844
rect 121828 291788 190120 291844
rect 339864 291564 341292 291620
rect 341348 291564 349468 291620
rect 349412 291508 349468 291564
rect 349412 291452 353948 291508
rect 354004 291452 354014 291508
rect -960 290836 480 291032
rect 339836 290892 343084 290948
rect 343140 290892 349468 290948
rect -960 290808 4172 290836
rect 392 290780 4172 290808
rect 4228 290780 4238 290836
rect 339836 290696 339892 290892
rect 349412 290836 349468 290892
rect 349412 290780 352044 290836
rect 352100 290780 352110 290836
rect 342038 290668 342076 290724
rect 342132 290668 358876 290724
rect 358932 290668 359492 290724
rect 359436 290612 360136 290668
rect 138562 290444 138572 290500
rect 138628 290444 190120 290500
rect 99960 290220 165676 290276
rect 165732 290220 165742 290276
rect 169138 289772 169148 289828
rect 169204 289772 187292 289828
rect 187348 289772 187358 289828
rect 339864 289772 342860 289828
rect 342916 289772 355516 289828
rect 355572 289772 355582 289828
rect 167122 289100 167132 289156
rect 167188 289100 190120 289156
rect 143602 288988 143612 289044
rect 143668 288988 149548 289044
rect 149492 288932 149548 288988
rect 149492 288876 151116 288932
rect 151172 288876 151182 288932
rect 339266 288876 339276 288932
rect 339332 288876 342860 288932
rect 342916 288876 342926 288932
rect 188066 288428 188076 288484
rect 188132 288428 190652 288484
rect 190708 288428 190718 288484
rect 339864 287980 342748 288036
rect 342804 287980 342814 288036
rect 120082 287756 120092 287812
rect 120148 287756 190120 287812
rect 339864 287084 341292 287140
rect 341348 287084 341358 287140
rect 168802 286636 168812 286692
rect 168868 286636 186508 286692
rect 186564 286636 188076 286692
rect 188132 286636 188142 286692
rect 103618 286524 103628 286580
rect 103684 286524 176428 286580
rect 176484 286524 176494 286580
rect 173012 286412 190120 286468
rect 173012 286356 173068 286412
rect 113362 286300 113372 286356
rect 113428 286300 173068 286356
rect 339836 285796 339892 286216
rect 187842 285740 187852 285796
rect 187908 285740 190540 285796
rect 190596 285740 190606 285796
rect 339836 285740 354508 285796
rect 354564 285740 354574 285796
rect 182354 285628 182364 285684
rect 182420 285628 183932 285684
rect 183988 285628 183998 285684
rect 187142 285628 187180 285684
rect 187236 285628 187246 285684
rect 118402 285404 118412 285460
rect 118468 285404 190148 285460
rect 151218 285292 151228 285348
rect 151284 285292 165452 285348
rect 165508 285292 165518 285348
rect 190092 285096 190148 285404
rect 339388 284788 339444 285320
rect 355394 284844 355404 284900
rect 355460 284844 356860 284900
rect 356916 284844 359492 284900
rect 359436 284788 360136 284844
rect 339378 284732 339388 284788
rect 339444 284732 342748 284788
rect 342804 284732 342814 284788
rect 346210 284732 346220 284788
rect 346276 284732 347564 284788
rect 347620 284732 347630 284788
rect 595560 284676 597000 284872
rect 565282 284620 565292 284676
rect 565348 284648 597000 284676
rect 565348 284620 595672 284648
rect 99960 284396 103404 284452
rect 103460 284396 103470 284452
rect 339836 284116 339892 284424
rect 339836 284060 346220 284116
rect 346276 284060 358876 284116
rect 358932 284060 358942 284116
rect 165928 283948 169148 284004
rect 169204 283948 169214 284004
rect 342738 283948 342748 284004
rect 342804 283948 355964 284004
rect 356020 283948 356030 284004
rect 185602 283836 185612 283892
rect 185668 283836 187404 283892
rect 187460 283836 187470 283892
rect 348002 283836 348012 283892
rect 348068 283836 349132 283892
rect 349188 283836 349198 283892
rect 172274 283724 172284 283780
rect 172340 283724 190120 283780
rect 348114 283724 348124 283780
rect 348180 283724 349356 283780
rect 349412 283724 349422 283780
rect 182466 283612 182476 283668
rect 182532 283612 187628 283668
rect 187684 283612 187694 283668
rect 339864 283500 348236 283556
rect 348292 283500 348302 283556
rect 339864 282604 341292 282660
rect 341348 282604 341358 282660
rect 167234 282380 167244 282436
rect 167300 282380 190120 282436
rect 186498 282156 186508 282212
rect 186564 282156 187964 282212
rect 188020 282156 188030 282212
rect 352818 282156 352828 282212
rect 352884 282156 354396 282212
rect 354452 282156 354462 282212
rect 165928 281932 182364 281988
rect 182420 281932 182430 281988
rect 175634 281372 175644 281428
rect 175700 281372 187516 281428
rect 187572 281372 187582 281428
rect 339276 281204 339332 281736
rect 339266 281148 339276 281204
rect 339332 281148 339948 281204
rect 340004 281148 340014 281204
rect 168802 281036 168812 281092
rect 168868 281036 190120 281092
rect 344372 280924 349468 280980
rect 339304 280840 341068 280868
rect 339276 280812 341068 280840
rect 187142 280476 187180 280532
rect 187236 280476 187246 280532
rect 186274 280364 186284 280420
rect 186340 280364 187292 280420
rect 187348 280364 187358 280420
rect 190642 280364 190652 280420
rect 190708 280364 190718 280420
rect 190652 279972 190708 280364
rect 339276 280196 339332 280812
rect 341012 280756 341068 280812
rect 344372 280756 344428 280924
rect 341012 280700 344428 280756
rect 349412 280756 349468 280924
rect 349412 280700 353836 280756
rect 353892 280700 353902 280756
rect 339938 280588 339948 280644
rect 340004 280588 358652 280644
rect 358708 280588 358718 280644
rect 354722 280476 354732 280532
rect 354788 280476 355964 280532
rect 356020 280476 356030 280532
rect 354610 280364 354620 280420
rect 354676 280364 356076 280420
rect 356132 280364 356142 280420
rect 339266 280140 339276 280196
rect 339332 280140 339342 280196
rect 165928 279916 190708 279972
rect 182242 279692 182252 279748
rect 182308 279692 190120 279748
rect 339388 279636 339444 279944
rect 339378 279580 339388 279636
rect 339444 279580 339454 279636
rect 339388 279300 339444 279580
rect 165442 279244 165452 279300
rect 165508 279244 168140 279300
rect 168196 279244 168206 279300
rect 339388 279244 349468 279300
rect 173012 279020 186284 279076
rect 186340 279020 186350 279076
rect 339864 279020 342748 279076
rect 342804 279020 342814 279076
rect 173012 278964 173068 279020
rect 168130 278908 168140 278964
rect 168196 278908 173068 278964
rect 349412 278964 349468 279244
rect 359436 278964 360136 279020
rect 349412 278908 355404 278964
rect 355460 278908 355470 278964
rect 358754 278908 358764 278964
rect 358820 278908 359492 278964
rect 165442 278796 165452 278852
rect 165508 278796 174636 278852
rect 174692 278796 174702 278852
rect 342850 278796 342860 278852
rect 342916 278796 344316 278852
rect 344372 278796 344382 278852
rect 99960 278572 113372 278628
rect 113428 278572 113438 278628
rect 177314 278348 177324 278404
rect 177380 278348 190120 278404
rect 339864 278124 341404 278180
rect 341460 278124 341470 278180
rect 168018 278012 168028 278068
rect 168084 278012 185388 278068
rect 185444 278012 185454 278068
rect 165928 277900 168812 277956
rect 168868 277900 168878 277956
rect 165666 277228 165676 277284
rect 165732 277228 168028 277284
rect 168084 277228 168094 277284
rect 185378 277228 185388 277284
rect 185444 277228 187292 277284
rect 187348 277228 187358 277284
rect 339864 277228 341740 277284
rect 341796 277228 341806 277284
rect 175522 277004 175532 277060
rect 175588 277004 190120 277060
rect -960 276724 480 276920
rect -960 276696 12572 276724
rect 392 276668 12572 276696
rect 12628 276668 12638 276724
rect 339864 276332 341516 276388
rect 341572 276332 341582 276388
rect 174626 275996 174636 276052
rect 174692 275996 177212 276052
rect 177268 275996 177278 276052
rect 165928 275884 190540 275940
rect 190596 275884 190606 275940
rect 180562 275660 180572 275716
rect 180628 275660 190120 275716
rect 342738 275548 342748 275604
rect 342804 275548 344652 275604
rect 344708 275548 344718 275604
rect 339714 275436 339724 275492
rect 339780 275436 339790 275492
rect 339826 274540 339836 274596
rect 339892 274540 339902 274596
rect 177202 274316 177212 274372
rect 177268 274316 190120 274372
rect 165928 273868 185724 273924
rect 185780 273868 185790 273924
rect 339864 273644 342860 273700
rect 342916 273644 342926 273700
rect 359436 273140 360136 273196
rect 356738 273084 356748 273140
rect 356804 273084 357420 273140
rect 357476 273084 359492 273140
rect 173954 272972 173964 273028
rect 174020 272972 190120 273028
rect 356850 272972 356860 273028
rect 356916 272972 358764 273028
rect 358820 272972 358830 273028
rect 99960 272748 103628 272804
rect 103684 272748 103694 272804
rect 339864 272748 342972 272804
rect 343028 272748 343038 272804
rect 173012 272076 181356 272132
rect 181412 272076 182476 272132
rect 182532 272076 182542 272132
rect 344530 272076 344540 272132
rect 344596 272076 345996 272132
rect 346052 272076 346062 272132
rect 173012 271908 173068 272076
rect 165928 271852 173068 271908
rect 339864 271852 349580 271908
rect 349636 271852 349646 271908
rect 175522 271628 175532 271684
rect 175588 271628 190120 271684
rect 595560 271460 597000 271656
rect 590594 271404 590604 271460
rect 590660 271432 597000 271460
rect 590660 271404 595672 271432
rect 339864 270956 342860 271012
rect 342916 270956 342926 271012
rect 177314 270284 177324 270340
rect 177380 270284 190120 270340
rect 339266 270060 339276 270116
rect 339332 270060 339342 270116
rect 165928 269836 170492 269892
rect 170548 269836 170558 269892
rect 339864 269164 342972 269220
rect 343028 269164 343038 269220
rect 189634 268940 189644 268996
rect 189700 268940 190120 268996
rect 174626 268716 174636 268772
rect 174692 268716 175644 268772
rect 175700 268716 175710 268772
rect 357410 268716 357420 268772
rect 357476 268716 357756 268772
rect 357812 268716 357822 268772
rect 339864 268268 351372 268324
rect 351428 268268 351438 268324
rect 165900 267204 165956 267848
rect 189522 267596 189532 267652
rect 189588 267596 190120 267652
rect 339266 267372 339276 267428
rect 339332 267372 339342 267428
rect 357410 267372 357420 267428
rect 357476 267372 359492 267428
rect 359436 267316 360136 267372
rect 165900 267148 174636 267204
rect 174692 267148 174702 267204
rect 99960 266924 140252 266980
rect 140308 266924 140318 266980
rect 339864 266476 343084 266532
rect 343140 266476 343150 266532
rect 189410 266252 189420 266308
rect 189476 266252 190120 266308
rect 165928 265804 186396 265860
rect 186452 265804 186462 265860
rect 339864 265580 354620 265636
rect 354676 265580 354686 265636
rect 177202 265468 177212 265524
rect 177268 265468 181468 265524
rect 181524 265468 181534 265524
rect 189746 264908 189756 264964
rect 189812 264908 190120 264964
rect 339864 264684 343308 264740
rect 343364 264684 343374 264740
rect 344306 264572 344316 264628
rect 344372 264572 359548 264628
rect 359604 264572 359614 264628
rect 165928 263788 168140 263844
rect 168196 263788 168206 263844
rect 339864 263788 346108 263844
rect 346164 263788 346174 263844
rect 184706 263564 184716 263620
rect 184772 263564 190120 263620
rect 339864 262892 342748 262948
rect 342804 262892 342814 262948
rect 392 262808 4172 262836
rect -960 262780 4172 262808
rect 4228 262780 4238 262836
rect -960 262584 480 262780
rect 180450 262220 180460 262276
rect 180516 262220 190120 262276
rect 165928 261772 168028 261828
rect 168084 261772 168094 261828
rect 339276 261492 339332 262024
rect 359436 261492 360136 261548
rect 339266 261436 339276 261492
rect 339332 261436 339342 261492
rect 357532 261436 359492 261492
rect 357532 261380 357588 261436
rect 357522 261324 357532 261380
rect 357588 261324 357598 261380
rect 99960 261100 115164 261156
rect 115220 261100 115230 261156
rect 339864 261100 341404 261156
rect 341460 261100 341470 261156
rect 183026 260876 183036 260932
rect 183092 260876 190120 260932
rect 339266 260204 339276 260260
rect 339332 260204 339342 260260
rect 339266 259980 339276 260036
rect 339332 259980 339388 260036
rect 339444 259980 339454 260036
rect 184706 259532 184716 259588
rect 184772 259532 190120 259588
rect 339500 258804 339556 259336
rect 339490 258748 339500 258804
rect 339556 258748 339566 258804
rect 186162 258188 186172 258244
rect 186228 258188 190120 258244
rect 339500 257908 339556 258440
rect 590482 258412 590492 258468
rect 590548 258440 595672 258468
rect 590548 258412 597000 258440
rect 595560 258216 597000 258412
rect 339490 257852 339500 257908
rect 339556 257852 339566 257908
rect 339864 257516 349468 257572
rect 349524 257516 349534 257572
rect 356962 256956 356972 257012
rect 357028 256956 357308 257012
rect 357364 256956 357374 257012
rect 185938 256844 185948 256900
rect 186004 256844 190120 256900
rect 339864 256620 351372 256676
rect 351428 256620 351438 256676
rect 341282 255836 341292 255892
rect 341348 255836 359324 255892
rect 359380 255836 359390 255892
rect 339864 255724 341180 255780
rect 341236 255724 341246 255780
rect 357298 255724 357308 255780
rect 357364 255724 359492 255780
rect 359436 255668 360136 255724
rect 186050 255500 186060 255556
rect 186116 255500 190120 255556
rect 181458 255388 181468 255444
rect 181524 255388 185612 255444
rect 185668 255388 185678 255444
rect 99960 255276 178332 255332
rect 178388 255276 178398 255332
rect 339266 254828 339276 254884
rect 339332 254828 339342 254884
rect 184594 254156 184604 254212
rect 184660 254156 190120 254212
rect 339864 253932 342748 253988
rect 342804 253932 342814 253988
rect 339864 253036 346220 253092
rect 346276 253036 346286 253092
rect 187170 252812 187180 252868
rect 187236 252812 190120 252868
rect 339266 252476 339276 252532
rect 339332 252476 345772 252532
rect 345828 252476 345838 252532
rect 339864 252140 341068 252196
rect 341124 252140 341134 252196
rect 344418 252028 344428 252084
rect 344484 252028 345100 252084
rect 345156 252028 345166 252084
rect 187842 251468 187852 251524
rect 187908 251468 190120 251524
rect 339864 251244 340396 251300
rect 340452 251244 340462 251300
rect 343522 251132 343532 251188
rect 343588 251132 356188 251188
rect 356244 251132 356254 251188
rect 339266 250348 339276 250404
rect 339332 250348 339342 250404
rect 190652 249844 190708 250152
rect 359436 249844 360136 249900
rect 190642 249788 190652 249844
rect 190708 249788 190718 249844
rect 356962 249788 356972 249844
rect 357028 249788 357420 249844
rect 357476 249788 359492 249844
rect 99960 249452 178220 249508
rect 178276 249452 179004 249508
rect 179060 249452 179070 249508
rect 339864 249452 343420 249508
rect 343476 249452 343486 249508
rect 357074 249452 357084 249508
rect 357140 249452 358764 249508
rect 358820 249452 358830 249508
rect 190642 248780 190652 248836
rect 190708 248780 190718 248836
rect -960 248500 480 248696
rect 339864 248556 343084 248612
rect 343140 248556 343150 248612
rect 347890 248556 347900 248612
rect 347956 248556 349244 248612
rect 349300 248556 349310 248612
rect -960 248472 4172 248500
rect 392 248444 4172 248472
rect 4228 248444 4238 248500
rect 342402 248444 342412 248500
rect 342468 248444 349132 248500
rect 349188 248444 349198 248500
rect 342178 247772 342188 247828
rect 342244 247772 352940 247828
rect 352996 247772 353006 247828
rect 190652 247268 190708 247464
rect 190642 247212 190652 247268
rect 190708 247212 190718 247268
rect 339276 247156 339332 247688
rect 339266 247100 339276 247156
rect 339332 247100 339342 247156
rect 339388 246372 339444 246792
rect 339378 246316 339388 246372
rect 339444 246316 339454 246372
rect 190652 245476 190708 246120
rect 339864 245868 341628 245924
rect 341684 245868 341694 245924
rect 190642 245420 190652 245476
rect 190708 245420 190718 245476
rect 356626 245196 356636 245252
rect 356692 245196 357196 245252
rect 357252 245196 357262 245252
rect 595560 245028 597000 245224
rect 587122 244972 587132 245028
rect 587188 245000 597000 245028
rect 587188 244972 595672 245000
rect 190530 244748 190540 244804
rect 190596 244748 190606 244804
rect 356626 244076 356636 244132
rect 356692 244076 359492 244132
rect 359436 244020 360136 244076
rect 99960 243628 179116 243684
rect 179172 243628 179182 243684
rect 185602 243516 185612 243572
rect 185668 243516 188188 243572
rect 188244 243516 188254 243572
rect 339266 243516 339276 243572
rect 339332 243516 341068 243572
rect 341124 243516 341134 243572
rect 190652 242676 190708 243432
rect 190642 242620 190652 242676
rect 190708 242620 190718 242676
rect 188066 242060 188076 242116
rect 188132 242060 190120 242116
rect 349122 241948 349132 242004
rect 349188 241948 349356 242004
rect 349412 241948 349422 242004
rect 338594 241836 338604 241892
rect 338660 241836 339276 241892
rect 339332 241836 339342 241892
rect 343298 241836 343308 241892
rect 343364 241836 343374 241892
rect 343308 241780 343364 241836
rect 335906 241724 335916 241780
rect 335972 241724 343364 241780
rect 198034 241612 198044 241668
rect 198100 241612 335804 241668
rect 335860 241612 335870 241668
rect 337698 241612 337708 241668
rect 337764 241612 342748 241668
rect 342804 241612 342814 241668
rect 322578 241388 322588 241444
rect 322644 241388 345548 241444
rect 345604 241388 345614 241444
rect 187058 241276 187068 241332
rect 187124 241276 273868 241332
rect 273924 241276 273934 241332
rect 318546 241276 318556 241332
rect 318612 241276 359212 241332
rect 359268 241276 359278 241332
rect 187394 241164 187404 241220
rect 187460 241164 278908 241220
rect 278964 241164 278974 241220
rect 288194 241164 288204 241220
rect 288260 241164 342972 241220
rect 343028 241164 343038 241220
rect 60844 241052 126812 241108
rect 126868 241052 126878 241108
rect 190642 241052 190652 241108
rect 190708 241052 290668 241108
rect 317874 241052 317884 241108
rect 317940 241052 359660 241108
rect 359716 241052 359726 241108
rect 60844 240772 60900 241052
rect 290612 240772 290668 241052
rect 334114 240940 334124 240996
rect 334180 240940 343084 240996
rect 343140 240940 343150 240996
rect 309092 240828 339892 240884
rect 343746 240828 343756 240884
rect 343812 240828 349580 240884
rect 349636 240828 349646 240884
rect 60834 240716 60844 240772
rect 60900 240716 60910 240772
rect 74946 240716 74956 240772
rect 75012 240716 180684 240772
rect 180740 240716 180750 240772
rect 290612 240716 304892 240772
rect 304948 240716 304958 240772
rect 309092 240660 309148 240828
rect 181346 240604 181356 240660
rect 181412 240604 309148 240660
rect 309260 240716 334236 240772
rect 334292 240716 334302 240772
rect 309260 240548 309316 240716
rect 339836 240660 339892 240828
rect 342178 240716 342188 240772
rect 342244 240716 351372 240772
rect 351428 240716 351438 240772
rect 64866 240492 64876 240548
rect 64932 240492 184156 240548
rect 184212 240492 184222 240548
rect 185714 240492 185724 240548
rect 185780 240492 309316 240548
rect 311612 240604 315644 240660
rect 315700 240604 315710 240660
rect 317846 240604 317884 240660
rect 317940 240604 317950 240660
rect 318518 240604 318556 240660
rect 318612 240604 318622 240660
rect 322550 240604 322588 240660
rect 322644 240604 322654 240660
rect 323222 240604 323260 240660
rect 323316 240604 323326 240660
rect 337138 240604 337148 240660
rect 337204 240604 339780 240660
rect 339836 240604 341292 240660
rect 341348 240604 350588 240660
rect 350644 240604 350654 240660
rect 311612 240436 311668 240604
rect 339724 240548 339780 240604
rect 62850 240380 62860 240436
rect 62916 240380 190540 240436
rect 190596 240380 190606 240436
rect 197474 240380 197484 240436
rect 197540 240380 311668 240436
rect 311724 240492 336924 240548
rect 336980 240492 336990 240548
rect 338258 240492 338268 240548
rect 338324 240492 338334 240548
rect 339724 240492 346108 240548
rect 346164 240492 346174 240548
rect 311724 240324 311780 240492
rect 338268 240436 338324 240492
rect 315634 240380 315644 240436
rect 315700 240380 321076 240436
rect 66882 240268 66892 240324
rect 66948 240268 183932 240324
rect 183988 240268 183998 240324
rect 197698 240268 197708 240324
rect 197764 240268 311780 240324
rect 321020 240324 321076 240380
rect 332612 240380 338324 240436
rect 343522 240380 343532 240436
rect 343588 240380 346220 240436
rect 346276 240380 346286 240436
rect 332612 240324 332668 240380
rect 321020 240268 332668 240324
rect 336018 240268 336028 240324
rect 336084 240268 337596 240324
rect 337652 240268 337662 240324
rect 344866 240268 344876 240324
rect 344932 240268 345100 240324
rect 345156 240268 345166 240324
rect 358418 240268 358428 240324
rect 358484 240268 358988 240324
rect 359044 240268 359054 240324
rect 48514 240156 48524 240212
rect 48580 240156 67228 240212
rect 68898 240156 68908 240212
rect 68964 240156 197372 240212
rect 197428 240156 197438 240212
rect 317202 240156 317212 240212
rect 317268 240156 320180 240212
rect 320534 240156 320572 240212
rect 320628 240156 320638 240212
rect 320852 240156 359772 240212
rect 359828 240156 359838 240212
rect 67172 240100 67228 240156
rect 320124 240100 320180 240156
rect 320852 240100 320908 240156
rect 56802 240044 56812 240100
rect 56868 240044 56878 240100
rect 67172 240044 214396 240100
rect 214452 240044 214462 240100
rect 303090 240044 303100 240100
rect 303156 240044 314972 240100
rect 315028 240044 315038 240100
rect 319862 240044 319900 240100
rect 319956 240044 319966 240100
rect 320124 240044 320908 240100
rect 325826 240044 325836 240100
rect 325892 240044 358988 240100
rect 359044 240044 359054 240100
rect 56812 239988 56868 240044
rect 56812 239932 120092 239988
rect 120148 239932 120158 239988
rect 174626 239932 174636 239988
rect 174692 239932 337036 239988
rect 337092 239932 337102 239988
rect 338370 239932 338380 239988
rect 338436 239932 358764 239988
rect 358820 239932 358830 239988
rect 58818 239820 58828 239876
rect 58884 239820 115052 239876
rect 115108 239820 115118 239876
rect 182354 239820 182364 239876
rect 182420 239820 341292 239876
rect 341348 239820 341358 239876
rect 80994 239708 81004 239764
rect 81060 239708 125132 239764
rect 125188 239708 125198 239764
rect 186274 239708 186284 239764
rect 186340 239708 344988 239764
rect 345044 239708 345054 239764
rect 187282 239596 187292 239652
rect 187348 239596 341068 239652
rect 341124 239596 341134 239652
rect 182578 239484 182588 239540
rect 182644 239484 318332 239540
rect 318388 239484 318398 239540
rect 319218 239484 319228 239540
rect 319284 239484 358764 239540
rect 358820 239484 358830 239540
rect 4162 239372 4172 239428
rect 4228 239372 290668 239428
rect 304854 239372 304892 239428
rect 304948 239372 304958 239428
rect 314962 239372 314972 239428
rect 315028 239372 325836 239428
rect 325892 239372 325902 239428
rect 326060 239372 339612 239428
rect 339668 239372 339678 239428
rect 290612 239316 290668 239372
rect 184370 239260 184380 239316
rect 184436 239260 272748 239316
rect 272804 239260 272814 239316
rect 288166 239260 288204 239316
rect 288260 239260 288270 239316
rect 290612 239260 307356 239316
rect 307412 239260 307422 239316
rect 326060 239204 326116 239372
rect 314850 239148 314860 239204
rect 314916 239148 326116 239204
rect 317426 239036 317436 239092
rect 317492 239036 341180 239092
rect 341236 239036 341246 239092
rect 341058 238588 341068 238644
rect 341124 238588 345772 238644
rect 345828 238588 345838 238644
rect 347778 238588 347788 238644
rect 347844 238588 349244 238644
rect 349300 238588 349310 238644
rect 38546 238476 38556 238532
rect 38612 238476 46732 238532
rect 46788 238476 46798 238532
rect 72902 238476 72940 238532
rect 72996 238476 73006 238532
rect 76934 238476 76972 238532
rect 77028 238476 77038 238532
rect 91074 238476 91084 238532
rect 91140 238476 91150 238532
rect 95106 238476 95116 238532
rect 95172 238476 99932 238532
rect 99988 238476 99998 238532
rect 188178 238476 188188 238532
rect 188244 238476 206332 238532
rect 206388 238476 206398 238532
rect 241910 238476 241948 238532
rect 242004 238476 242014 238532
rect 242582 238476 242620 238532
rect 242676 238476 242686 238532
rect 247314 238476 247324 238532
rect 247380 238476 270732 238532
rect 270788 238476 270798 238532
rect 286290 238476 286300 238532
rect 286356 238476 294812 238532
rect 294868 238476 294878 238532
rect 321206 238476 321244 238532
rect 321300 238476 321310 238532
rect 321878 238476 321916 238532
rect 321972 238476 321982 238532
rect 91084 238420 91140 238476
rect 40226 238364 40236 238420
rect 40292 238364 52780 238420
rect 52836 238364 52846 238420
rect 91084 238364 96852 238420
rect 97122 238364 97132 238420
rect 97188 238364 106652 238420
rect 106708 238364 106718 238420
rect 243282 238364 243292 238420
rect 243348 238364 267260 238420
rect 267316 238364 267326 238420
rect 288978 238364 288988 238420
rect 289044 238364 299964 238420
rect 300020 238364 300030 238420
rect 313170 238364 313180 238420
rect 313236 238364 356748 238420
rect 356804 238364 356814 238420
rect 38434 238252 38444 238308
rect 38500 238252 50764 238308
rect 50820 238252 50830 238308
rect 93090 238252 93100 238308
rect 93156 238252 96572 238308
rect 96628 238252 96638 238308
rect 96796 238196 96852 238364
rect 97010 238252 97020 238308
rect 97076 238252 111692 238308
rect 111748 238252 111758 238308
rect 244626 238252 244636 238308
rect 244692 238252 269724 238308
rect 269780 238252 269790 238308
rect 280914 238252 280924 238308
rect 280980 238252 293244 238308
rect 293300 238252 293310 238308
rect 312498 238252 312508 238308
rect 312564 238252 354172 238308
rect 354228 238252 354238 238308
rect 359436 238196 360136 238252
rect 38322 238140 38332 238196
rect 38388 238140 48748 238196
rect 48804 238140 48814 238196
rect 87042 238140 87052 238196
rect 87108 238140 96572 238196
rect 96628 238140 96638 238196
rect 96796 238140 103516 238196
rect 103572 238140 103582 238196
rect 249330 238140 249340 238196
rect 249396 238140 273868 238196
rect 273924 238140 273934 238196
rect 278898 238140 278908 238196
rect 278964 238140 301644 238196
rect 301700 238140 301710 238196
rect 311154 238140 311164 238196
rect 311220 238140 350700 238196
rect 350756 238140 350766 238196
rect 356962 238140 356972 238196
rect 357028 238140 359492 238196
rect 85026 238028 85036 238084
rect 85092 238028 118412 238084
rect 118468 238028 118478 238084
rect 248658 238028 248668 238084
rect 248724 238028 273980 238084
rect 274036 238028 274046 238084
rect 278226 238028 278236 238084
rect 278292 238028 303996 238084
rect 304052 238028 304062 238084
rect 315858 238028 315868 238084
rect 315924 238028 352268 238084
rect 352324 238028 352334 238084
rect 40674 237916 40684 237972
rect 40740 237916 54796 237972
rect 54852 237916 54862 237972
rect 78978 237916 78988 237972
rect 79044 237916 103292 237972
rect 103348 237916 103358 237972
rect 245970 237916 245980 237972
rect 246036 237916 279020 237972
rect 279076 237916 279086 237972
rect 282258 237916 282268 237972
rect 282324 237916 303548 237972
rect 303604 237916 303614 237972
rect 314514 237916 314524 237972
rect 314580 237916 350476 237972
rect 350532 237916 350542 237972
rect 83010 237804 83020 237860
rect 83076 237804 100380 237860
rect 100436 237804 100446 237860
rect 243954 237804 243964 237860
rect 244020 237804 277228 237860
rect 277284 237804 277294 237860
rect 277554 237804 277564 237860
rect 277620 237804 305004 237860
rect 305060 237804 305070 237860
rect 311826 237804 311836 237860
rect 311892 237804 345324 237860
rect 345380 237804 345390 237860
rect 89058 237692 89068 237748
rect 89124 237692 100156 237748
rect 100212 237692 100222 237748
rect 245298 237692 245308 237748
rect 245364 237692 278908 237748
rect 278964 237692 278974 237748
rect 279570 237692 279580 237748
rect 279636 237692 308700 237748
rect 308756 237692 308766 237748
rect 310482 237692 310492 237748
rect 310548 237692 341964 237748
rect 342020 237692 342030 237748
rect 96562 237580 96572 237636
rect 96628 237580 104972 237636
rect 105028 237580 105038 237636
rect 306450 237580 306460 237636
rect 306516 237580 350924 237636
rect 350980 237580 350990 237636
rect 247986 237468 247996 237524
rect 248052 237468 269836 237524
rect 269892 237468 269902 237524
rect 308466 237468 308476 237524
rect 308532 237468 312508 237524
rect 312564 237468 312574 237524
rect 313842 237468 313852 237524
rect 313908 237468 340172 237524
rect 340228 237468 340238 237524
rect 233174 237244 233212 237300
rect 233268 237244 233278 237300
rect 235862 237244 235900 237300
rect 235956 237244 235966 237300
rect 218418 237020 218428 237076
rect 218484 237020 219996 237076
rect 220052 237020 220062 237076
rect 267474 237020 267484 237076
rect 267540 237020 268716 237076
rect 268772 237020 268782 237076
rect 269490 237020 269500 237076
rect 269556 237020 270284 237076
rect 270340 237020 270350 237076
rect 292338 237020 292348 237076
rect 292404 237020 293916 237076
rect 293972 237020 293982 237076
rect 218278 236908 218316 236964
rect 218372 236908 218382 236964
rect 228498 236908 228508 236964
rect 228564 236908 229180 236964
rect 229236 236908 229246 236964
rect 236758 236908 236796 236964
rect 236852 236908 236862 236964
rect 268566 236908 268604 236964
rect 268660 236908 268670 236964
rect 270358 236908 270396 236964
rect 270452 236908 270462 236964
rect 293766 236908 293804 236964
rect 293860 236908 293870 236964
rect 295558 236908 295596 236964
rect 295652 236908 295662 236964
rect 297714 236908 297724 236964
rect 297780 236908 298956 236964
rect 299012 236908 299022 236964
rect 299730 236908 299740 236964
rect 299796 236908 300636 236964
rect 300692 236908 300702 236964
rect 316530 236796 316540 236852
rect 316596 236796 340060 236852
rect 340116 236796 340126 236852
rect 351810 236796 351820 236852
rect 351876 236796 356636 236852
rect 356692 236796 356702 236852
rect 305106 236684 305116 236740
rect 305172 236684 358652 236740
rect 358708 236684 358718 236740
rect 260082 236572 260092 236628
rect 260148 236572 306572 236628
rect 306628 236572 306638 236628
rect 307346 236572 307356 236628
rect 307412 236572 359884 236628
rect 359940 236572 359950 236628
rect 227826 236460 227836 236516
rect 227892 236460 269388 236516
rect 269444 236460 269454 236516
rect 304434 236460 304444 236516
rect 304500 236460 357308 236516
rect 357364 236460 357374 236516
rect 251346 236348 251356 236404
rect 251412 236348 298172 236404
rect 298228 236348 298238 236404
rect 305778 236348 305788 236404
rect 305844 236348 355516 236404
rect 355572 236348 355582 236404
rect 188066 236236 188076 236292
rect 188132 236236 279692 236292
rect 279748 236236 279758 236292
rect 303762 236236 303772 236292
rect 303828 236236 352380 236292
rect 352436 236236 352446 236292
rect 46946 236124 46956 236180
rect 47012 236124 210364 236180
rect 210420 236124 210430 236180
rect 250674 236124 250684 236180
rect 250740 236124 301532 236180
rect 301588 236124 301598 236180
rect 307122 236124 307132 236180
rect 307188 236124 347228 236180
rect 347284 236124 347294 236180
rect 46162 236012 46172 236068
rect 46228 236012 273756 236068
rect 273812 236012 273822 236068
rect 307318 236012 307356 236068
rect 307412 236012 307422 236068
rect 307794 236012 307804 236068
rect 307860 236012 340396 236068
rect 340452 236012 340462 236068
rect 197586 235900 197596 235956
rect 197652 235900 359660 235956
rect 359716 235900 359726 235956
rect 70914 235116 70924 235172
rect 70980 235116 180572 235172
rect 180628 235116 180638 235172
rect 225138 235116 225148 235172
rect 225204 235116 267484 235172
rect 267540 235116 267550 235172
rect 273746 235116 273756 235172
rect 273812 235116 340172 235172
rect 340228 235116 340238 235172
rect 356738 235116 356748 235172
rect 356804 235116 358540 235172
rect 358596 235116 358606 235172
rect 223794 235004 223804 235060
rect 223860 235004 266812 235060
rect 266868 235004 266878 235060
rect 312498 235004 312508 235060
rect 312564 235004 340956 235060
rect 341012 235004 341022 235060
rect 315186 234892 315196 234948
rect 315252 234892 340732 234948
rect 340788 234892 340798 234948
rect 181010 234780 181020 234836
rect 181076 234780 330652 234836
rect 330708 234780 330718 234836
rect 179666 234668 179676 234724
rect 179732 234668 341740 234724
rect 341796 234668 341806 234724
rect -960 234388 480 234584
rect 51762 234556 51772 234612
rect 51828 234556 215068 234612
rect 215124 234556 215134 234612
rect 217074 234556 217084 234612
rect 217140 234556 269276 234612
rect 269332 234556 269342 234612
rect 311154 234556 311164 234612
rect 311220 234556 342076 234612
rect 342132 234556 342142 234612
rect 50194 234444 50204 234500
rect 50260 234444 215740 234500
rect 215796 234444 215806 234500
rect 216402 234444 216412 234500
rect 216468 234444 271068 234500
rect 271124 234444 271134 234500
rect 315186 234444 315196 234500
rect 315252 234444 356748 234500
rect 356804 234444 356814 234500
rect -960 234360 130172 234388
rect 392 234332 130172 234360
rect 130228 234332 130238 234388
rect 206322 234332 206332 234388
rect 206388 234332 267148 234388
rect 267204 234332 267214 234388
rect 289762 234332 289772 234388
rect 289828 234332 342860 234388
rect 342916 234332 342926 234388
rect 225810 234220 225820 234276
rect 225876 234220 267372 234276
rect 267428 234220 267438 234276
rect 177874 234108 177884 234164
rect 177940 234108 321692 234164
rect 321748 234108 321758 234164
rect 301746 233436 301756 233492
rect 301812 233436 341852 233492
rect 341908 233436 341918 233492
rect 188738 233100 188748 233156
rect 188804 233100 311612 233156
rect 311668 233100 311678 233156
rect 175970 232988 175980 233044
rect 176036 232988 320572 233044
rect 320628 232988 320638 233044
rect 180898 232876 180908 232932
rect 180964 232876 326172 232932
rect 326228 232876 326238 232932
rect 179442 232764 179452 232820
rect 179508 232764 336252 232820
rect 336308 232764 336318 232820
rect 22754 232652 22764 232708
rect 22820 232652 207676 232708
rect 207732 232652 207742 232708
rect 240594 232652 240604 232708
rect 240660 232652 270620 232708
rect 270676 232652 270686 232708
rect 309922 232652 309932 232708
rect 309988 232652 352492 232708
rect 352548 232652 352558 232708
rect 359436 232372 360136 232428
rect 357186 232316 357196 232372
rect 357252 232316 359492 232372
rect 595560 231924 597000 232008
rect 590706 231868 590716 231924
rect 590772 231868 597000 231924
rect 227154 231756 227164 231812
rect 227220 231756 269612 231812
rect 269668 231756 269678 231812
rect 595560 231784 597000 231868
rect 219762 231644 219772 231700
rect 219828 231644 269612 231700
rect 269668 231644 269678 231700
rect 312386 231644 312396 231700
rect 312452 231644 337372 231700
rect 337428 231644 337438 231700
rect 220434 231532 220444 231588
rect 220500 231532 274428 231588
rect 274484 231532 274494 231588
rect 311714 231532 311724 231588
rect 311780 231532 337148 231588
rect 337204 231532 337214 231588
rect 219090 231420 219100 231476
rect 219156 231420 271180 231476
rect 271236 231420 271246 231476
rect 272962 231420 272972 231476
rect 273028 231420 340284 231476
rect 340340 231420 340350 231476
rect 179106 231308 179116 231364
rect 179172 231308 305116 231364
rect 305172 231308 305182 231364
rect 311938 231308 311948 231364
rect 312004 231308 351260 231364
rect 351316 231308 351326 231364
rect 188850 231196 188860 231252
rect 188916 231196 319452 231252
rect 319508 231196 319518 231252
rect 320002 231196 320012 231252
rect 320068 231196 343420 231252
rect 343476 231196 343486 231252
rect 186274 231084 186284 231140
rect 186340 231084 328412 231140
rect 328468 231084 328478 231140
rect 329186 231084 329196 231140
rect 329252 231084 336028 231140
rect 336084 231084 336094 231140
rect 189186 230972 189196 231028
rect 189252 230972 335132 231028
rect 335188 230972 335198 231028
rect 226482 230860 226492 230916
rect 226548 230860 267596 230916
rect 267652 230860 267662 230916
rect 309810 230860 309820 230916
rect 309876 230860 341964 230916
rect 342020 230860 342030 230916
rect 311042 230188 311052 230244
rect 311108 230188 357980 230244
rect 358036 230188 358764 230244
rect 358820 230188 358830 230244
rect 309138 230076 309148 230132
rect 309204 230076 340508 230132
rect 340564 230076 340574 230132
rect 182690 229852 182700 229908
rect 182756 229852 314972 229908
rect 315028 229852 315038 229908
rect 189074 229740 189084 229796
rect 189140 229740 325052 229796
rect 325108 229740 325118 229796
rect 181122 229628 181132 229684
rect 181188 229628 332892 229684
rect 332948 229628 332958 229684
rect 40226 229516 40236 229572
rect 40292 229516 212380 229572
rect 212436 229516 212446 229572
rect 309922 229516 309932 229572
rect 309988 229516 338940 229572
rect 338996 229516 339006 229572
rect 13234 229404 13244 229460
rect 13300 229404 207004 229460
rect 207060 229404 207070 229460
rect 258066 229404 258076 229460
rect 258132 229404 306796 229460
rect 306852 229404 306862 229460
rect 310146 229404 310156 229460
rect 310212 229404 345548 229460
rect 345604 229404 345614 229460
rect 20850 229292 20860 229348
rect 20916 229292 339836 229348
rect 339892 229292 339902 229348
rect 237234 228396 237244 228452
rect 237300 228396 270732 228452
rect 270788 228396 270798 228452
rect 302418 228396 302428 228452
rect 302484 228396 357084 228452
rect 357140 228396 357150 228452
rect 228498 228284 228508 228340
rect 228564 228284 271292 228340
rect 271348 228284 271358 228340
rect 222450 228172 222460 228228
rect 222516 228172 274092 228228
rect 274148 228172 274158 228228
rect 221106 228060 221116 228116
rect 221172 228060 274540 228116
rect 274596 228060 274606 228116
rect 186162 227948 186172 228004
rect 186228 227948 322812 228004
rect 322868 227948 322878 228004
rect 182802 227836 182812 227892
rect 182868 227836 329532 227892
rect 329588 227836 329598 227892
rect 181234 227724 181244 227780
rect 181300 227724 340732 227780
rect 340788 227724 340798 227780
rect 30370 227612 30380 227668
rect 30436 227612 208348 227668
rect 208404 227612 208414 227668
rect 221778 227612 221788 227668
rect 221844 227612 275772 227668
rect 275828 227612 275838 227668
rect 279794 227612 279804 227668
rect 279860 227612 354620 227668
rect 354676 227612 354686 227668
rect 237906 227500 237916 227556
rect 237972 227500 270620 227556
rect 270676 227500 270686 227556
rect 359436 226548 360136 226604
rect 259410 226492 259420 226548
rect 259476 226492 304892 226548
rect 304948 226492 304958 226548
rect 357074 226492 357084 226548
rect 357140 226492 359492 226548
rect 289874 226380 289884 226436
rect 289940 226380 338380 226436
rect 338436 226380 338446 226436
rect 286626 226268 286636 226324
rect 286692 226268 337260 226324
rect 337316 226268 337326 226324
rect 283154 226156 283164 226212
rect 283220 226156 338716 226212
rect 338772 226156 338782 226212
rect 286402 226044 286412 226100
rect 286468 226044 349468 226100
rect 349524 226044 349534 226100
rect 286850 225932 286860 225988
rect 286916 225932 351372 225988
rect 351428 225932 351438 225988
rect 239250 225036 239260 225092
rect 239316 225036 270956 225092
rect 271012 225036 271022 225092
rect 224466 224924 224476 224980
rect 224532 224924 274316 224980
rect 274372 224924 274382 224980
rect 184482 224812 184492 224868
rect 184548 224812 327292 224868
rect 327348 224812 327358 224868
rect 178882 224700 178892 224756
rect 178948 224700 321804 224756
rect 321860 224700 321870 224756
rect 177986 224588 177996 224644
rect 178052 224588 337372 224644
rect 337428 224588 337438 224644
rect 48626 224476 48636 224532
rect 48692 224476 213724 224532
rect 213780 224476 213790 224532
rect 257394 224476 257404 224532
rect 257460 224476 310044 224532
rect 310100 224476 310110 224532
rect 38546 224364 38556 224420
rect 38612 224364 209692 224420
rect 209748 224364 209758 224420
rect 223122 224364 223132 224420
rect 223188 224364 275884 224420
rect 275940 224364 275950 224420
rect 276322 224364 276332 224420
rect 276388 224364 336588 224420
rect 336644 224364 336654 224420
rect 51986 224252 51996 224308
rect 52052 224252 235228 224308
rect 235284 224252 235294 224308
rect 241266 224252 241276 224308
rect 241332 224252 275660 224308
rect 275716 224252 275726 224308
rect 278114 224252 278124 224308
rect 278180 224252 343756 224308
rect 343812 224252 343822 224308
rect 239922 224140 239932 224196
rect 239988 224140 269500 224196
rect 269556 224140 269566 224196
rect 253362 223244 253372 223300
rect 253428 223244 306572 223300
rect 306628 223244 306638 223300
rect 186386 223132 186396 223188
rect 186452 223132 338492 223188
rect 338548 223132 338558 223188
rect 179554 223020 179564 223076
rect 179620 223020 331772 223076
rect 331828 223020 331838 223076
rect 178994 222908 179004 222964
rect 179060 222908 331996 222964
rect 332052 222908 332062 222964
rect 37986 222796 37996 222852
rect 38052 222796 209020 222852
rect 209076 222796 209086 222852
rect 279906 222796 279916 222852
rect 279972 222796 336812 222852
rect 336868 222796 336878 222852
rect 39890 222684 39900 222740
rect 39956 222684 230524 222740
rect 230580 222684 230590 222740
rect 283042 222684 283052 222740
rect 283108 222684 341404 222740
rect 341460 222684 341470 222740
rect 26562 222572 26572 222628
rect 26628 222572 341628 222628
rect 341684 222572 341694 222628
rect 256050 221340 256060 221396
rect 256116 221340 303436 221396
rect 303492 221340 303502 221396
rect 255378 221228 255388 221284
rect 255444 221228 303212 221284
rect 303268 221228 303278 221284
rect 187730 221116 187740 221172
rect 187796 221116 274092 221172
rect 274148 221116 274158 221172
rect 176082 221004 176092 221060
rect 176148 221004 317212 221060
rect 317268 221004 317278 221060
rect 176306 220892 176316 220948
rect 176372 220892 339612 220948
rect 339668 220892 339678 220948
rect 359436 220724 360136 220780
rect 356850 220668 356860 220724
rect 356916 220668 359492 220724
rect -960 220276 480 220472
rect -960 220248 118412 220276
rect 392 220220 118412 220248
rect 118468 220220 118478 220276
rect 280354 219884 280364 219940
rect 280420 219884 337148 219940
rect 337204 219884 337214 219940
rect 181234 219772 181244 219828
rect 181300 219772 272524 219828
rect 272580 219772 272590 219828
rect 280018 219772 280028 219828
rect 280084 219772 338604 219828
rect 338660 219772 338670 219828
rect 177874 219660 177884 219716
rect 177940 219660 272860 219716
rect 272916 219660 272926 219716
rect 278002 219660 278012 219716
rect 278068 219660 338828 219716
rect 338884 219660 338894 219716
rect 199490 219548 199500 219604
rect 199556 219548 310268 219604
rect 310324 219548 310334 219604
rect 184370 219436 184380 219492
rect 184436 219436 316092 219492
rect 316148 219436 316158 219492
rect 183026 219324 183036 219380
rect 183092 219324 334012 219380
rect 334068 219324 334078 219380
rect 38434 219212 38444 219268
rect 38500 219212 211036 219268
rect 211092 219212 211102 219268
rect 276434 219212 276444 219268
rect 276500 219212 342188 219268
rect 342244 219212 342254 219268
rect 595560 218596 597000 218792
rect 577042 218540 577052 218596
rect 577108 218568 597000 218596
rect 577108 218540 595672 218568
rect 266130 218316 266140 218372
rect 266196 218316 303660 218372
rect 303716 218316 303726 218372
rect 264786 218204 264796 218260
rect 264852 218204 307020 218260
rect 307076 218204 307086 218260
rect 186834 218092 186844 218148
rect 186900 218092 271068 218148
rect 271124 218092 271134 218148
rect 186946 217980 186956 218036
rect 187012 217980 275884 218036
rect 275940 217980 275950 218036
rect 184258 217868 184268 217924
rect 184324 217868 312732 217924
rect 312788 217868 312798 217924
rect 176194 217756 176204 217812
rect 176260 217756 313852 217812
rect 313908 217756 313918 217812
rect 4274 217644 4284 217700
rect 4340 217644 138572 217700
rect 138628 217644 138638 217700
rect 154914 217644 154924 217700
rect 154980 217644 172172 217700
rect 172228 217644 172238 217700
rect 182914 217644 182924 217700
rect 182980 217644 323932 217700
rect 323988 217644 323998 217700
rect 51874 217532 51884 217588
rect 51940 217532 213052 217588
rect 213108 217532 213118 217588
rect 264114 217532 264124 217588
rect 264180 217532 306796 217588
rect 306852 217532 306862 217588
rect 266802 217420 266812 217476
rect 266868 217420 303884 217476
rect 303940 217420 303950 217476
rect 187618 216524 187628 216580
rect 187684 216524 270956 216580
rect 271012 216524 271022 216580
rect 187506 216412 187516 216468
rect 187572 216412 275772 216468
rect 275828 216412 275838 216468
rect 289986 216412 289996 216468
rect 290052 216412 339276 216468
rect 339332 216412 339342 216468
rect 199602 216300 199612 216356
rect 199668 216300 290220 216356
rect 290276 216300 290286 216356
rect 199714 216188 199724 216244
rect 199780 216188 307468 216244
rect 307524 216188 307534 216244
rect 190866 216076 190876 216132
rect 190932 216076 359660 216132
rect 359716 216076 359726 216132
rect 50306 215964 50316 216020
rect 50372 215964 234556 216020
rect 234612 215964 234622 216020
rect 252690 215964 252700 216020
rect 252756 215964 303324 216020
rect 303380 215964 303390 216020
rect 41122 215852 41132 215908
rect 41188 215852 233884 215908
rect 233940 215852 233950 215908
rect 274642 215852 274652 215908
rect 274708 215852 343532 215908
rect 343588 215852 343598 215908
rect 254706 214956 254716 215012
rect 254772 214956 296492 215012
rect 296548 214956 296558 215012
rect 359436 214900 360136 214956
rect 263442 214844 263452 214900
rect 263508 214844 307132 214900
rect 307188 214844 307198 214900
rect 349412 214844 357308 214900
rect 357364 214844 359492 214900
rect 182914 214732 182924 214788
rect 182980 214732 272188 214788
rect 272244 214732 272254 214788
rect 199378 214620 199388 214676
rect 199444 214620 310940 214676
rect 310996 214620 311006 214676
rect 194226 214508 194236 214564
rect 194292 214508 346556 214564
rect 346612 214508 346622 214564
rect 38322 214396 38332 214452
rect 38388 214396 231196 214452
rect 231252 214396 231262 214452
rect 262770 214396 262780 214452
rect 262836 214396 306684 214452
rect 306740 214396 306750 214452
rect 34962 214284 34972 214340
rect 35028 214284 231868 214340
rect 231924 214284 231934 214340
rect 262098 214284 262108 214340
rect 262164 214284 306908 214340
rect 306964 214284 306974 214340
rect 349412 214228 349468 214844
rect 32274 214172 32284 214228
rect 32340 214172 229852 214228
rect 229908 214172 229918 214228
rect 252018 214172 252028 214228
rect 252084 214172 308252 214228
rect 308308 214172 308318 214228
rect 321794 214172 321804 214228
rect 321860 214172 349468 214228
rect 261426 214060 261436 214116
rect 261492 214060 298172 214116
rect 298228 214060 298238 214116
rect 246642 213276 246652 213332
rect 246708 213276 270508 213332
rect 270564 213276 270574 213332
rect 184482 213164 184492 213220
rect 184548 213164 272412 213220
rect 272468 213164 272478 213220
rect 265458 213052 265468 213108
rect 265524 213052 303100 213108
rect 303156 213052 303166 213108
rect 179666 212940 179676 212996
rect 179732 212940 272972 212996
rect 273028 212940 273038 212996
rect 174514 212828 174524 212884
rect 174580 212828 272300 212884
rect 272356 212828 272366 212884
rect 4610 212716 4620 212772
rect 4676 212716 120092 212772
rect 120148 212716 120158 212772
rect 174402 212716 174412 212772
rect 174468 212716 273420 212772
rect 273476 212716 273486 212772
rect 4386 212604 4396 212660
rect 4452 212604 167132 212660
rect 167188 212604 167198 212660
rect 189298 212604 189308 212660
rect 189364 212604 345100 212660
rect 345156 212604 345166 212660
rect 39666 212492 39676 212548
rect 39732 212492 232540 212548
rect 232596 212492 232606 212548
rect 256722 212492 256732 212548
rect 256788 212492 299852 212548
rect 299908 212492 299918 212548
rect 49634 211708 49644 211764
rect 49700 211708 273980 211764
rect 274036 211708 274046 211764
rect 254034 211596 254044 211652
rect 254100 211596 293132 211652
rect 293188 211596 293198 211652
rect 260754 211484 260764 211540
rect 260820 211484 307244 211540
rect 307300 211484 307310 211540
rect 258738 211372 258748 211428
rect 258804 211372 308252 211428
rect 308308 211372 308318 211428
rect 190082 211260 190092 211316
rect 190148 211260 269500 211316
rect 269556 211260 269566 211316
rect 272374 211260 272412 211316
rect 272468 211260 272478 211316
rect 185714 211148 185724 211204
rect 185780 211148 272636 211204
rect 272692 211148 272702 211204
rect 4498 211036 4508 211092
rect 4564 211036 113372 211092
rect 113428 211036 113438 211092
rect 177986 211036 177996 211092
rect 178052 211036 272412 211092
rect 272468 211036 272478 211092
rect 273522 211036 273532 211092
rect 273588 211036 310380 211092
rect 310436 211036 310446 211092
rect 4162 210924 4172 210980
rect 4228 210924 121772 210980
rect 121828 210924 121838 210980
rect 272178 210924 272188 210980
rect 272244 210924 272300 210980
rect 272356 210924 272366 210980
rect 272850 210924 272860 210980
rect 272916 210924 310604 210980
rect 310660 210924 310670 210980
rect 33506 210812 33516 210868
rect 33572 210812 211708 210868
rect 211764 210812 211774 210868
rect 272178 210812 272188 210868
rect 272244 210812 355516 210868
rect 355572 210812 355582 210868
rect 250002 210700 250012 210756
rect 250068 210700 277340 210756
rect 277396 210700 277406 210756
rect 174290 210476 174300 210532
rect 174356 210476 273196 210532
rect 273252 210476 273262 210532
rect 49522 210028 49532 210084
rect 49588 210028 274652 210084
rect 274708 210028 274718 210084
rect 238578 209916 238588 209972
rect 238644 209916 272188 209972
rect 272244 209916 272254 209972
rect 272598 209916 272636 209972
rect 272692 209916 272702 209972
rect 349682 209916 349692 209972
rect 349748 209916 351036 209972
rect 351092 209916 351102 209972
rect 190418 209804 190428 209860
rect 190484 209804 272748 209860
rect 272804 209804 272814 209860
rect 185826 209692 185836 209748
rect 185892 209692 273084 209748
rect 273140 209692 273150 209748
rect 174626 209580 174636 209636
rect 174692 209580 272188 209636
rect 272244 209580 272254 209636
rect 184594 209468 184604 209524
rect 184660 209468 343980 209524
rect 344036 209468 344046 209524
rect 181346 209356 181356 209412
rect 181412 209356 349804 209412
rect 349860 209356 349870 209412
rect 359846 209244 359884 209300
rect 359940 209244 359950 209300
rect 272486 209132 272524 209188
rect 272580 209132 272590 209188
rect 331986 209132 331996 209188
rect 332052 209132 357420 209188
rect 357476 209132 359492 209188
rect 359436 209076 360136 209132
rect 4162 208684 4172 208740
rect 4228 208684 269164 208740
rect 269220 208684 269230 208740
rect 269864 207004 272300 207060
rect 272356 207004 272366 207060
rect 392 206360 4172 206388
rect -960 206332 4172 206360
rect 4228 206332 4238 206388
rect -960 206136 480 206332
rect 352772 205996 359884 206052
rect 359940 205996 359950 206052
rect 273074 205884 273084 205940
rect 273140 205884 350812 205940
rect 350868 205884 350878 205940
rect 352772 205828 352828 205996
rect 273298 205772 273308 205828
rect 273364 205772 352828 205828
rect 359846 205772 359884 205828
rect 359940 205772 359950 205828
rect 595560 205380 597000 205576
rect 560242 205324 560252 205380
rect 560308 205352 597000 205380
rect 560308 205324 595672 205352
rect 355842 204988 355852 205044
rect 355908 204988 356188 205044
rect 356244 204988 356254 205044
rect 269864 204092 272188 204148
rect 272244 204092 272254 204148
rect 305106 204092 305116 204148
rect 305172 204092 356748 204148
rect 356804 204092 356814 204148
rect 356738 203308 356748 203364
rect 356804 203308 359492 203364
rect 359436 203252 360136 203308
rect 342934 201516 342972 201572
rect 343028 201516 343038 201572
rect 269864 201180 273420 201236
rect 273476 201180 273486 201236
rect 269864 198268 272860 198324
rect 272916 198268 272926 198324
rect 345772 198268 346276 198324
rect 345772 198212 345828 198268
rect 346220 198212 346276 198268
rect 339378 198156 339388 198212
rect 339444 198156 345828 198212
rect 345958 198156 345996 198212
rect 346052 198156 346062 198212
rect 346220 198156 349468 198212
rect 349412 198100 349468 198156
rect 345202 198044 345212 198100
rect 345268 198044 347900 198100
rect 347956 198044 347966 198100
rect 349412 198044 359884 198100
rect 359940 198044 359950 198100
rect 336690 197932 336700 197988
rect 336756 197932 358988 197988
rect 359044 197932 359054 197988
rect 317202 197820 317212 197876
rect 317268 197820 339500 197876
rect 339556 197820 339566 197876
rect 317314 197708 317324 197764
rect 317380 197708 341516 197764
rect 341572 197708 341582 197764
rect 315298 197596 315308 197652
rect 315364 197596 340060 197652
rect 340116 197596 340126 197652
rect 344978 197484 344988 197540
rect 345044 197484 359324 197540
rect 359380 197484 359492 197540
rect 359436 197428 360136 197484
rect 270274 197372 270284 197428
rect 270340 197372 350700 197428
rect 350756 197372 350766 197428
rect 338146 197260 338156 197316
rect 338212 197260 351260 197316
rect 351316 197260 351326 197316
rect 276210 197148 276220 197204
rect 276276 197148 352268 197204
rect 352324 197148 352334 197204
rect 339602 197036 339612 197092
rect 339668 197036 356076 197092
rect 356132 197036 356142 197092
rect 345650 196700 345660 196756
rect 345716 196700 349468 196756
rect 349412 196644 349468 196700
rect 345510 196588 345548 196644
rect 345604 196588 345614 196644
rect 349412 196588 352604 196644
rect 352660 196588 352670 196644
rect 341618 196476 341628 196532
rect 341684 196476 344596 196532
rect 344978 196476 344988 196532
rect 345044 196476 347788 196532
rect 347844 196476 347854 196532
rect 343186 196364 343196 196420
rect 343252 196364 343262 196420
rect 344204 196364 344316 196420
rect 344372 196364 344382 196420
rect 343196 195860 343252 196364
rect 344204 196196 344260 196364
rect 344194 196140 344204 196196
rect 344260 196140 344270 196196
rect 344540 196084 344596 196476
rect 344754 196364 344764 196420
rect 344820 196364 344830 196420
rect 345650 196364 345660 196420
rect 345716 196364 345726 196420
rect 345874 196364 345884 196420
rect 345940 196364 346556 196420
rect 346612 196364 346622 196420
rect 344764 196196 344820 196364
rect 345660 196308 345716 196364
rect 345660 196252 349580 196308
rect 349636 196252 349646 196308
rect 344764 196140 359772 196196
rect 359828 196140 359838 196196
rect 344540 196028 356188 196084
rect 356244 196028 356254 196084
rect 345538 195916 345548 195972
rect 345604 195916 354172 195972
rect 354228 195916 354238 195972
rect 343196 195804 354508 195860
rect 354564 195804 354574 195860
rect 344194 195692 344204 195748
rect 344260 195692 357868 195748
rect 357924 195692 357934 195748
rect 269864 195356 272972 195412
rect 273028 195356 273038 195412
rect 345090 194908 345100 194964
rect 345156 194908 346444 194964
rect 346500 194908 346510 194964
rect 345762 194796 345772 194852
rect 345828 194796 346948 194852
rect 313394 194684 313404 194740
rect 313460 194684 336028 194740
rect 336084 194684 336094 194740
rect 346892 194628 346948 194796
rect 346892 194600 351036 194628
rect 346920 194572 351036 194600
rect 351092 194572 351102 194628
rect 349570 193228 349580 193284
rect 349636 193228 350924 193284
rect 350980 193228 350990 193284
rect 269864 192444 272748 192500
rect 272804 192444 272814 192500
rect 346434 192444 346444 192500
rect 346500 192444 346510 192500
rect -960 192052 480 192248
rect -960 192024 14252 192052
rect 392 191996 14252 192024
rect 14308 191996 14318 192052
rect 346444 191912 346500 192444
rect 595560 192164 597000 192360
rect 590818 192108 590828 192164
rect 590884 192136 597000 192164
rect 590884 192108 595672 192136
rect 351026 191772 351036 191828
rect 351092 191772 359492 191828
rect 351138 191660 351148 191716
rect 351204 191660 352716 191716
rect 352772 191660 352782 191716
rect 359436 191660 359492 191772
rect 359436 191604 359772 191660
rect 359828 191604 360136 191660
rect 351250 191548 351260 191604
rect 351316 191548 352604 191604
rect 352660 191548 352670 191604
rect 346892 189756 350476 189812
rect 350532 189756 350812 189812
rect 350868 189756 350878 189812
rect 269864 189532 272524 189588
rect 272580 189532 272590 189588
rect 346892 189224 346948 189756
rect 350802 188076 350812 188132
rect 350868 188076 351820 188132
rect 351876 188076 351886 188132
rect 269864 186620 273196 186676
rect 273252 186620 273262 186676
rect 346920 186508 350812 186564
rect 350868 186508 350878 186564
rect 359874 186172 359884 186228
rect 359940 186172 359950 186228
rect 359884 186004 359940 186172
rect 359874 185948 359884 186004
rect 359940 185948 359950 186004
rect 356178 185836 356188 185892
rect 356244 185836 359492 185892
rect 359436 185780 360136 185836
rect 346920 183820 356972 183876
rect 357028 183820 358652 183876
rect 358708 183820 358718 183876
rect 269864 183708 273084 183764
rect 273140 183708 273150 183764
rect 356738 181356 356748 181412
rect 356804 181356 359772 181412
rect 359828 181356 359838 181412
rect 346920 181132 356972 181188
rect 357028 181132 357196 181188
rect 357252 181132 357262 181188
rect 269864 180796 272748 180852
rect 272804 180796 272814 180852
rect 359436 179956 360136 180012
rect 357746 179900 357756 179956
rect 357812 179900 359492 179956
rect 595560 178948 597000 179144
rect 570322 178892 570332 178948
rect 570388 178920 597000 178948
rect 570388 178892 595672 178920
rect 346920 178444 357084 178500
rect 357140 178444 357150 178500
rect -960 178052 480 178136
rect -960 177996 4508 178052
rect 4564 177996 4574 178052
rect 350690 177996 350700 178052
rect 350756 177996 359772 178052
rect 359828 177996 359838 178052
rect -960 177912 480 177996
rect 269864 177884 272636 177940
rect 272692 177884 272702 177940
rect 346920 175756 356972 175812
rect 357028 175756 357038 175812
rect 346546 175420 346556 175476
rect 346612 175420 590716 175476
rect 590772 175420 590782 175476
rect 356962 175308 356972 175364
rect 357028 175308 361228 175364
rect 361284 175308 361294 175364
rect 361442 175308 361452 175364
rect 361508 175308 590492 175364
rect 590548 175308 590558 175364
rect 354050 175196 354060 175252
rect 354116 175196 369180 175252
rect 369236 175196 369246 175252
rect 375190 175196 375228 175252
rect 375284 175196 375294 175252
rect 352706 175084 352716 175140
rect 352772 175084 399420 175140
rect 399476 175084 399486 175140
rect 269864 174972 272524 175028
rect 272580 174972 272590 175028
rect 358390 174636 358428 174692
rect 358484 174636 358494 174692
rect 417526 174636 417564 174692
rect 417620 174636 417630 174692
rect 361666 174524 361676 174580
rect 361732 174524 520380 174580
rect 520436 174524 520446 174580
rect 362114 174412 362124 174468
rect 362180 174412 465948 174468
rect 466004 174412 466014 174468
rect 354162 174300 354172 174356
rect 354228 174300 453852 174356
rect 453908 174300 453918 174356
rect 349010 174188 349020 174244
rect 349076 174188 393372 174244
rect 393428 174188 393438 174244
rect 359090 174076 359100 174132
rect 359156 174076 489132 174132
rect 489188 174076 489198 174132
rect 359426 173964 359436 174020
rect 359492 173964 495852 174020
rect 495908 173964 495918 174020
rect 359426 173852 359436 173908
rect 359492 173852 497196 173908
rect 497252 173852 497262 173908
rect 352146 173628 352156 173684
rect 352212 173628 387324 173684
rect 387380 173628 387390 173684
rect 355170 173516 355180 173572
rect 355236 173516 590604 173572
rect 590660 173516 590670 173572
rect 346920 173068 357308 173124
rect 357364 173068 361340 173124
rect 361396 173068 361406 173124
rect 355842 172956 355852 173012
rect 355908 172956 363132 173012
rect 363188 172956 363198 173012
rect 538514 172956 538524 173012
rect 538580 172956 549556 173012
rect 550610 172956 550620 173012
rect 550676 172956 559468 173012
rect 559524 172956 559534 173012
rect 561092 172956 562828 173012
rect 562884 172956 562894 173012
rect 355394 172844 355404 172900
rect 355460 172844 447804 172900
rect 447860 172844 447870 172900
rect 544562 172844 544572 172900
rect 544628 172844 549388 172900
rect 350354 172732 350364 172788
rect 350420 172732 435708 172788
rect 435764 172732 435774 172788
rect 549332 172676 549388 172844
rect 549500 172788 549556 172956
rect 561092 172900 561148 172956
rect 556658 172844 556668 172900
rect 556724 172844 561148 172900
rect 549500 172732 559692 172788
rect 559748 172732 559758 172788
rect 348786 172620 348796 172676
rect 348852 172620 423612 172676
rect 423668 172620 423678 172676
rect 549332 172620 559580 172676
rect 559636 172620 559646 172676
rect 359874 172508 359884 172564
rect 359940 172508 429660 172564
rect 429716 172508 429726 172564
rect 347106 172396 347116 172452
rect 347172 172396 405468 172452
rect 405524 172396 405534 172452
rect 355618 172284 355628 172340
rect 355684 172284 381276 172340
rect 381332 172284 381342 172340
rect 469522 172284 469532 172340
rect 469588 172284 559020 172340
rect 559076 172284 559086 172340
rect 360322 172172 360332 172228
rect 360388 172172 559468 172228
rect 559524 172172 559534 172228
rect 269864 172060 272412 172116
rect 272468 172060 272478 172116
rect 360546 172060 360556 172116
rect 360612 172060 490140 172116
rect 490196 172060 490206 172116
rect 348562 171276 348572 171332
rect 348628 171276 532476 171332
rect 532532 171276 532542 171332
rect 358530 171164 358540 171220
rect 358596 171164 484092 171220
rect 484148 171164 484158 171220
rect 346994 171052 347004 171108
rect 347060 171052 471996 171108
rect 472052 171052 472062 171108
rect 352034 170940 352044 170996
rect 352100 170940 459900 170996
rect 459956 170940 459966 170996
rect 353714 170828 353724 170884
rect 353780 170828 441756 170884
rect 441812 170828 441822 170884
rect 355954 170716 355964 170772
rect 356020 170716 457772 170772
rect 457828 170716 457838 170772
rect 358866 170604 358876 170660
rect 358932 170604 486444 170660
rect 486500 170604 486510 170660
rect 359090 170492 359100 170548
rect 359156 170492 494508 170548
rect 494564 170492 494574 170548
rect 346920 170380 357420 170436
rect 357476 170380 420812 170436
rect 420868 170380 420878 170436
rect 351922 169596 351932 169652
rect 351988 169596 514332 169652
rect 514388 169596 514398 169652
rect 350242 169484 350252 169540
rect 350308 169484 496188 169540
rect 496244 169484 496254 169540
rect 348674 169372 348684 169428
rect 348740 169372 478044 169428
rect 478100 169372 478110 169428
rect 355842 169260 355852 169316
rect 355908 169260 457884 169316
rect 457940 169260 457950 169316
rect 467842 169260 467852 169316
rect 467908 169260 587132 169316
rect 587188 169260 587198 169316
rect 269864 169148 274092 169204
rect 274148 169148 274158 169204
rect 358754 169148 358764 169204
rect 358820 169148 483756 169204
rect 483812 169148 483822 169204
rect 355506 169036 355516 169092
rect 355572 169036 516012 169092
rect 516068 169036 516078 169092
rect 352370 168924 352380 168980
rect 352436 168924 559804 168980
rect 559860 168924 559870 168980
rect 354050 168812 354060 168868
rect 354116 168812 563164 168868
rect 563220 168812 563230 168868
rect 348898 168700 348908 168756
rect 348964 168700 411516 168756
rect 411572 168700 411582 168756
rect 354386 167916 354396 167972
rect 354452 167916 590828 167972
rect 590884 167916 590894 167972
rect 346994 167804 347004 167860
rect 347060 167804 526428 167860
rect 526484 167804 526494 167860
rect 346892 167412 346948 167720
rect 355282 167692 355292 167748
rect 355348 167692 508284 167748
rect 508340 167692 508350 167748
rect 353602 167580 353612 167636
rect 353668 167580 502236 167636
rect 502292 167580 502302 167636
rect 361218 167468 361228 167524
rect 361284 167468 423164 167524
rect 423220 167468 423230 167524
rect 346892 167356 356748 167412
rect 356804 167356 420924 167412
rect 420980 167356 420990 167412
rect 350466 167244 350476 167300
rect 350532 167244 562828 167300
rect 562884 167244 562894 167300
rect 349412 167132 559916 167188
rect 559972 167132 559982 167188
rect 349412 167076 349468 167132
rect 346658 167020 346668 167076
rect 346724 167020 349468 167076
rect 357634 166348 357644 166404
rect 357700 166348 498540 166404
rect 498596 166348 498606 166404
rect 269864 166236 275884 166292
rect 275940 166236 275950 166292
rect 356850 166236 356860 166292
rect 356916 166236 357532 166292
rect 357588 166236 357598 166292
rect 361330 165788 361340 165844
rect 361396 165788 422940 165844
rect 422996 165788 423006 165844
rect 358530 165676 358540 165732
rect 358596 165676 482412 165732
rect 482468 165676 482478 165732
rect 595560 165704 597000 165928
rect 352258 165564 352268 165620
rect 352324 165564 563052 165620
rect 563108 165564 563118 165620
rect 359650 165452 359660 165508
rect 359716 165452 590604 165508
rect 590660 165452 590670 165508
rect 346920 165004 349692 165060
rect 349748 165004 349758 165060
rect 357074 164892 357084 164948
rect 357140 164892 477036 164948
rect 477092 164892 477102 164948
rect 357298 164780 357308 164836
rect 357364 164780 478380 164836
rect 478436 164780 478446 164836
rect 357522 164668 357532 164724
rect 357588 164668 485100 164724
rect 485156 164668 485166 164724
rect 356962 164556 356972 164612
rect 357028 164556 357532 164612
rect 357588 164556 357598 164612
rect 468962 164332 468972 164388
rect 469028 164332 565292 164388
rect 565348 164332 565358 164388
rect 350690 164220 350700 164276
rect 350756 164220 510636 164276
rect 510692 164220 510702 164276
rect 352258 164108 352268 164164
rect 352324 164108 524076 164164
rect 524132 164108 524142 164164
rect 392 164024 4172 164052
rect -960 163996 4172 164024
rect 4228 163996 4238 164052
rect 355618 163996 355628 164052
rect 355684 163996 563388 164052
rect 563444 163996 563454 164052
rect -960 163800 480 163996
rect 346434 163884 346444 163940
rect 346500 163884 559692 163940
rect 559748 163884 559758 163940
rect 346770 163772 346780 163828
rect 346836 163772 562940 163828
rect 562996 163772 563006 163828
rect 269864 163324 271068 163380
rect 271124 163324 271134 163380
rect 421586 163212 421596 163268
rect 421652 163212 474348 163268
rect 474404 163212 474414 163268
rect 356962 163100 356972 163156
rect 357028 163100 479724 163156
rect 479780 163100 479790 163156
rect 357746 162988 357756 163044
rect 357812 162988 499884 163044
rect 499940 162988 499950 163044
rect 358642 162876 358652 162932
rect 358708 162876 421596 162932
rect 421652 162876 421662 162932
rect 361666 162540 361676 162596
rect 361732 162540 421708 162596
rect 421764 162540 421774 162596
rect 352482 162428 352492 162484
rect 352548 162428 457996 162484
rect 458052 162428 458062 162484
rect 466274 162428 466284 162484
rect 466340 162428 560252 162484
rect 560308 162428 560318 162484
rect 346920 162316 350588 162372
rect 350644 162316 350654 162372
rect 359314 162316 359324 162372
rect 359380 162316 487788 162372
rect 487844 162316 487854 162372
rect 350354 162204 350364 162260
rect 350420 162204 563276 162260
rect 563332 162204 563342 162260
rect 293010 162092 293020 162148
rect 293076 162092 560364 162148
rect 560420 162092 560430 162148
rect 298386 161980 298396 162036
rect 298452 161980 564508 162036
rect 564564 161980 564574 162036
rect 290322 161868 290332 161924
rect 290388 161868 546588 161924
rect 546644 161868 546654 161924
rect 270386 161756 270396 161812
rect 270452 161756 511980 161812
rect 512036 161756 512046 161812
rect 290612 160748 314188 160804
rect 290612 160692 290668 160748
rect 314132 160692 314188 160748
rect 274866 160636 274876 160692
rect 274932 160636 290668 160692
rect 313366 160636 313404 160692
rect 313460 160636 313470 160692
rect 314132 160636 521388 160692
rect 521444 160636 521454 160692
rect 275538 160524 275548 160580
rect 275604 160524 522732 160580
rect 522788 160524 522798 160580
rect 269864 160412 272300 160468
rect 272356 160412 272366 160468
rect 301074 160412 301084 160468
rect 301140 160412 566188 160468
rect 566244 160412 566254 160468
rect 274194 160300 274204 160356
rect 274260 160300 520044 160356
rect 520100 160300 520110 160356
rect 310370 160188 310380 160244
rect 310436 160188 518700 160244
rect 518756 160188 518766 160244
rect 314850 160076 314860 160132
rect 314916 160076 314972 160132
rect 315028 160076 315038 160132
rect 317398 160076 317436 160132
rect 317492 160076 317502 160132
rect 329074 160076 329084 160132
rect 329140 160076 337708 160132
rect 344754 160076 344764 160132
rect 344820 160076 349580 160132
rect 349636 160076 350700 160132
rect 350756 160076 350766 160132
rect 337652 160020 337708 160076
rect 337652 159964 347900 160020
rect 347956 159964 347966 160020
rect 310594 159852 310604 159908
rect 310660 159852 517356 159908
rect 517412 159852 517422 159908
rect 343186 159740 343196 159796
rect 343252 159740 346220 159796
rect 346276 159740 346286 159796
rect 340050 159516 340060 159572
rect 340116 159516 351372 159572
rect 351428 159516 352492 159572
rect 352548 159516 352558 159572
rect 286962 159404 286972 159460
rect 287028 159404 524188 159460
rect 524244 159404 524254 159460
rect 270834 159292 270844 159348
rect 270900 159292 513324 159348
rect 513380 159292 513390 159348
rect 299954 159180 299964 159236
rect 300020 159180 549612 159236
rect 549668 159180 549678 159236
rect 287634 159068 287644 159124
rect 287700 159068 540876 159124
rect 540932 159068 540942 159124
rect 289650 158956 289660 159012
rect 289716 158956 544348 159012
rect 544404 158956 544414 159012
rect 288306 158844 288316 158900
rect 288372 158844 548268 158900
rect 548324 158844 548334 158900
rect 300402 158732 300412 158788
rect 300468 158732 561372 158788
rect 561428 158732 561438 158788
rect 338482 158620 338492 158676
rect 338548 158620 357868 158676
rect 357924 158620 357934 158676
rect 324342 157836 324380 157892
rect 324436 157836 324446 157892
rect 330614 157836 330652 157892
rect 330708 157836 330718 157892
rect 332182 157836 332220 157892
rect 332276 157836 332286 157892
rect 335346 157836 335356 157892
rect 335412 157836 346108 157892
rect 346164 157836 346174 157892
rect 357858 157836 357868 157892
rect 357924 157836 560140 157892
rect 560196 157836 560206 157892
rect 317314 157724 317324 157780
rect 317380 157724 327516 157780
rect 327572 157724 327582 157780
rect 341618 157724 341628 157780
rect 341684 157724 354508 157780
rect 354564 157724 561148 157780
rect 561204 157724 561214 157780
rect 310258 157612 310268 157668
rect 310324 157612 319676 157668
rect 319732 157612 319742 157668
rect 321234 157612 321244 157668
rect 321300 157612 346444 157668
rect 346500 157612 346510 157668
rect 352482 157612 352492 157668
rect 352548 157612 560252 157668
rect 560308 157612 560318 157668
rect 269864 157500 273868 157556
rect 273924 157500 273934 157556
rect 317090 157500 317100 157556
rect 317156 157500 325948 157556
rect 326004 157500 326014 157556
rect 336914 157500 336924 157556
rect 336980 157500 347788 157556
rect 347844 157500 559916 157556
rect 559972 157500 559982 157556
rect 346098 157388 346108 157444
rect 346164 157388 346780 157444
rect 346836 157388 559804 157444
rect 559860 157388 559870 157444
rect 333778 157276 333788 157332
rect 333844 157276 351484 157332
rect 351540 157276 564732 157332
rect 564788 157276 564798 157332
rect 350690 157164 350700 157220
rect 350756 157164 559692 157220
rect 559748 157164 559758 157220
rect 346210 157052 346220 157108
rect 346276 157052 560028 157108
rect 560084 157052 560094 157108
rect 318098 156940 318108 156996
rect 318164 156940 351148 156996
rect 351204 156940 351214 156996
rect 322802 156828 322812 156884
rect 322868 156828 352828 156884
rect 352884 156828 352894 156884
rect 420914 156380 420924 156436
rect 420980 156380 422492 156436
rect 422548 156380 422558 156436
rect 421698 156268 421708 156324
rect 421764 156268 422604 156324
rect 422660 156268 473004 156324
rect 473060 156268 473070 156324
rect 304994 156156 305004 156212
rect 305060 156156 526764 156212
rect 526820 156156 526830 156212
rect 308690 156044 308700 156100
rect 308756 156044 530796 156100
rect 530852 156044 530862 156100
rect 280242 155932 280252 155988
rect 280308 155932 503916 155988
rect 503972 155932 503982 155988
rect 303986 155820 303996 155876
rect 304052 155820 528108 155876
rect 528164 155820 528174 155876
rect 301634 155708 301644 155764
rect 301700 155708 529452 155764
rect 529508 155708 529518 155764
rect 294802 155596 294812 155652
rect 294868 155596 544236 155652
rect 544292 155596 544302 155652
rect 282930 155484 282940 155540
rect 282996 155484 537516 155540
rect 537572 155484 537582 155540
rect 297042 155372 297052 155428
rect 297108 155372 564620 155428
rect 564676 155372 564686 155428
rect 420802 154924 420812 154980
rect 420868 154924 422716 154980
rect 422772 154924 422782 154980
rect 269864 154588 270956 154644
rect 271012 154588 271022 154644
rect 273410 154476 273420 154532
rect 273476 154476 273868 154532
rect 275426 154476 275436 154532
rect 275492 154476 356188 154532
rect 356244 154476 357196 154532
rect 357252 154476 357262 154532
rect 472994 154476 473004 154532
rect 473060 154476 559468 154532
rect 559524 154476 559534 154532
rect 273812 154420 273868 154476
rect 273812 154364 274652 154420
rect 274708 154364 356972 154420
rect 357028 154364 361228 154420
rect 474338 154364 474348 154420
rect 474404 154364 558908 154420
rect 558964 154364 558974 154420
rect 273186 154252 273196 154308
rect 273252 154252 273980 154308
rect 274036 154252 275436 154308
rect 275492 154252 275502 154308
rect 345202 153804 345212 153860
rect 345268 153804 357756 153860
rect 357812 153804 357822 153860
rect 361172 153748 361228 154364
rect 490578 154252 490588 154308
rect 490644 154252 491820 154308
rect 491876 154252 491886 154308
rect 544338 154252 544348 154308
rect 544404 154252 550956 154308
rect 551012 154252 551022 154308
rect 422482 154140 422492 154196
rect 422548 154140 466284 154196
rect 466340 154140 466350 154196
rect 546578 154140 546588 154196
rect 546644 154140 552300 154196
rect 552356 154140 552366 154196
rect 422706 154028 422716 154084
rect 422772 154028 467852 154084
rect 467908 154028 467918 154084
rect 488898 154028 488908 154084
rect 488964 154028 490476 154084
rect 490532 154028 490542 154084
rect 540866 154028 540876 154084
rect 540932 154028 546924 154084
rect 546980 154028 546990 154084
rect 422930 153916 422940 153972
rect 422996 153916 468972 153972
rect 469028 153916 469038 153972
rect 503906 153916 503916 153972
rect 503972 153916 532140 153972
rect 532196 153916 532206 153972
rect 423154 153804 423164 153860
rect 423220 153804 469532 153860
rect 469588 153804 469598 153860
rect 471650 153804 471660 153860
rect 471716 153804 559580 153860
rect 559636 153804 559646 153860
rect 361172 153692 505260 153748
rect 505316 153692 505326 153748
rect 524178 153692 524188 153748
rect 524244 153692 545580 153748
rect 545636 153692 545646 153748
rect 272486 153580 272524 153636
rect 272580 153580 273756 153636
rect 273812 153580 273822 153636
rect 502292 153580 509292 153636
rect 509348 153580 509358 153636
rect 502292 153524 502348 153580
rect 350578 153468 350588 153524
rect 350644 153468 502348 153524
rect 356178 153356 356188 153412
rect 356244 153356 357644 153412
rect 357700 153356 506604 153412
rect 506660 153356 506670 153412
rect 506818 153356 506828 153412
rect 506884 153356 542892 153412
rect 542948 153356 542958 153412
rect 423266 153244 423276 153300
rect 423332 153244 471660 153300
rect 471716 153244 471726 153300
rect 493126 153244 493164 153300
rect 493220 153244 493230 153300
rect 503906 153244 503916 153300
rect 503972 153244 525420 153300
rect 525476 153244 525486 153300
rect 505586 153132 505596 153188
rect 505652 153132 534828 153188
rect 534884 153132 534894 153188
rect 350466 153020 350476 153076
rect 350532 153020 507948 153076
rect 508004 153020 508014 153076
rect 508162 153020 508172 153076
rect 508228 153020 540204 153076
rect 540260 153020 540270 153076
rect 502534 152908 502572 152964
rect 502628 152908 502638 152964
rect 503094 152908 503132 152964
rect 503188 152908 503198 152964
rect 532578 152908 532588 152964
rect 532644 152908 541548 152964
rect 541604 152908 541614 152964
rect 281586 152796 281596 152852
rect 281652 152796 505596 152852
rect 505652 152796 505662 152852
rect 353938 152684 353948 152740
rect 354004 152684 563612 152740
rect 563668 152684 563678 152740
rect 348562 152572 348572 152628
rect 348628 152572 563724 152628
rect 563780 152572 563790 152628
rect 595560 152516 597000 152712
rect 304882 152460 304892 152516
rect 304948 152488 597000 152516
rect 304948 152460 595672 152488
rect 293234 152348 293244 152404
rect 293300 152348 533484 152404
rect 533540 152348 533550 152404
rect 271506 152236 271516 152292
rect 271572 152236 514668 152292
rect 514724 152236 514734 152292
rect 283602 152124 283612 152180
rect 283668 152124 538860 152180
rect 538916 152124 538926 152180
rect 294354 152012 294364 152068
rect 294420 152012 561596 152068
rect 561652 152012 561662 152068
rect 357074 151900 357084 151956
rect 357140 151900 421708 151956
rect 421764 151900 423276 151956
rect 423332 151900 423342 151956
rect 345314 151788 345324 151844
rect 345380 151788 356188 151844
rect 356244 151788 356254 151844
rect 269864 151676 278908 151732
rect 278964 151676 278974 151732
rect 459442 151228 459452 151284
rect 459508 151228 475692 151284
rect 475748 151228 475758 151284
rect 352902 151116 352940 151172
rect 352996 151116 353006 151172
rect 284946 151004 284956 151060
rect 285012 151004 532588 151060
rect 532644 151004 532654 151060
rect 276882 150892 276892 150948
rect 276948 150892 503916 150948
rect 503972 150892 503982 150948
rect 284274 150780 284284 150836
rect 284340 150780 508172 150836
rect 508228 150780 508238 150836
rect 290994 150668 291004 150724
rect 291060 150668 552636 150724
rect 552692 150668 552702 150724
rect 349234 150556 349244 150612
rect 349300 150556 563164 150612
rect 563220 150556 563230 150612
rect 348674 150444 348684 150500
rect 348740 150444 563500 150500
rect 563556 150444 563566 150500
rect 291666 150332 291676 150388
rect 291732 150332 561484 150388
rect 561540 150332 561550 150388
rect 506790 150220 506828 150276
rect 506884 150220 506894 150276
rect -960 149716 480 149912
rect 463362 149772 463372 149828
rect 463428 149772 481068 149828
rect 481124 149772 481134 149828
rect -960 149688 32732 149716
rect 392 149660 32732 149688
rect 32788 149660 32798 149716
rect 482066 149660 482076 149716
rect 482132 149660 562828 149716
rect 562884 149660 562894 149716
rect 303538 149548 303548 149604
rect 303604 149548 536172 149604
rect 536228 149548 536238 149604
rect 295698 149436 295708 149492
rect 295764 149436 561260 149492
rect 561316 149436 561326 149492
rect 478772 149324 502348 149380
rect 478772 149268 478828 149324
rect 502292 149268 502348 149324
rect 296370 149212 296380 149268
rect 296436 149212 478828 149268
rect 501218 149212 501228 149268
rect 501284 149212 501294 149268
rect 502292 149212 559468 149268
rect 559524 149212 559534 149268
rect 285618 149100 285628 149156
rect 285684 149100 501004 149156
rect 501060 149100 501070 149156
rect 501228 149044 501284 149212
rect 501442 149100 501452 149156
rect 501508 149100 506828 149156
rect 506884 149100 506894 149156
rect 462018 148988 462028 149044
rect 462084 148988 501284 149044
rect 349346 148876 349356 148932
rect 349412 148876 562940 148932
rect 562996 148876 563006 148932
rect 269864 148764 275772 148820
rect 275828 148764 275838 148820
rect 348786 148764 348796 148820
rect 348852 148764 563052 148820
rect 563108 148764 563118 148820
rect 299058 148652 299068 148708
rect 299124 148652 559580 148708
rect 559636 148652 559646 148708
rect 457986 148540 457996 148596
rect 458052 148540 460068 148596
rect 460012 147896 460068 148540
rect 341842 146972 341852 147028
rect 341908 146972 357644 147028
rect 357700 146972 357710 147028
rect 269836 145348 269892 145880
rect 273298 145404 273308 145460
rect 273364 145404 307356 145460
rect 307412 145404 307422 145460
rect 269836 145292 272300 145348
rect 272356 145292 350700 145348
rect 350756 145292 350766 145348
rect 358978 145068 358988 145124
rect 359044 145068 459396 145124
rect 459340 145012 460040 145068
rect 273522 143724 273532 143780
rect 273588 143724 350252 143780
rect 350308 143724 350318 143780
rect 269266 143612 269276 143668
rect 269332 143612 417116 143668
rect 417172 143612 417182 143668
rect 269864 142940 272412 142996
rect 272468 142940 273532 142996
rect 273588 142940 273598 142996
rect 559944 142940 561260 142996
rect 561316 142940 561326 142996
rect 354274 142156 354284 142212
rect 354340 142156 459396 142212
rect 459340 142100 460040 142156
rect 559682 142044 559692 142100
rect 559748 142044 559758 142100
rect 274642 141932 274652 141988
rect 274708 141932 356972 141988
rect 357028 141932 357038 141988
rect 559692 141400 559748 142044
rect 559916 140588 560028 140644
rect 560084 140588 560094 140644
rect 269378 140028 269388 140084
rect 269444 140028 345324 140084
rect 345380 140028 345390 140084
rect 559916 139832 559972 140588
rect 595560 139300 597000 139496
rect 356066 139244 356076 139300
rect 356132 139244 459396 139300
rect 575362 139244 575372 139300
rect 575428 139272 597000 139300
rect 575428 139244 595672 139272
rect 459340 139188 460040 139244
rect 276546 138572 276556 138628
rect 276612 138572 357084 138628
rect 357140 138572 357150 138628
rect 559944 138236 561148 138292
rect 561204 138236 561214 138292
rect 269864 137116 273420 137172
rect 273476 137116 273486 137172
rect 559944 136668 560252 136724
rect 560308 136668 560318 136724
rect 354162 136332 354172 136388
rect 354228 136332 459396 136388
rect 459340 136276 460040 136332
rect 392 135800 4620 135828
rect -960 135772 4620 135800
rect 4676 135772 4686 135828
rect -960 135576 480 135772
rect 559944 135100 560140 135156
rect 560196 135100 560206 135156
rect 559906 134316 559916 134372
rect 559972 134316 559982 134372
rect 269864 134204 273196 134260
rect 273252 134204 273262 134260
rect 307010 133868 307020 133924
rect 307076 133868 405020 133924
rect 405076 133868 405086 133924
rect 303090 133756 303100 133812
rect 303156 133756 407036 133812
rect 407092 133756 407102 133812
rect 303650 133644 303660 133700
rect 303716 133644 409052 133700
rect 409108 133644 409118 133700
rect 303874 133532 303884 133588
rect 303940 133532 411068 133588
rect 411124 133532 411134 133588
rect 559916 133560 559972 134316
rect 352146 133420 352156 133476
rect 352212 133420 459396 133476
rect 459340 133364 460040 133420
rect 559794 132524 559804 132580
rect 559860 132524 559870 132580
rect 278226 131964 278236 132020
rect 278292 131964 357308 132020
rect 357364 131964 357374 132020
rect 559804 131992 559860 132524
rect 355730 131852 355740 131908
rect 355796 131852 457660 131908
rect 457716 131852 457726 131908
rect 269864 131292 272524 131348
rect 272580 131292 272590 131348
rect 457650 130508 457660 130564
rect 457716 130508 459396 130564
rect 459340 130452 460040 130508
rect 303426 130396 303436 130452
rect 303492 130396 378812 130452
rect 378868 130396 378878 130452
rect 559944 130396 564732 130452
rect 564788 130396 564798 130452
rect 307122 130284 307132 130340
rect 307188 130284 400988 130340
rect 401044 130284 401054 130340
rect 306786 130172 306796 130228
rect 306852 130172 403004 130228
rect 403060 130172 403070 130228
rect 559944 128828 566188 128884
rect 566244 128828 566254 128884
rect 348450 128492 348460 128548
rect 348516 128492 458108 128548
rect 458164 128492 458174 128548
rect 269864 128380 273308 128436
rect 273364 128380 273374 128436
rect 356738 127596 356748 127652
rect 356804 127596 459396 127652
rect 459340 127540 460040 127596
rect 303202 127372 303212 127428
rect 303268 127372 376796 127428
rect 376852 127372 376862 127428
rect 307234 127260 307244 127316
rect 307300 127260 392924 127316
rect 392980 127260 392990 127316
rect 559944 127260 561372 127316
rect 561428 127260 561438 127316
rect 306898 127148 306908 127204
rect 306964 127148 396956 127204
rect 397012 127148 397022 127204
rect 306674 127036 306684 127092
rect 306740 127036 398972 127092
rect 399028 127036 399038 127092
rect 358866 126924 358876 126980
rect 358932 126924 458220 126980
rect 458276 126924 458286 126980
rect 273746 126812 273756 126868
rect 273812 126812 345212 126868
rect 345268 126812 345278 126868
rect 350578 126812 350588 126868
rect 350644 126812 457996 126868
rect 458052 126812 458062 126868
rect 595560 126056 597000 126280
rect 559944 125692 561260 125748
rect 561316 125692 561326 125748
rect 269864 125468 273756 125524
rect 273812 125468 273822 125524
rect 352594 124684 352604 124740
rect 352660 124684 459396 124740
rect 459340 124628 460040 124684
rect 559570 124348 559580 124404
rect 559636 124348 559646 124404
rect 301522 124236 301532 124292
rect 301588 124236 362684 124292
rect 362740 124236 362750 124292
rect 306562 124124 306572 124180
rect 306628 124124 370748 124180
rect 370804 124124 370814 124180
rect 559580 124152 559636 124348
rect 303314 124012 303324 124068
rect 303380 124012 368732 124068
rect 368788 124012 368798 124068
rect 298162 123900 298172 123956
rect 298228 123900 364700 123956
rect 364756 123900 364766 123956
rect 310034 123788 310044 123844
rect 310100 123788 382844 123844
rect 382900 123788 382910 123844
rect 296482 123676 296492 123732
rect 296548 123676 374780 123732
rect 374836 123676 374846 123732
rect 293122 123564 293132 123620
rect 293188 123564 372764 123620
rect 372820 123564 372830 123620
rect 299842 123452 299852 123508
rect 299908 123452 380828 123508
rect 380884 123452 380894 123508
rect 308242 123340 308252 123396
rect 308308 123340 366716 123396
rect 366772 123340 366782 123396
rect 384822 122668 384860 122724
rect 384916 122668 384926 122724
rect 386838 122668 386876 122724
rect 386932 122668 386942 122724
rect 388854 122668 388892 122724
rect 388948 122668 388958 122724
rect 390870 122668 390908 122724
rect 390964 122668 390974 122724
rect 394902 122668 394940 122724
rect 394996 122668 395006 122724
rect 411618 122668 411628 122724
rect 411684 122668 413084 122724
rect 413140 122668 413150 122724
rect 414950 122668 414988 122724
rect 415044 122668 415054 122724
rect 269864 122556 341852 122612
rect 341908 122556 341918 122612
rect 559944 122556 564508 122612
rect 564564 122556 564574 122612
rect 355954 122108 355964 122164
rect 356020 122108 457996 122164
rect 458052 122108 458062 122164
rect 353826 121996 353836 122052
rect 353892 121996 458220 122052
rect 458276 121996 458286 122052
rect 346882 121884 346892 121940
rect 346948 121884 457660 121940
rect 457716 121884 457726 121940
rect 349122 121772 349132 121828
rect 349188 121772 459396 121828
rect 459340 121716 460040 121772
rect 392 121688 4172 121716
rect -960 121660 4172 121688
rect 4228 121660 4238 121716
rect -960 121464 480 121660
rect 559944 120988 566188 121044
rect 566244 120988 566254 121044
rect 359314 120428 359324 120484
rect 359380 120428 421708 120484
rect 421764 120428 421774 120484
rect 353938 120316 353948 120372
rect 354004 120316 457884 120372
rect 457940 120316 457950 120372
rect 352594 120204 352604 120260
rect 352660 120204 458108 120260
rect 458164 120204 458174 120260
rect 352034 120092 352044 120148
rect 352100 120092 458332 120148
rect 458388 120092 458398 120148
rect 269864 119644 310156 119700
rect 310212 119644 310222 119700
rect 559944 119420 564620 119476
rect 564676 119420 564686 119476
rect 350242 119308 350252 119364
rect 350308 119308 421932 119364
rect 421988 119308 421998 119364
rect 457650 118860 457660 118916
rect 457716 118860 459396 118916
rect 459340 118804 460040 118860
rect 359986 118748 359996 118804
rect 360052 118748 421820 118804
rect 421876 118748 421886 118804
rect 362002 118636 362012 118692
rect 362068 118636 458556 118692
rect 458612 118636 458622 118692
rect 361778 118524 361788 118580
rect 361844 118524 457660 118580
rect 457716 118524 457726 118580
rect 355506 118412 355516 118468
rect 355572 118412 457548 118468
rect 457604 118412 457614 118468
rect 559458 118412 559468 118468
rect 559524 118412 559534 118468
rect 559468 117880 559524 118412
rect 458518 117516 458556 117572
rect 458612 117516 458622 117572
rect 360434 117068 360444 117124
rect 360500 117068 458332 117124
rect 458388 117068 458398 117124
rect 359538 116956 359548 117012
rect 359604 116956 457772 117012
rect 457828 116956 457838 117012
rect 457650 116844 457660 116900
rect 457716 116844 458444 116900
rect 458500 116844 458510 116900
rect 269864 116732 309932 116788
rect 309988 116732 309998 116788
rect 559944 116284 564732 116340
rect 564788 116284 564798 116340
rect 419944 116060 421708 116116
rect 421764 116060 425852 116116
rect 425908 116060 425918 116116
rect 459340 115892 460040 115948
rect 457650 115836 457660 115892
rect 457716 115836 459396 115892
rect 559944 114716 561596 114772
rect 561652 114716 561662 114772
rect 269864 113820 312060 113876
rect 312116 113820 312126 113876
rect 559944 113148 564620 113204
rect 564676 113148 564686 113204
rect 458098 113036 458108 113092
rect 458164 113036 459396 113092
rect 590594 113036 590604 113092
rect 590660 113064 595672 113092
rect 590660 113036 597000 113064
rect 459340 112980 460040 113036
rect 595560 112840 597000 113036
rect 559944 111580 560364 111636
rect 560420 111580 560430 111636
rect 269864 110908 273308 110964
rect 273364 110908 273374 110964
rect 458210 110124 458220 110180
rect 458276 110124 459396 110180
rect 459340 110068 460040 110124
rect 559944 110012 564508 110068
rect 564564 110012 564574 110068
rect 419944 109116 421820 109172
rect 421876 109116 424172 109172
rect 424228 109116 424238 109172
rect 559944 108444 561484 108500
rect 561540 108444 561550 108500
rect 356962 108220 356972 108276
rect 357028 108220 357532 108276
rect 357588 108220 360136 108276
rect 269864 107996 311948 108052
rect 312004 107996 312014 108052
rect -960 107380 480 107576
rect -960 107352 29372 107380
rect 392 107324 29372 107352
rect 29428 107324 29438 107380
rect 457986 107212 457996 107268
rect 458052 107212 459396 107268
rect 459340 107156 460040 107212
rect 559944 106876 563164 106932
rect 563220 106876 563230 106932
rect 559944 105308 561148 105364
rect 561204 105308 561214 105364
rect 269864 105084 311052 105140
rect 311108 105084 311118 105140
rect 458546 104300 458556 104356
rect 458612 104300 459396 104356
rect 459340 104244 460040 104300
rect 559944 103740 563388 103796
rect 563444 103740 563454 103796
rect 419916 102396 421932 102452
rect 421988 102396 459452 102452
rect 459508 102396 459518 102452
rect 269864 102172 273084 102228
rect 273140 102172 273150 102228
rect 419916 102200 419972 102396
rect 559944 102172 563276 102228
rect 563332 102172 563342 102228
rect 273298 101612 273308 101668
rect 273364 101612 350252 101668
rect 350308 101612 350318 101668
rect 457874 101388 457884 101444
rect 457940 101388 459396 101444
rect 459340 101332 460040 101388
rect 559944 100604 563052 100660
rect 563108 100604 563118 100660
rect 585442 99820 585452 99876
rect 585508 99848 595672 99876
rect 585508 99820 597000 99848
rect 595560 99624 597000 99820
rect 269864 99260 272972 99316
rect 273028 99260 273038 99316
rect 559944 99036 563724 99092
rect 563780 99036 563790 99092
rect 458546 98476 458556 98532
rect 458612 98476 459396 98532
rect 459340 98420 460040 98476
rect 559944 97468 562940 97524
rect 562996 97468 563006 97524
rect 269864 96348 311164 96404
rect 311220 96348 311230 96404
rect 559906 95900 559916 95956
rect 559972 95900 559982 95956
rect 457650 95564 457660 95620
rect 457716 95564 459396 95620
rect 459340 95508 460040 95564
rect 419944 95228 420140 95284
rect 420196 95228 421820 95284
rect 421876 95228 421886 95284
rect 559944 94332 563612 94388
rect 563668 94332 563678 94388
rect 392 93464 4396 93492
rect -960 93436 4396 93464
rect 4452 93436 4462 93492
rect 269864 93436 356972 93492
rect 357028 93436 357038 93492
rect -960 93240 480 93436
rect 559944 92764 562828 92820
rect 562884 92764 562894 92820
rect 457762 92652 457772 92708
rect 457828 92652 459396 92708
rect 459340 92596 460040 92652
rect 559944 91196 563500 91252
rect 563556 91196 563566 91252
rect 269864 90524 279692 90580
rect 279748 90524 279758 90580
rect 458434 89740 458444 89796
rect 458500 89740 459396 89796
rect 459340 89684 460040 89740
rect 559794 89628 559804 89684
rect 559860 89628 559870 89684
rect 419944 88284 420140 88340
rect 420196 88284 422604 88340
rect 422660 88284 422670 88340
rect 559944 88060 563164 88116
rect 563220 88060 563230 88116
rect 269864 87612 315196 87668
rect 315252 87612 315262 87668
rect 458322 86828 458332 86884
rect 458388 86828 459396 86884
rect 459340 86772 460040 86828
rect 559944 86492 563052 86548
rect 563108 86492 563118 86548
rect 595560 86408 597000 86632
rect 350242 84924 350252 84980
rect 350308 84924 360136 84980
rect 559794 84924 559804 84980
rect 559860 84924 559870 84980
rect 269864 84700 330092 84756
rect 330148 84700 330158 84756
rect 457874 83916 457884 83972
rect 457940 83916 459396 83972
rect 459340 83860 460040 83916
rect 559944 83356 562828 83412
rect 562884 83356 562894 83412
rect 269864 81788 274652 81844
rect 274708 81788 274718 81844
rect 559944 81788 563500 81844
rect 563556 81788 563566 81844
rect 419944 81340 421708 81396
rect 421764 81340 421774 81396
rect 457762 81004 457772 81060
rect 457828 81004 459396 81060
rect 459340 80948 460040 81004
rect 559944 80220 562940 80276
rect 562996 80220 563006 80276
rect -960 79156 480 79352
rect -960 79128 14252 79156
rect 392 79100 14252 79128
rect 14308 79100 14318 79156
rect 269864 78876 278236 78932
rect 278292 78876 278302 78932
rect 559570 78652 559580 78708
rect 559636 78652 559646 78708
rect 458210 78092 458220 78148
rect 458276 78092 459396 78148
rect 459340 78036 460040 78092
rect 559682 77084 559692 77140
rect 559748 77084 559758 77140
rect 269864 75964 276556 76020
rect 276612 75964 276622 76020
rect 559458 75516 559468 75572
rect 559524 75516 559534 75572
rect 458098 75180 458108 75236
rect 458164 75180 459396 75236
rect 459340 75124 460040 75180
rect 419944 74396 420252 74452
rect 420308 74396 423164 74452
rect 423220 74396 423230 74452
rect 559944 73948 562940 74004
rect 562996 73948 563006 74004
rect 590482 73388 590492 73444
rect 590548 73416 595672 73444
rect 590548 73388 597000 73416
rect 595560 73192 597000 73388
rect 269864 73052 273308 73108
rect 273364 73052 273374 73108
rect 559944 72380 563388 72436
rect 563444 72380 563454 72436
rect 459340 72212 460040 72268
rect 457986 72156 457996 72212
rect 458052 72156 459396 72212
rect 559944 70812 562828 70868
rect 562884 70812 562894 70868
rect 269864 70140 273084 70196
rect 273140 70140 273150 70196
rect 459340 69300 460040 69356
rect 457762 69244 457772 69300
rect 457828 69244 459396 69300
rect 559944 69244 563724 69300
rect 563780 69244 563790 69300
rect 421810 68796 421820 68852
rect 421876 68796 422940 68852
rect 422996 68796 423006 68852
rect 559944 67676 563164 67732
rect 563220 67676 563230 67732
rect 419944 67452 421820 67508
rect 421876 67452 421886 67508
rect 269864 67228 272972 67284
rect 273028 67228 273038 67284
rect 459340 66388 460040 66444
rect 424162 66332 424172 66388
rect 424228 66332 457660 66388
rect 457716 66332 457726 66388
rect 457874 66332 457884 66388
rect 457940 66332 459396 66388
rect 559944 66108 563052 66164
rect 563108 66108 563118 66164
rect -960 65044 480 65240
rect -960 65016 20972 65044
rect 392 64988 20972 65016
rect 21028 64988 21038 65044
rect 559944 64540 563164 64596
rect 563220 64540 563230 64596
rect 269864 64316 276556 64372
rect 276612 64316 276622 64372
rect 459340 63476 460040 63532
rect 457986 63420 457996 63476
rect 458052 63420 459396 63476
rect 559944 62972 563276 63028
rect 563332 62972 563342 63028
rect 357746 61628 357756 61684
rect 357812 61628 360136 61684
rect 269864 61404 273196 61460
rect 273252 61404 273262 61460
rect 559944 61404 563612 61460
rect 563668 61404 563678 61460
rect 425842 60620 425852 60676
rect 425908 60620 459396 60676
rect 459340 60564 460040 60620
rect 419944 60508 421932 60564
rect 421988 60508 422716 60564
rect 422772 60508 422782 60564
rect 595560 60004 597000 60200
rect 573682 59948 573692 60004
rect 573748 59976 597000 60004
rect 573748 59948 595672 59976
rect 559944 59836 562940 59892
rect 562996 59836 563006 59892
rect 269864 58492 275436 58548
rect 275492 58492 275502 58548
rect 559944 58268 562828 58324
rect 562884 58268 562894 58324
rect 457650 57708 457660 57764
rect 457716 57708 459396 57764
rect 459340 57652 460040 57708
rect 559468 56084 559524 56728
rect 559458 56028 559468 56084
rect 559524 56028 559534 56084
rect 269864 55580 288988 55636
rect 289044 55580 289054 55636
rect 459340 54740 460040 54796
rect 457650 54684 457660 54740
rect 457716 54684 459396 54740
rect 419384 53592 422492 53620
rect 419356 53564 422492 53592
rect 422548 53564 422558 53620
rect 419356 53060 419412 53564
rect 419234 53004 419244 53060
rect 419300 53004 419412 53060
rect 355394 52892 355404 52948
rect 355460 52892 457996 52948
rect 458052 52892 458062 52948
rect 273074 52780 273084 52836
rect 273140 52780 420028 52836
rect 420084 52780 420094 52836
rect 269864 52668 275548 52724
rect 275604 52668 275614 52724
rect 358642 52668 358652 52724
rect 358708 52668 457772 52724
rect 457828 52668 457838 52724
rect 289762 51996 289772 52052
rect 289828 51996 457660 52052
rect 457716 51996 457726 52052
rect 356178 51884 356188 51940
rect 356244 51884 357756 51940
rect 357812 51884 459396 51940
rect 459340 51828 460040 51884
rect 353826 51436 353836 51492
rect 353892 51436 457884 51492
rect 457940 51436 457950 51492
rect 392 51128 4284 51156
rect -960 51100 4284 51128
rect 4340 51100 4350 51156
rect -960 50904 480 51100
rect 275538 50652 275548 50708
rect 275604 50652 419244 50708
rect 419300 50652 419310 50708
rect 272962 50540 272972 50596
rect 273028 50540 420140 50596
rect 420196 50540 420206 50596
rect 288978 50428 288988 50484
rect 289044 50428 421932 50484
rect 421988 50428 421998 50484
rect 14242 50316 14252 50372
rect 14308 50316 272412 50372
rect 272468 50316 272478 50372
rect 307430 50316 307468 50372
rect 307524 50316 307534 50372
rect 315270 50316 315308 50372
rect 315364 50316 315374 50372
rect 347666 50316 347676 50372
rect 347732 50316 563276 50372
rect 563332 50316 563342 50372
rect 351026 50204 351036 50260
rect 351092 50204 559468 50260
rect 559524 50204 559534 50260
rect 351922 50092 351932 50148
rect 351988 50092 563052 50148
rect 563108 50092 563118 50148
rect 353714 49980 353724 50036
rect 353780 49980 562940 50036
rect 562996 49980 563006 50036
rect 356066 49868 356076 49924
rect 356132 49868 562828 49924
rect 562884 49868 562894 49924
rect 197922 49756 197932 49812
rect 197988 49756 273980 49812
rect 274036 49756 274046 49812
rect 275426 49756 275436 49812
rect 275492 49756 421820 49812
rect 421876 49756 421886 49812
rect 123666 49644 123676 49700
rect 123732 49644 269500 49700
rect 269556 49644 269566 49700
rect 273186 49644 273196 49700
rect 273252 49644 420252 49700
rect 420308 49644 420318 49700
rect 46946 49532 46956 49588
rect 47012 49532 53228 49588
rect 53284 49532 53294 49588
rect 95106 49532 95116 49588
rect 95172 49532 269836 49588
rect 269892 49532 269902 49588
rect 276546 49532 276556 49588
rect 276612 49532 422044 49588
rect 422100 49532 422110 49588
rect 184772 48748 267148 48804
rect 267204 48748 267214 48804
rect 184772 48692 184828 48748
rect 97346 48636 97356 48692
rect 97412 48636 184828 48692
rect 267092 48692 267148 48748
rect 267092 48636 293580 48692
rect 293636 48636 356188 48692
rect 356244 48636 356254 48692
rect 201730 48524 201740 48580
rect 201796 48524 269388 48580
rect 269444 48524 269454 48580
rect 290210 48524 290220 48580
rect 290276 48524 300748 48580
rect 300804 48524 300814 48580
rect 315074 48524 315084 48580
rect 315140 48524 322252 48580
rect 322308 48524 322318 48580
rect 347554 48524 347564 48580
rect 347620 48524 563388 48580
rect 563444 48524 563454 48580
rect 190306 48412 190316 48468
rect 190372 48412 267596 48468
rect 267652 48412 267662 48468
rect 350914 48412 350924 48468
rect 350980 48412 563724 48468
rect 563780 48412 563790 48468
rect 186498 48300 186508 48356
rect 186564 48300 270732 48356
rect 270788 48300 270798 48356
rect 352706 48300 352716 48356
rect 352772 48300 562940 48356
rect 562996 48300 563006 48356
rect 48514 48188 48524 48244
rect 48580 48188 87500 48244
rect 87556 48188 87566 48244
rect 138898 48188 138908 48244
rect 138964 48188 274428 48244
rect 274484 48188 274494 48244
rect 354386 48188 354396 48244
rect 354452 48188 563164 48244
rect 563220 48188 563230 48244
rect 51762 48076 51772 48132
rect 51828 48076 93212 48132
rect 93268 48076 93278 48132
rect 116050 48076 116060 48132
rect 116116 48076 270844 48132
rect 270900 48076 270910 48132
rect 355282 48076 355292 48132
rect 355348 48076 563164 48132
rect 563220 48076 563230 48132
rect 50194 47964 50204 48020
rect 50260 47964 98924 48020
rect 98980 47964 98990 48020
rect 110338 47964 110348 48020
rect 110404 47964 269276 48020
rect 269332 47964 269342 48020
rect 349234 47964 349244 48020
rect 349300 47964 563612 48020
rect 563668 47964 563678 48020
rect 11330 47852 11340 47908
rect 11396 47852 97356 47908
rect 97412 47852 97422 47908
rect 104626 47852 104636 47908
rect 104692 47852 271068 47908
rect 271124 47852 271134 47908
rect 207442 47740 207452 47796
rect 207508 47740 271292 47796
rect 271348 47740 271358 47796
rect 212258 47628 212268 47684
rect 212324 47628 269500 47684
rect 269556 47628 269566 47684
rect 595560 46760 597000 46984
rect 184594 45276 184604 45332
rect 184660 45276 267372 45332
rect 267428 45276 267438 45332
rect 349346 45276 349356 45332
rect 349412 45276 563500 45332
rect 563556 45276 563566 45332
rect 178882 45164 178892 45220
rect 178948 45164 267484 45220
rect 267540 45164 267550 45220
rect 353602 45164 353612 45220
rect 353668 45164 562828 45220
rect 562884 45164 562894 45220
rect 167458 45052 167468 45108
rect 167524 45052 266812 45108
rect 266868 45052 266878 45108
rect 359762 45052 359772 45108
rect 359828 45052 559804 45108
rect 559860 45052 559870 45108
rect 144610 44940 144620 44996
rect 144676 44940 274540 44996
rect 274596 44940 274606 44996
rect 148418 44828 148428 44884
rect 148484 44828 280364 44884
rect 280420 44828 280430 44884
rect 133186 44716 133196 44772
rect 133252 44716 269612 44772
rect 269668 44716 269678 44772
rect 127474 44604 127484 44660
rect 127540 44604 271180 44660
rect 271236 44604 271246 44660
rect 121762 44492 121772 44548
rect 121828 44492 269724 44548
rect 269780 44492 269790 44548
rect 203634 44380 203644 44436
rect 203700 44380 273868 44436
rect 273924 44380 273934 44436
rect 175074 42924 175084 42980
rect 175140 42924 279020 42980
rect 279076 42924 279086 42980
rect 41794 42812 41804 42868
rect 41860 42812 280028 42868
rect 280084 42812 280094 42868
rect 199938 41916 199948 41972
rect 200004 41916 278124 41972
rect 278180 41916 278190 41972
rect 173170 41804 173180 41860
rect 173236 41804 274316 41860
rect 274372 41804 274382 41860
rect 161746 41692 161756 41748
rect 161812 41692 275884 41748
rect 275940 41692 275950 41748
rect 156034 41580 156044 41636
rect 156100 41580 274092 41636
rect 274148 41580 274158 41636
rect 150322 41468 150332 41524
rect 150388 41468 275772 41524
rect 275828 41468 275838 41524
rect 129378 41356 129388 41412
rect 129444 41356 270620 41412
rect 270676 41356 270686 41412
rect 100818 41244 100828 41300
rect 100884 41244 270732 41300
rect 270788 41244 270798 41300
rect 89394 41132 89404 41188
rect 89460 41132 270508 41188
rect 270564 41132 270574 41188
rect 196018 41020 196028 41076
rect 196084 41020 269612 41076
rect 269668 41020 269678 41076
rect 176978 38444 176988 38500
rect 177044 38444 276444 38500
rect 276500 38444 276510 38500
rect 135090 38332 135100 38388
rect 135156 38332 275660 38388
rect 275716 38332 275726 38388
rect 136994 38220 137004 38276
rect 137060 38220 279916 38276
rect 279972 38220 279982 38276
rect 117954 38108 117964 38164
rect 118020 38108 270956 38164
rect 271012 38108 271022 38164
rect 106530 37996 106540 38052
rect 106596 37996 270620 38052
rect 270676 37996 270686 38052
rect 85698 37884 85708 37940
rect 85764 37884 311612 37940
rect 311668 37884 311678 37940
rect 57138 37772 57148 37828
rect 57204 37772 311836 37828
rect 311892 37772 311902 37828
rect -960 36820 480 37016
rect -960 36792 272300 36820
rect 392 36764 272300 36792
rect 272356 36764 272366 36820
rect 125570 34748 125580 34804
rect 125636 34748 283164 34804
rect 283220 34748 283230 34804
rect 108434 34636 108444 34692
rect 108500 34636 286412 34692
rect 286468 34636 286478 34692
rect 102722 34524 102732 34580
rect 102788 34524 286860 34580
rect 286916 34524 286926 34580
rect 97010 34412 97020 34468
rect 97076 34412 286636 34468
rect 286692 34412 286702 34468
rect 595560 33684 597000 33768
rect 279682 33628 279692 33684
rect 279748 33628 597000 33684
rect 595560 33544 597000 33628
rect 188402 31388 188412 31444
rect 188468 31388 278012 31444
rect 278068 31388 278078 31444
rect 159842 31276 159852 31332
rect 159908 31276 279804 31332
rect 279860 31276 279870 31332
rect 131282 31164 131292 31220
rect 131348 31164 283052 31220
rect 283108 31164 283118 31220
rect 119858 31052 119868 31108
rect 119924 31052 289884 31108
rect 289940 31052 289950 31108
rect 169362 29372 169372 29428
rect 169428 29372 278908 29428
rect 278964 29372 278974 29428
rect 62738 27692 62748 27748
rect 62804 27692 309932 27748
rect 309988 27692 309998 27748
rect 140802 26012 140812 26068
rect 140868 26012 275660 26068
rect 275716 26012 275726 26068
rect 192210 24668 192220 24724
rect 192276 24668 269836 24724
rect 269892 24668 269902 24724
rect 79874 24556 79884 24612
rect 79940 24556 274652 24612
rect 274708 24556 274718 24612
rect 68450 24444 68460 24500
rect 68516 24444 276332 24500
rect 276388 24444 276398 24500
rect 74162 24332 74172 24388
rect 74228 24332 289996 24388
rect 290052 24332 290062 24388
rect -960 22708 480 22904
rect -960 22680 27692 22708
rect 392 22652 27692 22680
rect 27748 22652 27758 22708
rect 595560 20356 597000 20552
rect 572002 20300 572012 20356
rect 572068 20328 597000 20356
rect 572068 20300 595672 20328
rect 152226 17612 152236 17668
rect 152292 17612 267260 17668
rect 267316 17612 267326 17668
rect 163650 12572 163660 12628
rect 163716 12572 269724 12628
rect 269780 12572 269790 12628
rect 392 8792 4172 8820
rect -960 8764 4172 8792
rect 4228 8764 4238 8820
rect -960 8568 480 8764
rect 146738 7532 146748 7588
rect 146804 7532 275548 7588
rect 275604 7532 275614 7588
rect 595560 7140 597000 7336
rect 288082 7084 288092 7140
rect 288148 7112 597000 7140
rect 288148 7084 595672 7112
rect 158162 5852 158172 5908
rect 158228 5852 277228 5908
rect 277284 5852 277294 5908
rect 38546 4956 38556 5012
rect 38612 4956 45612 5012
rect 45668 4956 45678 5012
rect 51874 4956 51884 5012
rect 51940 4956 76076 5012
rect 76132 4956 76142 5012
rect 205762 4956 205772 5012
rect 205828 4956 288204 5012
rect 288260 4956 288270 5012
rect 41346 4844 41356 4900
rect 41412 4844 66556 4900
rect 66612 4844 66622 4900
rect 181010 4844 181020 4900
rect 181076 4844 270508 4900
rect 270564 4844 270574 4900
rect 50306 4732 50316 4788
rect 50372 4732 77980 4788
rect 78036 4732 78046 4788
rect 194338 4732 194348 4788
rect 194404 4732 285180 4788
rect 285236 4732 285246 4788
rect 40226 4620 40236 4676
rect 40292 4620 70364 4676
rect 70420 4620 70430 4676
rect 114370 4620 114380 4676
rect 114436 4620 209132 4676
rect 209188 4620 209198 4676
rect 211474 4620 211484 4676
rect 211540 4620 289772 4676
rect 289828 4620 289838 4676
rect 41122 4508 41132 4564
rect 41188 4508 72268 4564
rect 72324 4508 72334 4564
rect 182914 4508 182924 4564
rect 182980 4508 283052 4564
rect 283108 4508 283118 4564
rect 33506 4396 33516 4452
rect 33572 4396 64652 4452
rect 64708 4396 64718 4452
rect 165778 4396 165788 4452
rect 165844 4396 281372 4452
rect 281428 4396 281438 4452
rect 35186 4284 35196 4340
rect 35252 4284 49420 4340
rect 49476 4284 49486 4340
rect 51986 4284 51996 4340
rect 52052 4284 83692 4340
rect 83748 4284 83758 4340
rect 154354 4284 154364 4340
rect 154420 4284 284956 4340
rect 285012 4284 285022 4340
rect 15362 4172 15372 4228
rect 15428 4172 16716 4228
rect 16772 4172 16782 4228
rect 17266 4172 17276 4228
rect 17332 4172 18396 4228
rect 18452 4172 18462 4228
rect 19170 4172 19180 4228
rect 19236 4172 20076 4228
rect 20132 4172 20142 4228
rect 25078 4172 25116 4228
rect 25172 4172 25182 4228
rect 34402 4172 34412 4228
rect 34468 4172 35084 4228
rect 35140 4172 35150 4228
rect 38322 4172 38332 4228
rect 38388 4172 47516 4228
rect 47572 4172 47582 4228
rect 48626 4172 48636 4228
rect 48692 4172 81788 4228
rect 81844 4172 81854 4228
rect 112466 4172 112476 4228
rect 112532 4172 272188 4228
rect 272244 4172 272254 4228
rect 579618 4172 579628 4228
rect 579684 4172 580636 4228
rect 580692 4172 580702 4228
rect 581298 4172 581308 4228
rect 581364 4172 582540 4228
rect 582596 4172 582606 4228
rect 582978 4172 582988 4228
rect 583044 4172 584444 4228
rect 584500 4172 584510 4228
rect 38434 4060 38444 4116
rect 38500 4060 58940 4116
rect 58996 4060 59006 4116
rect 171490 4060 171500 4116
rect 171556 4060 172956 4116
rect 173012 4060 173022 4116
rect 209570 4060 209580 4116
rect 209636 4060 277340 4116
rect 277396 4060 277406 4116
rect 55094 3388 55132 3444
rect 55188 3388 55198 3444
rect 60806 3388 60844 3444
rect 60900 3388 60910 3444
rect 91494 3388 91532 3444
rect 91588 3388 91598 3444
rect 142902 3388 142940 3444
rect 142996 3388 143006 3444
<< via3 >>
rect 560252 591276 560308 591332
rect 193116 591052 193172 591108
rect 193340 590828 193396 590884
rect 194236 590604 194292 590660
rect 511308 590604 511364 590660
rect 514892 590156 514948 590212
rect 584668 590156 584724 590212
rect 590492 588588 590548 588644
rect 183036 575484 183092 575540
rect 590492 575484 590548 575540
rect 184716 567868 184772 567924
rect 590492 567868 590548 567924
rect 511420 566972 511476 567028
rect 556108 565068 556164 565124
rect 585452 562156 585508 562212
rect 4172 558908 4228 558964
rect 552748 555660 552804 555716
rect 556220 550956 556276 551012
rect 590492 549164 590548 549220
rect 556444 536844 556500 536900
rect 565292 535724 565348 535780
rect 186396 529228 186452 529284
rect 556332 527436 556388 527492
rect 549388 522732 549444 522788
rect 568652 522508 568708 522564
rect 184492 522060 184548 522116
rect 4284 516572 4340 516628
rect 590492 509292 590548 509348
rect 183932 500556 183988 500612
rect 551068 494508 551124 494564
rect 549500 489804 549556 489860
rect 187516 486220 187572 486276
rect 566972 482860 567028 482916
rect 187964 479052 188020 479108
rect 4396 474236 4452 474292
rect 590604 469644 590660 469700
rect 4172 469532 4228 469588
rect 177212 469532 177268 469588
rect 4284 467852 4340 467908
rect 180572 467852 180628 467908
rect 4396 466172 4452 466228
rect 175532 466172 175588 466228
rect 187852 457548 187908 457604
rect 570332 456428 570388 456484
rect 187292 436044 187348 436100
rect 177324 431900 177380 431956
rect 590716 430108 590772 430164
rect 185388 428876 185444 428932
rect 190652 421820 190708 421876
rect 551180 414540 551236 414596
rect 359884 410060 359940 410116
rect 193340 409052 193396 409108
rect 339276 408940 339332 408996
rect 359548 408380 359604 408436
rect 243516 407932 243572 407988
rect 357308 407932 357364 407988
rect 193116 407708 193172 407764
rect 533820 407596 533876 407652
rect 539196 407596 539252 407652
rect 248892 407484 248948 407540
rect 356188 407372 356244 407428
rect 362012 407372 362068 407428
rect 557788 407372 557844 407428
rect 357196 407036 357252 407092
rect 357308 406700 357364 406756
rect 227612 406588 227668 406644
rect 266252 406588 266308 406644
rect 270396 406588 270452 406644
rect 276332 406588 276388 406644
rect 281372 406588 281428 406644
rect 286412 406588 286468 406644
rect 323372 406588 323428 406644
rect 335916 406588 335972 406644
rect 357196 406588 357252 406644
rect 194236 405804 194292 405860
rect 359772 404908 359828 404964
rect 357196 404348 357252 404404
rect 511308 404348 511364 404404
rect 359996 403452 360052 403508
rect 186060 402332 186116 402388
rect 590716 402332 590772 402388
rect 348908 401660 348964 401716
rect 184604 401548 184660 401604
rect 590940 401548 590996 401604
rect 361900 399980 361956 400036
rect 360556 399868 360612 399924
rect 471996 398188 472052 398244
rect 519148 398076 519204 398132
rect 375452 397292 375508 397348
rect 511420 397292 511476 397348
rect 526428 396844 526484 396900
rect 532476 396732 532532 396788
rect 359660 396620 359716 396676
rect 556668 396620 556724 396676
rect 550620 396508 550676 396564
rect 227612 395724 227668 395780
rect 362908 395052 362964 395108
rect 538524 394828 538580 394884
rect 405468 394492 405524 394548
rect 441756 394492 441812 394548
rect 438508 394156 438564 394212
rect 438508 393932 438564 393988
rect 362908 392700 362964 392756
rect 360444 392588 360500 392644
rect 361900 392588 361956 392644
rect 405468 392476 405524 392532
rect 361788 392364 361844 392420
rect 471996 392364 472052 392420
rect 362124 392252 362180 392308
rect 216636 391356 216692 391412
rect 215068 390908 215124 390964
rect 358988 390908 359044 390964
rect 590940 390572 590996 390628
rect 359884 389900 359940 389956
rect 4396 389564 4452 389620
rect 359884 389452 359940 389508
rect 359548 389340 359604 389396
rect 359884 388892 359940 388948
rect 329084 388108 329140 388164
rect 342300 385980 342356 386036
rect 338492 385756 338548 385812
rect 110012 385196 110068 385252
rect 186396 383852 186452 383908
rect 343084 383852 343140 383908
rect 197372 383740 197428 383796
rect 199500 383628 199556 383684
rect 99932 383404 99988 383460
rect 340060 383180 340116 383236
rect 349468 383068 349524 383124
rect 231644 382284 231700 382340
rect 198156 382172 198212 382228
rect 199836 382172 199892 382228
rect 201516 382172 201572 382228
rect 208236 382172 208292 382228
rect 209916 382172 209972 382228
rect 230076 382172 230132 382228
rect 231756 382172 231812 382228
rect 277116 382060 277172 382116
rect 305676 382060 305732 382116
rect 307356 382060 307412 382116
rect 319116 382060 319172 382116
rect 320796 382060 320852 382116
rect 324156 382060 324212 382116
rect 329196 382060 329252 382116
rect 330876 382060 330932 382116
rect 334236 382060 334292 382116
rect 196476 381948 196532 382004
rect 198044 381948 198100 382004
rect 199724 381948 199780 382004
rect 201404 381948 201460 382004
rect 204876 381948 204932 382004
rect 206556 381948 206612 382004
rect 206780 381948 206836 382004
rect 199836 381836 199892 381892
rect 199612 381388 199668 381444
rect 206780 381388 206836 381444
rect 336924 380492 336980 380548
rect 346108 380044 346164 380100
rect 347788 379932 347844 379988
rect 210364 379708 210420 379764
rect 236124 379708 236180 379764
rect 196364 379596 196420 379652
rect 202412 379596 202468 379652
rect 342972 379596 343028 379652
rect 253372 379484 253428 379540
rect 336812 379484 336868 379540
rect 196140 379372 196196 379428
rect 196364 379372 196420 379428
rect 221564 379372 221620 379428
rect 221788 379372 221844 379428
rect 222684 379372 222740 379428
rect 235228 379372 235284 379428
rect 237020 379372 237076 379428
rect 238476 379372 238532 379428
rect 250124 379372 250180 379428
rect 249116 379260 249172 379316
rect 264460 379372 264516 379428
rect 192332 379148 192388 379204
rect 202412 379148 202468 379204
rect 221900 379148 221956 379204
rect 249340 379148 249396 379204
rect 250012 379148 250068 379204
rect 264460 379036 264516 379092
rect 222684 378924 222740 378980
rect 253372 378924 253428 378980
rect 197596 378812 197652 378868
rect 210364 378812 210420 378868
rect 221788 378812 221844 378868
rect 182476 377804 182532 377860
rect 590492 377356 590548 377412
rect 4396 377132 4452 377188
rect 182252 377132 182308 377188
rect 187404 376460 187460 376516
rect 354284 376236 354340 376292
rect 357868 376236 357924 376292
rect 4172 375676 4228 375732
rect 184156 375116 184212 375172
rect 180684 373772 180740 373828
rect 344092 373100 344148 373156
rect 184044 372428 184100 372484
rect 344204 372204 344260 372260
rect 185612 371084 185668 371140
rect 339948 367948 340004 368004
rect 357196 367052 357252 367108
rect 185500 364364 185556 364420
rect 345324 363244 345380 363300
rect 182476 363020 182532 363076
rect 345436 360556 345492 360612
rect 187404 359660 187460 359716
rect 340172 359548 340228 359604
rect 178892 358652 178948 358708
rect 185612 358652 185668 358708
rect 184156 356300 184212 356356
rect 356524 354732 356580 354788
rect 345212 353388 345268 353444
rect 180684 352940 180740 352996
rect 341852 350700 341908 350756
rect 184044 350364 184100 350420
rect 357084 348796 357140 348852
rect 357084 347788 357140 347844
rect 357756 347788 357812 347844
rect 4172 347228 4228 347284
rect 345884 347116 345940 347172
rect 342972 344428 343028 344484
rect 344428 343532 344484 343588
rect 348572 343084 348628 343140
rect 357644 343084 357700 343140
rect 344092 341740 344148 341796
rect 344316 339948 344372 340004
rect 178108 339500 178164 339556
rect 339276 337260 339332 337316
rect 339388 336364 339444 336420
rect 354060 335468 354116 335524
rect 344428 334572 344484 334628
rect 355628 333676 355684 333732
rect 350364 332780 350420 332836
rect 352268 331884 352324 331940
rect 348572 330988 348628 331044
rect 359436 330988 359492 331044
rect 346780 330092 346836 330148
rect 346668 329196 346724 329252
rect 353948 328300 354004 328356
rect 350476 327404 350532 327460
rect 348684 326508 348740 326564
rect 178892 326060 178948 326116
rect 352380 325612 352436 325668
rect 356188 325612 356244 325668
rect 357868 325612 357924 325668
rect 181356 325388 181412 325444
rect 347900 324716 347956 324772
rect 348796 323820 348852 323876
rect 190652 323372 190708 323428
rect 350700 322924 350756 322980
rect 175308 322700 175364 322756
rect 187404 322700 187460 322756
rect 353612 322028 353668 322084
rect 175308 321804 175364 321860
rect 174524 321356 174580 321412
rect 348012 321132 348068 321188
rect 348124 320236 348180 320292
rect 178108 320124 178164 320180
rect 174636 320012 174692 320068
rect 360108 319732 360164 319788
rect 344540 319340 344596 319396
rect 174412 318668 174468 318724
rect 339276 318444 339332 318500
rect 359884 317548 359940 317604
rect 177884 317324 177940 317380
rect 353724 316652 353780 316708
rect 179676 315980 179732 316036
rect 346220 315756 346276 315812
rect 342188 314860 342244 314916
rect 184380 314636 184436 314692
rect 349580 313964 349636 314020
rect 177996 313292 178052 313348
rect 339388 313292 339444 313348
rect 358988 313292 359044 313348
rect 352828 313068 352884 313124
rect 351932 312172 351988 312228
rect 174300 311948 174356 312004
rect 355292 311276 355348 311332
rect 590492 311052 590548 311108
rect 185836 310604 185892 310660
rect 346332 310380 346388 310436
rect 339276 309820 339332 309876
rect 339500 309820 339556 309876
rect 190428 309260 190484 309316
rect 351148 308588 351204 308644
rect 357308 308028 357364 308084
rect 185724 307916 185780 307972
rect 357980 307916 358036 307972
rect 354620 307692 354676 307748
rect 349692 306796 349748 306852
rect 4172 306572 4228 306628
rect 168812 306572 168868 306628
rect 181244 306572 181300 306628
rect 352492 305900 352548 305956
rect 184492 305228 184548 305284
rect 339276 305004 339332 305060
rect 167244 304892 167300 304948
rect 354284 304108 354340 304164
rect 63756 303996 63812 304052
rect 78876 303996 78932 304052
rect 93996 303996 94052 304052
rect 187740 303884 187796 303940
rect 339612 303212 339668 303268
rect 186956 302540 187012 302596
rect 354172 302316 354228 302372
rect 350588 302204 350644 302260
rect 350812 302204 350868 302260
rect 352156 301420 352212 301476
rect 186844 301196 186900 301252
rect 355740 300524 355796 300580
rect 182924 299852 182980 299908
rect 356524 299516 356580 299572
rect 345660 298732 345716 298788
rect 187068 298508 187124 298564
rect 342412 297836 342468 297892
rect 187628 297164 187684 297220
rect 346892 296940 346948 296996
rect 4172 296604 4228 296660
rect 172284 296604 172340 296660
rect 187516 296492 187572 296548
rect 346332 296492 346388 296548
rect 165452 296044 165508 296100
rect 359884 296044 359940 296100
rect 187404 295820 187460 295876
rect 340284 295708 340340 295764
rect 187964 295596 188020 295652
rect 351260 295148 351316 295204
rect 187516 294476 187572 294532
rect 354732 293132 354788 293188
rect 342748 292460 342804 292516
rect 121772 291788 121828 291844
rect 343084 290892 343140 290948
rect 352044 290780 352100 290836
rect 342076 290668 342132 290724
rect 138572 290444 138628 290500
rect 165676 290220 165732 290276
rect 187292 289772 187348 289828
rect 342860 289772 342916 289828
rect 355516 289772 355572 289828
rect 167132 289100 167188 289156
rect 339276 288876 339332 288932
rect 342860 288876 342916 288932
rect 190652 288428 190708 288484
rect 342748 287980 342804 288036
rect 120092 287756 120148 287812
rect 341292 287084 341348 287140
rect 188076 286636 188132 286692
rect 113372 286300 113428 286356
rect 190540 285740 190596 285796
rect 354508 285740 354564 285796
rect 182364 285628 182420 285684
rect 183932 285628 183988 285684
rect 187180 285628 187236 285684
rect 118412 285404 118468 285460
rect 355404 284844 355460 284900
rect 339388 284732 339444 284788
rect 342748 284732 342804 284788
rect 346220 284732 346276 284788
rect 346220 284060 346276 284116
rect 358876 284060 358932 284116
rect 342748 283948 342804 284004
rect 355964 283948 356020 284004
rect 348012 283836 348068 283892
rect 172284 283724 172340 283780
rect 348124 283724 348180 283780
rect 182476 283612 182532 283668
rect 348236 283500 348292 283556
rect 167244 282380 167300 282436
rect 186508 282156 186564 282212
rect 352828 282156 352884 282212
rect 182364 281932 182420 281988
rect 175644 281372 175700 281428
rect 339276 281148 339332 281204
rect 168812 281036 168868 281092
rect 187180 280476 187236 280532
rect 186284 280364 186340 280420
rect 187292 280364 187348 280420
rect 190652 280364 190708 280420
rect 353836 280700 353892 280756
rect 358652 280588 358708 280644
rect 354732 280476 354788 280532
rect 354620 280364 354676 280420
rect 339276 280140 339332 280196
rect 182252 279692 182308 279748
rect 339388 279580 339444 279636
rect 165452 279244 165508 279300
rect 168140 279244 168196 279300
rect 186284 279020 186340 279076
rect 342748 279020 342804 279076
rect 168140 278908 168196 278964
rect 355404 278908 355460 278964
rect 342860 278796 342916 278852
rect 177324 278348 177380 278404
rect 341404 278124 341460 278180
rect 168028 278012 168084 278068
rect 185388 278012 185444 278068
rect 165676 277228 165732 277284
rect 168028 277228 168084 277284
rect 185388 277228 185444 277284
rect 187292 277228 187348 277284
rect 341740 277228 341796 277284
rect 175532 277004 175588 277060
rect 341516 276332 341572 276388
rect 190540 275884 190596 275940
rect 180572 275660 180628 275716
rect 342748 275548 342804 275604
rect 344652 275548 344708 275604
rect 339724 275436 339780 275492
rect 339836 274540 339892 274596
rect 177212 274316 177268 274372
rect 356748 273084 356804 273140
rect 357420 273084 357476 273140
rect 356860 272972 356916 273028
rect 182476 272076 182532 272132
rect 344540 272076 344596 272132
rect 590604 271404 590660 271460
rect 342860 270956 342916 271012
rect 339276 270060 339332 270116
rect 170492 269836 170548 269892
rect 342972 269164 343028 269220
rect 175644 268716 175700 268772
rect 357420 268716 357476 268772
rect 339276 267372 339332 267428
rect 357420 267372 357476 267428
rect 186396 265804 186452 265860
rect 359548 264572 359604 264628
rect 168140 263788 168196 263844
rect 4172 262780 4228 262836
rect 168028 261772 168084 261828
rect 357532 261324 357588 261380
rect 183036 260876 183092 260932
rect 339276 260204 339332 260260
rect 339388 259980 339444 260036
rect 184716 259532 184772 259588
rect 339500 258748 339556 258804
rect 186172 258188 186228 258244
rect 339500 257852 339556 257908
rect 356972 256956 357028 257012
rect 357308 256956 357364 257012
rect 185948 256844 186004 256900
rect 351372 256620 351428 256676
rect 341292 255836 341348 255892
rect 359324 255836 359380 255892
rect 341180 255724 341236 255780
rect 357308 255724 357364 255780
rect 186060 255500 186116 255556
rect 339276 254828 339332 254884
rect 184604 254156 184660 254212
rect 342748 253932 342804 253988
rect 187180 252812 187236 252868
rect 339276 252476 339332 252532
rect 344428 252028 344484 252084
rect 187852 251468 187908 251524
rect 340396 251244 340452 251300
rect 339276 250348 339332 250404
rect 190652 249788 190708 249844
rect 356972 249788 357028 249844
rect 357084 249452 357140 249508
rect 190652 248780 190708 248836
rect 343084 248556 343140 248612
rect 347900 248556 347956 248612
rect 4172 248444 4228 248500
rect 342412 248444 342468 248500
rect 349132 248444 349188 248500
rect 342188 247772 342244 247828
rect 190652 247212 190708 247268
rect 339276 247100 339332 247156
rect 339388 246316 339444 246372
rect 341628 245868 341684 245924
rect 190540 244748 190596 244804
rect 190652 242620 190708 242676
rect 349356 241948 349412 242004
rect 338604 241836 338660 241892
rect 339276 241836 339332 241892
rect 335916 241724 335972 241780
rect 198044 241612 198100 241668
rect 335804 241612 335860 241668
rect 337708 241612 337764 241668
rect 322588 241388 322644 241444
rect 345548 241388 345604 241444
rect 187068 241276 187124 241332
rect 273868 241276 273924 241332
rect 318556 241276 318612 241332
rect 187404 241164 187460 241220
rect 278908 241164 278964 241220
rect 288204 241164 288260 241220
rect 317884 241052 317940 241108
rect 359660 241052 359716 241108
rect 334124 240940 334180 240996
rect 304892 240716 304948 240772
rect 334236 240716 334292 240772
rect 317884 240604 317940 240660
rect 318556 240604 318612 240660
rect 322588 240604 322644 240660
rect 323260 240604 323316 240660
rect 350588 240604 350644 240660
rect 197484 240380 197540 240436
rect 336924 240492 336980 240548
rect 338268 240492 338324 240548
rect 197708 240268 197764 240324
rect 337596 240268 337652 240324
rect 344876 240268 344932 240324
rect 358988 240268 359044 240324
rect 48524 240156 48580 240212
rect 197372 240156 197428 240212
rect 320572 240156 320628 240212
rect 359772 240156 359828 240212
rect 314972 240044 315028 240100
rect 319900 240044 319956 240100
rect 337036 239932 337092 239988
rect 338380 239932 338436 239988
rect 182364 239820 182420 239876
rect 341292 239820 341348 239876
rect 186284 239708 186340 239764
rect 344988 239708 345044 239764
rect 187292 239596 187348 239652
rect 341068 239596 341124 239652
rect 358764 239484 358820 239540
rect 304892 239372 304948 239428
rect 314972 239372 315028 239428
rect 184380 239260 184436 239316
rect 272748 239260 272804 239316
rect 288204 239260 288260 239316
rect 314860 239148 314916 239204
rect 317436 239036 317492 239092
rect 341068 238588 341124 238644
rect 345772 238588 345828 238644
rect 349244 238588 349300 238644
rect 72940 238476 72996 238532
rect 76972 238476 77028 238532
rect 241948 238476 242004 238532
rect 242620 238476 242676 238532
rect 321244 238476 321300 238532
rect 321916 238476 321972 238532
rect 267260 238364 267316 238420
rect 96572 238252 96628 238308
rect 97020 238252 97076 238308
rect 356972 238140 357028 238196
rect 341964 237692 342020 237748
rect 233212 237244 233268 237300
rect 235900 237244 235956 237300
rect 219996 237020 220052 237076
rect 268716 237020 268772 237076
rect 270284 237020 270340 237076
rect 293916 237020 293972 237076
rect 218316 236908 218372 236964
rect 228508 236908 228564 236964
rect 236796 236908 236852 236964
rect 268604 236908 268660 236964
rect 270396 236908 270452 236964
rect 293804 236908 293860 236964
rect 295596 236908 295652 236964
rect 298956 236908 299012 236964
rect 300636 236908 300692 236964
rect 306572 236572 306628 236628
rect 46956 236124 47012 236180
rect 46172 236012 46228 236068
rect 307356 236012 307412 236068
rect 197596 235900 197652 235956
rect 359660 235900 359716 235956
rect 267484 235116 267540 235172
rect 340172 235116 340228 235172
rect 356748 235116 356804 235172
rect 266812 235004 266868 235060
rect 51772 234556 51828 234612
rect 269276 234556 269332 234612
rect 50204 234444 50260 234500
rect 315196 234444 315252 234500
rect 356748 234444 356804 234500
rect 267148 234332 267204 234388
rect 267372 234220 267428 234276
rect 590716 231868 590772 231924
rect 269612 231644 269668 231700
rect 312396 231644 312452 231700
rect 337372 231644 337428 231700
rect 311724 231532 311780 231588
rect 337148 231532 337204 231588
rect 340284 231420 340340 231476
rect 311948 231308 312004 231364
rect 320012 231196 320068 231252
rect 329196 231084 329252 231140
rect 267596 230860 267652 230916
rect 357980 230188 358036 230244
rect 358764 230188 358820 230244
rect 309932 229516 309988 229572
rect 338940 229516 338996 229572
rect 306796 229404 306852 229460
rect 339836 229292 339892 229348
rect 270732 228396 270788 228452
rect 270620 227500 270676 227556
rect 304892 226492 304948 226548
rect 338380 226380 338436 226436
rect 337260 226268 337316 226324
rect 338716 226156 338772 226212
rect 351372 225932 351428 225988
rect 48636 224476 48692 224532
rect 336588 224364 336644 224420
rect 51996 224252 52052 224308
rect 269500 224140 269556 224196
rect 336812 222796 336868 222852
rect 341628 222572 341684 222628
rect 187740 221116 187796 221172
rect 274092 221116 274148 221172
rect 356860 220668 356916 220724
rect 118412 220220 118468 220276
rect 181244 219772 181300 219828
rect 272524 219772 272580 219828
rect 338604 219772 338660 219828
rect 177884 219660 177940 219716
rect 272860 219660 272916 219716
rect 338828 219660 338884 219716
rect 199500 219548 199556 219604
rect 577052 218540 577108 218596
rect 186844 218092 186900 218148
rect 271068 218092 271124 218148
rect 186956 217980 187012 218036
rect 275884 217980 275940 218036
rect 4284 217644 4340 217700
rect 138572 217644 138628 217700
rect 172172 217644 172228 217700
rect 51884 217532 51940 217588
rect 187628 216524 187684 216580
rect 270956 216524 271012 216580
rect 187516 216412 187572 216468
rect 275772 216412 275828 216468
rect 199612 216300 199668 216356
rect 199724 216188 199780 216244
rect 307468 216188 307524 216244
rect 190876 216076 190932 216132
rect 359660 216076 359716 216132
rect 50316 215964 50372 216020
rect 274652 215852 274708 215908
rect 182924 214732 182980 214788
rect 272188 214732 272244 214788
rect 199388 214620 199444 214676
rect 194236 214508 194292 214564
rect 346556 214508 346612 214564
rect 34972 214284 35028 214340
rect 298172 214060 298228 214116
rect 184492 213164 184548 213220
rect 272412 213164 272468 213220
rect 179676 212940 179732 212996
rect 272972 212940 273028 212996
rect 174524 212828 174580 212884
rect 272300 212828 272356 212884
rect 4620 212716 4676 212772
rect 120092 212716 120148 212772
rect 174412 212716 174468 212772
rect 273420 212716 273476 212772
rect 4396 212604 4452 212660
rect 167132 212604 167188 212660
rect 39676 212492 39732 212548
rect 49644 211708 49700 211764
rect 273980 211708 274036 211764
rect 308252 211372 308308 211428
rect 272412 211260 272468 211316
rect 185724 211148 185780 211204
rect 272636 211148 272692 211204
rect 4508 211036 4564 211092
rect 113372 211036 113428 211092
rect 177996 211036 178052 211092
rect 272412 211036 272468 211092
rect 4172 210924 4228 210980
rect 121772 210924 121828 210980
rect 272188 210924 272244 210980
rect 174300 210476 174356 210532
rect 273196 210476 273252 210532
rect 49532 210028 49588 210084
rect 272636 209916 272692 209972
rect 349692 209916 349748 209972
rect 190428 209804 190484 209860
rect 185836 209692 185892 209748
rect 273084 209692 273140 209748
rect 174636 209580 174692 209636
rect 272188 209580 272244 209636
rect 181356 209356 181412 209412
rect 349804 209356 349860 209412
rect 359884 209244 359940 209300
rect 272524 209132 272580 209188
rect 269164 208684 269220 208740
rect 272300 207004 272356 207060
rect 4172 206332 4228 206388
rect 359884 205996 359940 206052
rect 350812 205884 350868 205940
rect 273308 205772 273364 205828
rect 359884 205772 359940 205828
rect 272188 204092 272244 204148
rect 342972 201516 343028 201572
rect 273420 201180 273476 201236
rect 272860 198268 272916 198324
rect 345996 198156 346052 198212
rect 336700 197932 336756 197988
rect 358988 197932 359044 197988
rect 317212 197820 317268 197876
rect 317324 197708 317380 197764
rect 315308 197596 315364 197652
rect 340060 197596 340116 197652
rect 344988 197484 345044 197540
rect 359324 197484 359380 197540
rect 270284 197372 270340 197428
rect 338156 197260 338212 197316
rect 339612 197036 339668 197092
rect 356076 197036 356132 197092
rect 345660 196700 345716 196756
rect 345548 196588 345604 196644
rect 352604 196588 352660 196644
rect 344204 196140 344260 196196
rect 359772 196140 359828 196196
rect 345548 195916 345604 195972
rect 344204 195692 344260 195748
rect 272972 195356 273028 195412
rect 345100 194908 345156 194964
rect 346444 194908 346500 194964
rect 345772 194796 345828 194852
rect 313404 194684 313460 194740
rect 336028 194684 336084 194740
rect 351036 194572 351092 194628
rect 349580 193228 349636 193284
rect 272748 192444 272804 192500
rect 346444 192444 346500 192500
rect 590828 192108 590884 192164
rect 351036 191772 351092 191828
rect 351148 191660 351204 191716
rect 359772 191604 359828 191660
rect 351260 191548 351316 191604
rect 272524 189532 272580 189588
rect 273196 186620 273252 186676
rect 359884 186172 359940 186228
rect 359884 185948 359940 186004
rect 356972 183820 357028 183876
rect 273084 183708 273140 183764
rect 356748 181356 356804 181412
rect 359772 181356 359828 181412
rect 356972 181132 357028 181188
rect 570332 178892 570388 178948
rect 4508 177996 4564 178052
rect 350700 177996 350756 178052
rect 359772 177996 359828 178052
rect 356972 175756 357028 175812
rect 346556 175420 346612 175476
rect 590716 175420 590772 175476
rect 356972 175308 357028 175364
rect 361452 175308 361508 175364
rect 590492 175308 590548 175364
rect 375228 175196 375284 175252
rect 352716 175084 352772 175140
rect 358428 174636 358484 174692
rect 417564 174636 417620 174692
rect 361676 174524 361732 174580
rect 362124 174412 362180 174468
rect 359436 173964 359492 174020
rect 355180 173516 355236 173572
rect 590604 173516 590660 173572
rect 559468 172956 559524 173012
rect 559580 172620 559636 172676
rect 360332 172172 360388 172228
rect 559468 172172 559524 172228
rect 360556 172060 360612 172116
rect 358540 171164 358596 171220
rect 355964 170716 356020 170772
rect 457772 170716 457828 170772
rect 359100 170492 359156 170548
rect 355852 169260 355908 169316
rect 457884 169260 457940 169316
rect 274092 169148 274148 169204
rect 352380 168924 352436 168980
rect 559804 168924 559860 168980
rect 354060 168812 354116 168868
rect 563164 168812 563220 168868
rect 354396 167916 354452 167972
rect 590828 167916 590884 167972
rect 350476 167244 350532 167300
rect 562828 167244 562884 167300
rect 559916 167132 559972 167188
rect 346668 167020 346724 167076
rect 357644 166348 357700 166404
rect 275884 166236 275940 166292
rect 352268 165564 352324 165620
rect 563052 165564 563108 165620
rect 359660 165452 359716 165508
rect 590604 165452 590660 165508
rect 349692 165004 349748 165060
rect 357084 164892 357140 164948
rect 357308 164780 357364 164836
rect 356972 164556 357028 164612
rect 357532 164556 357588 164612
rect 4172 163996 4228 164052
rect 355628 163996 355684 164052
rect 563388 163996 563444 164052
rect 346444 163884 346500 163940
rect 559692 163884 559748 163940
rect 346780 163772 346836 163828
rect 562940 163772 562996 163828
rect 271068 163324 271124 163380
rect 356972 163100 357028 163156
rect 357756 162988 357812 163044
rect 361676 162540 361732 162596
rect 352492 162428 352548 162484
rect 457996 162428 458052 162484
rect 350364 162204 350420 162260
rect 563276 162204 563332 162260
rect 270396 161756 270452 161812
rect 313404 160636 313460 160692
rect 314860 160076 314916 160132
rect 317436 160076 317492 160132
rect 346220 159740 346276 159796
rect 351372 159516 351428 159572
rect 324380 157836 324436 157892
rect 330652 157836 330708 157892
rect 332220 157836 332276 157892
rect 317324 157724 317380 157780
rect 273868 157500 273924 157556
rect 317100 157500 317156 157556
rect 346220 157052 346276 157108
rect 270956 154588 271012 154644
rect 275436 154476 275492 154532
rect 356188 154476 356244 154532
rect 357196 154476 357252 154532
rect 273980 154252 274036 154308
rect 275436 154252 275492 154308
rect 357756 153804 357812 153860
rect 490588 154252 490644 154308
rect 488908 154028 488964 154084
rect 272524 153580 272580 153636
rect 493164 153244 493220 153300
rect 502572 152908 502628 152964
rect 503132 152908 503188 152964
rect 353948 152684 354004 152740
rect 563612 152684 563668 152740
rect 348572 152572 348628 152628
rect 563724 152572 563780 152628
rect 278908 151676 278964 151732
rect 352940 151116 352996 151172
rect 348684 150444 348740 150500
rect 563500 150444 563556 150500
rect 506828 150220 506884 150276
rect 463372 149772 463428 149828
rect 482076 149660 482132 149716
rect 501004 149100 501060 149156
rect 501452 149100 501508 149156
rect 506828 149100 506884 149156
rect 462028 148988 462084 149044
rect 275772 148764 275828 148820
rect 348796 148764 348852 148820
rect 457996 148540 458052 148596
rect 357644 146972 357700 147028
rect 307356 145404 307412 145460
rect 358988 145068 359044 145124
rect 354284 142156 354340 142212
rect 356972 141932 357028 141988
rect 269388 140028 269444 140084
rect 356076 139244 356132 139300
rect 575372 139244 575428 139300
rect 357084 138572 357140 138628
rect 354172 136332 354228 136388
rect 4620 135772 4676 135828
rect 352156 133420 352212 133476
rect 357308 131964 357364 132020
rect 355740 131852 355796 131908
rect 457660 131852 457716 131908
rect 457660 130508 457716 130564
rect 348460 128492 348516 128548
rect 458108 128492 458164 128548
rect 356748 127596 356804 127652
rect 358876 126924 358932 126980
rect 458220 126924 458276 126980
rect 350588 126812 350644 126868
rect 457996 126812 458052 126868
rect 561260 125692 561316 125748
rect 352604 124684 352660 124740
rect 384860 122668 384916 122724
rect 386876 122668 386932 122724
rect 388892 122668 388948 122724
rect 390908 122668 390964 122724
rect 394940 122668 394996 122724
rect 411628 122668 411684 122724
rect 414988 122668 415044 122724
rect 346892 121884 346948 121940
rect 457660 121884 457716 121940
rect 349132 121772 349188 121828
rect 566188 120988 566244 121044
rect 359324 120428 359380 120484
rect 421708 120428 421764 120484
rect 352044 120092 352100 120148
rect 458332 120092 458388 120148
rect 457660 118860 457716 118916
rect 359996 118748 360052 118804
rect 421820 118748 421876 118804
rect 362012 118636 362068 118692
rect 458556 118636 458612 118692
rect 361788 118524 361844 118580
rect 457660 118524 457716 118580
rect 355516 118412 355572 118468
rect 457548 118412 457604 118468
rect 458556 117516 458612 117572
rect 360444 117068 360500 117124
rect 458332 117068 458388 117124
rect 359548 116956 359604 117012
rect 457660 116844 457716 116900
rect 458444 116844 458500 116900
rect 564732 116284 564788 116340
rect 421708 116060 421764 116116
rect 425852 116060 425908 116116
rect 457660 115836 457716 115892
rect 312060 113820 312116 113876
rect 564620 113148 564676 113204
rect 590604 113036 590660 113092
rect 273308 110908 273364 110964
rect 564508 110012 564564 110068
rect 421820 109116 421876 109172
rect 424172 109116 424228 109172
rect 311948 107996 312004 108052
rect 563164 106876 563220 106932
rect 561148 105308 561204 105364
rect 563388 103740 563444 103796
rect 563276 102172 563332 102228
rect 563052 100604 563108 100660
rect 585452 99820 585508 99876
rect 563724 99036 563780 99092
rect 458556 98476 458612 98532
rect 562940 97468 562996 97524
rect 559916 95900 559972 95956
rect 457660 95564 457716 95620
rect 563612 94332 563668 94388
rect 4396 93436 4452 93492
rect 562828 92764 562884 92820
rect 563500 91196 563556 91252
rect 279692 90524 279748 90580
rect 458444 89740 458500 89796
rect 559804 89628 559860 89684
rect 315196 87612 315252 87668
rect 458332 86828 458388 86884
rect 350252 84924 350308 84980
rect 559804 84924 559860 84980
rect 330092 84700 330148 84756
rect 457884 83916 457940 83972
rect 562828 83356 562884 83412
rect 457772 81004 457828 81060
rect 559580 78652 559636 78708
rect 458220 78092 458276 78148
rect 559692 77084 559748 77140
rect 559468 75516 559524 75572
rect 458108 75180 458164 75236
rect 562940 73948 562996 74004
rect 590492 73388 590548 73444
rect 457996 72156 458052 72212
rect 457772 69244 457828 69300
rect 424172 66332 424228 66388
rect 457660 66332 457716 66388
rect 457884 66332 457940 66388
rect 563052 66108 563108 66164
rect 563164 64540 563220 64596
rect 457996 63420 458052 63476
rect 425852 60620 425908 60676
rect 573692 59948 573748 60004
rect 457660 57708 457716 57764
rect 559468 56028 559524 56084
rect 457660 54684 457716 54740
rect 355404 52892 355460 52948
rect 457996 52892 458052 52948
rect 358652 52668 358708 52724
rect 457772 52668 457828 52724
rect 289772 51996 289828 52052
rect 457660 51996 457716 52052
rect 353836 51436 353892 51492
rect 457884 51436 457940 51492
rect 4284 51100 4340 51156
rect 307468 50316 307524 50372
rect 315308 50316 315364 50372
rect 559468 50204 559524 50260
rect 351932 50092 351988 50148
rect 563052 50092 563108 50148
rect 353724 49980 353780 50036
rect 562940 49980 562996 50036
rect 269500 49644 269556 49700
rect 46956 49532 47012 49588
rect 269836 49532 269892 49588
rect 267148 48748 267204 48804
rect 315084 48524 315140 48580
rect 267596 48412 267652 48468
rect 48524 48188 48580 48244
rect 51772 48076 51828 48132
rect 270844 48076 270900 48132
rect 355292 48076 355348 48132
rect 563164 48076 563220 48132
rect 50204 47964 50260 48020
rect 269276 47964 269332 48020
rect 349244 47964 349300 48020
rect 267372 45276 267428 45332
rect 349356 45276 349412 45332
rect 267484 45164 267540 45220
rect 353612 45164 353668 45220
rect 562828 45164 562884 45220
rect 266812 45052 266868 45108
rect 359772 45052 359828 45108
rect 559804 45052 559860 45108
rect 269612 44716 269668 44772
rect 269724 44492 269780 44548
rect 270732 41244 270788 41300
rect 270508 41132 270564 41188
rect 270620 37996 270676 38052
rect 311612 37884 311668 37940
rect 311836 37772 311892 37828
rect 309932 27692 309988 27748
rect 275660 26012 275716 26068
rect 274652 24556 274708 24612
rect 572012 20300 572068 20356
rect 267260 17612 267316 17668
rect 4172 8764 4228 8820
rect 275548 7532 275604 7588
rect 288092 7084 288148 7140
rect 51884 4956 51940 5012
rect 41356 4844 41412 4900
rect 50316 4732 50372 4788
rect 285180 4732 285236 4788
rect 209132 4620 209188 4676
rect 283052 4508 283108 4564
rect 281372 4396 281428 4452
rect 35196 4284 35252 4340
rect 51996 4284 52052 4340
rect 284956 4284 285012 4340
rect 16716 4172 16772 4228
rect 18396 4172 18452 4228
rect 20076 4172 20132 4228
rect 25116 4172 25172 4228
rect 35084 4172 35140 4228
rect 48636 4172 48692 4228
rect 579628 4172 579684 4228
rect 581308 4172 581364 4228
rect 582988 4172 583044 4228
rect 172956 4060 173012 4116
rect 55132 3388 55188 3444
rect 60844 3388 60900 3444
rect 91532 3388 91588 3444
rect 142940 3388 142996 3444
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect 5418 580350 6038 596784
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect 5418 562350 6038 579922
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect 4172 558964 4228 558974
rect 4172 469588 4228 558908
rect 5418 544350 6038 561922
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect 5418 526350 6038 543922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect 4172 469522 4228 469532
rect 4284 516628 4340 516638
rect 4284 467908 4340 516572
rect 5418 508350 6038 525922
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect 5418 490350 6038 507922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 4284 467842 4340 467852
rect 4396 474292 4452 474302
rect 4396 466228 4452 474236
rect 4396 466162 4452 466172
rect 5418 472350 6038 489922
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect 5418 454350 6038 471922
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect 5418 436350 6038 453922
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect 5418 418350 6038 435922
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect 5418 400350 6038 417922
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect 4396 389620 4452 389630
rect 4396 377188 4452 389564
rect 4396 377122 4452 377132
rect 5418 382350 6038 399922
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect 4172 376318 4228 376328
rect 4172 375732 4228 376262
rect 4172 375666 4228 375676
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect 5418 364350 6038 381922
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect 4172 347284 4228 347294
rect 4172 306628 4228 347228
rect 4172 306562 4228 306572
rect 5418 346350 6038 363922
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect 5418 328350 6038 345922
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect 5418 310350 6038 327922
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect 4172 296660 4228 296670
rect 4172 262836 4228 296604
rect 4172 262770 4228 262780
rect 5418 292350 6038 309922
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect 5418 274350 6038 291922
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect 5418 256350 6038 273922
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 4172 248500 4228 248510
rect 4172 247078 4228 248444
rect 4172 247012 4228 247022
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect 5418 238350 6038 255922
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect 5418 220350 6038 237922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect 4284 217700 4340 217710
rect 4172 210980 4228 210990
rect 4172 208348 4228 210924
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect 4060 208292 4228 208348
rect 4060 196588 4116 208292
rect 4172 206578 4228 206588
rect 4172 206388 4228 206522
rect 4172 206322 4228 206332
rect 4060 196532 4228 196588
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect 4172 173068 4228 196532
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect 4060 173012 4228 173068
rect 4060 161308 4116 173012
rect 4172 164638 4228 164648
rect 4172 164052 4228 164582
rect 4172 163986 4228 163996
rect 4060 161252 4228 161308
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect 4172 8820 4228 161252
rect 4284 51156 4340 217644
rect 4620 212772 4676 212782
rect 4396 212660 4452 212670
rect 4396 93492 4452 212604
rect 4508 211092 4564 211102
rect 4508 178052 4564 211036
rect 4508 177986 4564 177996
rect 4620 135828 4676 212716
rect 4620 135762 4676 135772
rect 5418 202350 6038 219922
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect 5418 184350 6038 201922
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 5418 166350 6038 183922
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect 5418 148350 6038 165922
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 4396 93426 4452 93436
rect 5418 130350 6038 147922
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect 5418 112350 6038 129922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect 5418 94350 6038 111922
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 4284 51090 4340 51100
rect 5418 76350 6038 93922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 5418 58350 6038 75922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 4172 8754 4228 8764
rect 5418 40350 6038 57922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect 5418 22350 6038 39922
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 4350 6038 21922
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 9138 568350 9758 585922
rect 9138 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 9758 568350
rect 9138 568226 9758 568294
rect 9138 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 9758 568226
rect 9138 568102 9758 568170
rect 9138 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 9758 568102
rect 9138 567978 9758 568046
rect 9138 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 9758 567978
rect 9138 550350 9758 567922
rect 9138 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 9758 550350
rect 9138 550226 9758 550294
rect 9138 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 9758 550226
rect 9138 550102 9758 550170
rect 9138 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 9758 550102
rect 9138 549978 9758 550046
rect 9138 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 9758 549978
rect 9138 532350 9758 549922
rect 9138 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 9758 532350
rect 9138 532226 9758 532294
rect 9138 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 9758 532226
rect 9138 532102 9758 532170
rect 9138 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 9758 532102
rect 9138 531978 9758 532046
rect 9138 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 9758 531978
rect 9138 514350 9758 531922
rect 9138 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 9758 514350
rect 9138 514226 9758 514294
rect 9138 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 9758 514226
rect 9138 514102 9758 514170
rect 9138 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 9758 514102
rect 9138 513978 9758 514046
rect 9138 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 9758 513978
rect 9138 496350 9758 513922
rect 9138 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 9758 496350
rect 9138 496226 9758 496294
rect 9138 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 9758 496226
rect 9138 496102 9758 496170
rect 9138 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 9758 496102
rect 9138 495978 9758 496046
rect 9138 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 9758 495978
rect 9138 478350 9758 495922
rect 9138 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 9758 478350
rect 9138 478226 9758 478294
rect 9138 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 9758 478226
rect 9138 478102 9758 478170
rect 9138 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 9758 478102
rect 9138 477978 9758 478046
rect 9138 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 9758 477978
rect 9138 460350 9758 477922
rect 9138 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 9758 460350
rect 9138 460226 9758 460294
rect 9138 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 9758 460226
rect 9138 460102 9758 460170
rect 9138 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 9758 460102
rect 9138 459978 9758 460046
rect 9138 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 9758 459978
rect 9138 442350 9758 459922
rect 9138 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 9758 442350
rect 9138 442226 9758 442294
rect 9138 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 9758 442226
rect 9138 442102 9758 442170
rect 9138 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 9758 442102
rect 9138 441978 9758 442046
rect 9138 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 9758 441978
rect 9138 424350 9758 441922
rect 9138 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 9758 424350
rect 9138 424226 9758 424294
rect 9138 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 9758 424226
rect 9138 424102 9758 424170
rect 9138 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 9758 424102
rect 9138 423978 9758 424046
rect 9138 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 9758 423978
rect 9138 406350 9758 423922
rect 9138 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 9758 406350
rect 9138 406226 9758 406294
rect 9138 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 9758 406226
rect 9138 406102 9758 406170
rect 9138 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 9758 406102
rect 9138 405978 9758 406046
rect 9138 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 9758 405978
rect 9138 388350 9758 405922
rect 9138 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 9758 388350
rect 9138 388226 9758 388294
rect 9138 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 9758 388226
rect 9138 388102 9758 388170
rect 9138 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 9758 388102
rect 9138 387978 9758 388046
rect 9138 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 9758 387978
rect 9138 370350 9758 387922
rect 9138 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 9758 370350
rect 9138 370226 9758 370294
rect 9138 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 9758 370226
rect 9138 370102 9758 370170
rect 9138 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 9758 370102
rect 9138 369978 9758 370046
rect 9138 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 9758 369978
rect 9138 352350 9758 369922
rect 9138 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 9758 352350
rect 9138 352226 9758 352294
rect 9138 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 9758 352226
rect 9138 352102 9758 352170
rect 9138 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 9758 352102
rect 9138 351978 9758 352046
rect 9138 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 9758 351978
rect 9138 334350 9758 351922
rect 9138 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 9758 334350
rect 9138 334226 9758 334294
rect 9138 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 9758 334226
rect 9138 334102 9758 334170
rect 9138 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 9758 334102
rect 9138 333978 9758 334046
rect 9138 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 9758 333978
rect 9138 316350 9758 333922
rect 9138 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 9758 316350
rect 9138 316226 9758 316294
rect 9138 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 9758 316226
rect 9138 316102 9758 316170
rect 9138 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 9758 316102
rect 9138 315978 9758 316046
rect 9138 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 9758 315978
rect 9138 298350 9758 315922
rect 9138 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 9758 298350
rect 9138 298226 9758 298294
rect 9138 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 9758 298226
rect 9138 298102 9758 298170
rect 9138 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 9758 298102
rect 9138 297978 9758 298046
rect 9138 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 9758 297978
rect 9138 280350 9758 297922
rect 9138 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 9758 280350
rect 9138 280226 9758 280294
rect 9138 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 9758 280226
rect 9138 280102 9758 280170
rect 9138 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 9758 280102
rect 9138 279978 9758 280046
rect 9138 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 9758 279978
rect 9138 262350 9758 279922
rect 9138 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 9758 262350
rect 9138 262226 9758 262294
rect 9138 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 9758 262226
rect 9138 262102 9758 262170
rect 9138 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 9758 262102
rect 9138 261978 9758 262046
rect 9138 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 9758 261978
rect 9138 244350 9758 261922
rect 9138 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 9758 244350
rect 9138 244226 9758 244294
rect 9138 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 9758 244226
rect 9138 244102 9758 244170
rect 9138 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 9758 244102
rect 9138 243978 9758 244046
rect 9138 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 9758 243978
rect 9138 226350 9758 243922
rect 36138 597212 36758 598268
rect 36138 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 36758 597212
rect 36138 597088 36758 597156
rect 36138 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 36758 597088
rect 36138 596964 36758 597032
rect 36138 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 36758 596964
rect 36138 596840 36758 596908
rect 36138 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 36758 596840
rect 36138 580350 36758 596784
rect 36138 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 36758 580350
rect 36138 580226 36758 580294
rect 36138 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 36758 580226
rect 36138 580102 36758 580170
rect 36138 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 36758 580102
rect 36138 579978 36758 580046
rect 36138 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 36758 579978
rect 36138 562350 36758 579922
rect 36138 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 36758 562350
rect 36138 562226 36758 562294
rect 36138 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 36758 562226
rect 36138 562102 36758 562170
rect 36138 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 36758 562102
rect 36138 561978 36758 562046
rect 36138 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 36758 561978
rect 36138 544350 36758 561922
rect 36138 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 36758 544350
rect 36138 544226 36758 544294
rect 36138 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 36758 544226
rect 36138 544102 36758 544170
rect 36138 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 36758 544102
rect 36138 543978 36758 544046
rect 36138 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 36758 543978
rect 36138 526350 36758 543922
rect 36138 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 36758 526350
rect 36138 526226 36758 526294
rect 36138 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 36758 526226
rect 36138 526102 36758 526170
rect 36138 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 36758 526102
rect 36138 525978 36758 526046
rect 36138 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 36758 525978
rect 36138 508350 36758 525922
rect 36138 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 36758 508350
rect 36138 508226 36758 508294
rect 36138 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 36758 508226
rect 36138 508102 36758 508170
rect 36138 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 36758 508102
rect 36138 507978 36758 508046
rect 36138 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 36758 507978
rect 36138 490350 36758 507922
rect 36138 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 36758 490350
rect 36138 490226 36758 490294
rect 36138 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 36758 490226
rect 36138 490102 36758 490170
rect 36138 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 36758 490102
rect 36138 489978 36758 490046
rect 36138 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 36758 489978
rect 36138 472350 36758 489922
rect 36138 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 36758 472350
rect 36138 472226 36758 472294
rect 36138 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 36758 472226
rect 36138 472102 36758 472170
rect 36138 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 36758 472102
rect 36138 471978 36758 472046
rect 36138 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 36758 471978
rect 36138 454350 36758 471922
rect 36138 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 36758 454350
rect 36138 454226 36758 454294
rect 36138 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 36758 454226
rect 36138 454102 36758 454170
rect 36138 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 36758 454102
rect 36138 453978 36758 454046
rect 36138 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 36758 453978
rect 36138 436350 36758 453922
rect 36138 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 36758 436350
rect 36138 436226 36758 436294
rect 36138 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 36758 436226
rect 36138 436102 36758 436170
rect 36138 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 36758 436102
rect 36138 435978 36758 436046
rect 36138 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 36758 435978
rect 36138 418350 36758 435922
rect 36138 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 36758 418350
rect 36138 418226 36758 418294
rect 36138 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 36758 418226
rect 36138 418102 36758 418170
rect 36138 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 36758 418102
rect 36138 417978 36758 418046
rect 36138 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 36758 417978
rect 36138 400350 36758 417922
rect 36138 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 36758 400350
rect 36138 400226 36758 400294
rect 36138 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 36758 400226
rect 36138 400102 36758 400170
rect 36138 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 36758 400102
rect 36138 399978 36758 400046
rect 36138 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 36758 399978
rect 36138 382350 36758 399922
rect 36138 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 36758 382350
rect 36138 382226 36758 382294
rect 36138 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 36758 382226
rect 36138 382102 36758 382170
rect 36138 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 36758 382102
rect 36138 381978 36758 382046
rect 36138 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 36758 381978
rect 36138 364350 36758 381922
rect 36138 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 36758 364350
rect 36138 364226 36758 364294
rect 36138 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 36758 364226
rect 36138 364102 36758 364170
rect 36138 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 36758 364102
rect 36138 363978 36758 364046
rect 36138 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 36758 363978
rect 36138 346350 36758 363922
rect 36138 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 36758 346350
rect 36138 346226 36758 346294
rect 36138 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 36758 346226
rect 36138 346102 36758 346170
rect 36138 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 36758 346102
rect 36138 345978 36758 346046
rect 36138 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 36758 345978
rect 36138 328350 36758 345922
rect 36138 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 36758 328350
rect 36138 328226 36758 328294
rect 36138 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 36758 328226
rect 36138 328102 36758 328170
rect 36138 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 36758 328102
rect 36138 327978 36758 328046
rect 36138 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 36758 327978
rect 36138 310350 36758 327922
rect 36138 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 36758 310350
rect 36138 310226 36758 310294
rect 36138 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 36758 310226
rect 36138 310102 36758 310170
rect 36138 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 36758 310102
rect 36138 309978 36758 310046
rect 36138 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 36758 309978
rect 36138 292350 36758 309922
rect 36138 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 36758 292350
rect 36138 292226 36758 292294
rect 36138 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 36758 292226
rect 36138 292102 36758 292170
rect 36138 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 36758 292102
rect 36138 291978 36758 292046
rect 36138 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 36758 291978
rect 36138 274350 36758 291922
rect 36138 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 36758 274350
rect 36138 274226 36758 274294
rect 36138 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 36758 274226
rect 36138 274102 36758 274170
rect 36138 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 36758 274102
rect 36138 273978 36758 274046
rect 36138 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 36758 273978
rect 36138 256350 36758 273922
rect 36138 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 36758 256350
rect 36138 256226 36758 256294
rect 36138 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 36758 256226
rect 36138 256102 36758 256170
rect 36138 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 36758 256102
rect 36138 255978 36758 256046
rect 36138 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 36758 255978
rect 35196 241138 35252 241148
rect 9138 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 9758 226350
rect 9138 226226 9758 226294
rect 9138 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 9758 226226
rect 9138 226102 9758 226170
rect 9138 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 9758 226102
rect 9138 225978 9758 226046
rect 9138 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 9758 225978
rect 9138 208350 9758 225922
rect 9138 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 9758 208350
rect 9138 208226 9758 208294
rect 9138 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 9758 208226
rect 9138 208102 9758 208170
rect 9138 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 9758 208102
rect 9138 207978 9758 208046
rect 9138 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 9758 207978
rect 9138 190350 9758 207922
rect 9138 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 9758 190350
rect 9138 190226 9758 190294
rect 9138 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 9758 190226
rect 9138 190102 9758 190170
rect 9138 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 9758 190102
rect 9138 189978 9758 190046
rect 9138 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 9758 189978
rect 9138 172350 9758 189922
rect 9138 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 9758 172350
rect 9138 172226 9758 172294
rect 9138 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 9758 172226
rect 9138 172102 9758 172170
rect 9138 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 9758 172102
rect 9138 171978 9758 172046
rect 9138 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 9758 171978
rect 9138 154350 9758 171922
rect 9138 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 9758 154350
rect 9138 154226 9758 154294
rect 9138 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 9758 154226
rect 9138 154102 9758 154170
rect 9138 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 9758 154102
rect 9138 153978 9758 154046
rect 9138 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 9758 153978
rect 9138 136350 9758 153922
rect 9138 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 9758 136350
rect 9138 136226 9758 136294
rect 9138 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 9758 136226
rect 9138 136102 9758 136170
rect 9138 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 9758 136102
rect 9138 135978 9758 136046
rect 9138 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 9758 135978
rect 9138 118350 9758 135922
rect 9138 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 9758 118350
rect 9138 118226 9758 118294
rect 9138 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 9758 118226
rect 9138 118102 9758 118170
rect 9138 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 9758 118102
rect 9138 117978 9758 118046
rect 9138 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 9758 117978
rect 9138 100350 9758 117922
rect 9138 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 9758 100350
rect 9138 100226 9758 100294
rect 9138 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 9758 100226
rect 9138 100102 9758 100170
rect 9138 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 9758 100102
rect 9138 99978 9758 100046
rect 9138 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 9758 99978
rect 9138 82350 9758 99922
rect 9138 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 9758 82350
rect 9138 82226 9758 82294
rect 9138 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 9758 82226
rect 9138 82102 9758 82170
rect 9138 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 9758 82102
rect 9138 81978 9758 82046
rect 9138 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 9758 81978
rect 9138 64350 9758 81922
rect 9138 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 9758 64350
rect 9138 64226 9758 64294
rect 9138 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 9758 64226
rect 9138 64102 9758 64170
rect 9138 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 9758 64102
rect 9138 63978 9758 64046
rect 9138 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 9758 63978
rect 9138 46350 9758 63922
rect 9138 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 9758 46350
rect 9138 46226 9758 46294
rect 9138 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 9758 46226
rect 9138 46102 9758 46170
rect 9138 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 9758 46102
rect 9138 45978 9758 46046
rect 9138 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 9758 45978
rect 9138 28350 9758 45922
rect 9138 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 9758 28350
rect 9138 28226 9758 28294
rect 9138 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 9758 28226
rect 9138 28102 9758 28170
rect 9138 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 9758 28102
rect 9138 27978 9758 28046
rect 9138 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 9758 27978
rect 9138 10350 9758 27922
rect 9138 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 9758 10350
rect 9138 10226 9758 10294
rect 9138 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 9758 10226
rect 9138 10102 9758 10170
rect 9138 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 9758 10102
rect 9138 9978 9758 10046
rect 9138 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 9758 9978
rect 9138 -1120 9758 9922
rect 16716 234298 16772 234308
rect 16716 4228 16772 234242
rect 25116 231058 25172 231068
rect 16716 4162 16772 4172
rect 18396 227638 18452 227648
rect 18396 4228 18452 227582
rect 18396 4162 18452 4172
rect 20076 224218 20132 224228
rect 20076 4228 20132 224162
rect 20076 4162 20132 4172
rect 25116 4228 25172 231002
rect 35084 230338 35140 230348
rect 34972 214340 35028 214350
rect 34972 4798 35028 214284
rect 34972 4732 35028 4742
rect 25116 4162 25172 4172
rect 35084 4228 35140 230282
rect 35196 4340 35252 241082
rect 35196 4274 35252 4284
rect 36138 238350 36758 255922
rect 36138 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 36758 238350
rect 36138 238226 36758 238294
rect 36138 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 36758 238226
rect 36138 238102 36758 238170
rect 36138 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 36758 238102
rect 36138 237978 36758 238046
rect 36138 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 36758 237978
rect 36138 220350 36758 237922
rect 36138 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 36758 220350
rect 36138 220226 36758 220294
rect 36138 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 36758 220226
rect 36138 220102 36758 220170
rect 36138 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 36758 220102
rect 36138 219978 36758 220046
rect 36138 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 36758 219978
rect 36138 202350 36758 219922
rect 39858 598172 40478 598268
rect 39858 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 40478 598172
rect 39858 598048 40478 598116
rect 39858 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 40478 598048
rect 39858 597924 40478 597992
rect 39858 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 40478 597924
rect 39858 597800 40478 597868
rect 39858 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 40478 597800
rect 39858 586350 40478 597744
rect 39858 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 40478 586350
rect 39858 586226 40478 586294
rect 39858 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 40478 586226
rect 39858 586102 40478 586170
rect 39858 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 40478 586102
rect 39858 585978 40478 586046
rect 39858 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 40478 585978
rect 39858 568350 40478 585922
rect 39858 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 40478 568350
rect 39858 568226 40478 568294
rect 39858 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 40478 568226
rect 39858 568102 40478 568170
rect 39858 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 40478 568102
rect 39858 567978 40478 568046
rect 39858 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 40478 567978
rect 39858 550350 40478 567922
rect 39858 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 40478 550350
rect 39858 550226 40478 550294
rect 39858 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 40478 550226
rect 39858 550102 40478 550170
rect 39858 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 40478 550102
rect 39858 549978 40478 550046
rect 39858 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 40478 549978
rect 39858 532350 40478 549922
rect 39858 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532294 40478 532350
rect 39858 532226 40478 532294
rect 39858 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 40478 532226
rect 39858 532102 40478 532170
rect 39858 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 40478 532102
rect 39858 531978 40478 532046
rect 39858 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 40478 531978
rect 39858 514350 40478 531922
rect 66858 597212 67478 598268
rect 66858 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 67478 597212
rect 66858 597088 67478 597156
rect 66858 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 67478 597088
rect 66858 596964 67478 597032
rect 66858 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 67478 596964
rect 66858 596840 67478 596908
rect 66858 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 67478 596840
rect 66858 580350 67478 596784
rect 66858 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 67478 580350
rect 66858 580226 67478 580294
rect 66858 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 67478 580226
rect 66858 580102 67478 580170
rect 66858 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 67478 580102
rect 66858 579978 67478 580046
rect 66858 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 67478 579978
rect 66858 562350 67478 579922
rect 66858 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 67478 562350
rect 66858 562226 67478 562294
rect 66858 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 67478 562226
rect 66858 562102 67478 562170
rect 66858 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 67478 562102
rect 66858 561978 67478 562046
rect 66858 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 67478 561978
rect 66858 544350 67478 561922
rect 66858 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 67478 544350
rect 66858 544226 67478 544294
rect 66858 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 67478 544226
rect 66858 544102 67478 544170
rect 66858 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 67478 544102
rect 66858 543978 67478 544046
rect 66858 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 67478 543978
rect 66858 530232 67478 543922
rect 70578 598172 71198 598268
rect 70578 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 71198 598172
rect 70578 598048 71198 598116
rect 70578 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 71198 598048
rect 70578 597924 71198 597992
rect 70578 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 71198 597924
rect 70578 597800 71198 597868
rect 70578 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 71198 597800
rect 70578 586350 71198 597744
rect 70578 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 71198 586350
rect 70578 586226 71198 586294
rect 70578 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 71198 586226
rect 70578 586102 71198 586170
rect 70578 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 71198 586102
rect 70578 585978 71198 586046
rect 70578 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 71198 585978
rect 70578 568350 71198 585922
rect 70578 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 71198 568350
rect 70578 568226 71198 568294
rect 70578 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 71198 568226
rect 70578 568102 71198 568170
rect 70578 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 71198 568102
rect 70578 567978 71198 568046
rect 70578 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 71198 567978
rect 70578 550350 71198 567922
rect 70578 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 71198 550350
rect 70578 550226 71198 550294
rect 70578 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 71198 550226
rect 70578 550102 71198 550170
rect 70578 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 71198 550102
rect 70578 549978 71198 550046
rect 70578 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 71198 549978
rect 70578 533912 71198 549922
rect 97578 597212 98198 598268
rect 97578 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 98198 597212
rect 97578 597088 98198 597156
rect 97578 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 98198 597088
rect 97578 596964 98198 597032
rect 97578 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 98198 596964
rect 97578 596840 98198 596908
rect 97578 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 98198 596840
rect 97578 580350 98198 596784
rect 97578 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 98198 580350
rect 97578 580226 98198 580294
rect 97578 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 98198 580226
rect 97578 580102 98198 580170
rect 97578 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 98198 580102
rect 97578 579978 98198 580046
rect 97578 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 98198 579978
rect 97578 562350 98198 579922
rect 97578 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 98198 562350
rect 97578 562226 98198 562294
rect 97578 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 98198 562226
rect 97578 562102 98198 562170
rect 97578 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 98198 562102
rect 97578 561978 98198 562046
rect 97578 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 98198 561978
rect 97578 544350 98198 561922
rect 97578 544294 97674 544350
rect 97730 544294 97798 544350
rect 97854 544294 97922 544350
rect 97978 544294 98046 544350
rect 98102 544294 98198 544350
rect 97578 544226 98198 544294
rect 97578 544170 97674 544226
rect 97730 544170 97798 544226
rect 97854 544170 97922 544226
rect 97978 544170 98046 544226
rect 98102 544170 98198 544226
rect 97578 544102 98198 544170
rect 97578 544046 97674 544102
rect 97730 544046 97798 544102
rect 97854 544046 97922 544102
rect 97978 544046 98046 544102
rect 98102 544046 98198 544102
rect 97578 543978 98198 544046
rect 97578 543922 97674 543978
rect 97730 543922 97798 543978
rect 97854 543922 97922 543978
rect 97978 543922 98046 543978
rect 98102 543922 98198 543978
rect 97578 541432 98198 543922
rect 101298 598172 101918 598268
rect 101298 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 101918 598172
rect 101298 598048 101918 598116
rect 101298 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 101918 598048
rect 101298 597924 101918 597992
rect 101298 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 101918 597924
rect 101298 597800 101918 597868
rect 101298 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 101918 597800
rect 101298 586350 101918 597744
rect 101298 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 101918 586350
rect 101298 586226 101918 586294
rect 101298 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 101918 586226
rect 101298 586102 101918 586170
rect 101298 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 101918 586102
rect 101298 585978 101918 586046
rect 101298 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 101918 585978
rect 101298 568350 101918 585922
rect 101298 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 101918 568350
rect 101298 568226 101918 568294
rect 101298 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 101918 568226
rect 101298 568102 101918 568170
rect 101298 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 101918 568102
rect 101298 567978 101918 568046
rect 101298 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 101918 567978
rect 101298 550350 101918 567922
rect 128298 597212 128918 598268
rect 128298 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 128918 597212
rect 128298 597088 128918 597156
rect 128298 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 128918 597088
rect 128298 596964 128918 597032
rect 128298 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 128918 596964
rect 128298 596840 128918 596908
rect 128298 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 128918 596840
rect 128298 580350 128918 596784
rect 128298 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 128918 580350
rect 128298 580226 128918 580294
rect 128298 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 128918 580226
rect 128298 580102 128918 580170
rect 128298 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 128918 580102
rect 128298 579978 128918 580046
rect 128298 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 128918 579978
rect 128298 562350 128918 579922
rect 128298 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 128918 562350
rect 128298 562226 128918 562294
rect 128298 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 128918 562226
rect 128298 562102 128918 562170
rect 128298 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 128918 562102
rect 117280 561988 124640 562040
rect 117280 561932 117336 561988
rect 117392 561932 117460 561988
rect 117516 561932 117584 561988
rect 117640 561932 117708 561988
rect 117764 561932 117832 561988
rect 117888 561932 117956 561988
rect 118012 561932 118080 561988
rect 118136 561932 118204 561988
rect 118260 561932 118328 561988
rect 118384 561932 118452 561988
rect 118508 561932 118576 561988
rect 118632 561932 118700 561988
rect 118756 561932 118824 561988
rect 118880 561932 118948 561988
rect 119004 561932 119072 561988
rect 119128 561932 119196 561988
rect 119252 561932 119320 561988
rect 119376 561932 119444 561988
rect 119500 561932 119568 561988
rect 119624 561932 119692 561988
rect 119748 561932 119816 561988
rect 119872 561932 119940 561988
rect 119996 561932 120064 561988
rect 120120 561932 120188 561988
rect 120244 561932 120312 561988
rect 120368 561932 120436 561988
rect 120492 561932 120560 561988
rect 120616 561932 120684 561988
rect 120740 561932 120808 561988
rect 120864 561932 120932 561988
rect 120988 561932 121056 561988
rect 121112 561932 121180 561988
rect 121236 561932 121304 561988
rect 121360 561932 121428 561988
rect 121484 561932 121552 561988
rect 121608 561932 121676 561988
rect 121732 561932 121800 561988
rect 121856 561932 121924 561988
rect 121980 561932 122048 561988
rect 122104 561932 122172 561988
rect 122228 561932 122296 561988
rect 122352 561932 122420 561988
rect 122476 561932 122544 561988
rect 122600 561932 122668 561988
rect 122724 561932 122792 561988
rect 122848 561932 122916 561988
rect 122972 561932 123040 561988
rect 123096 561932 123164 561988
rect 123220 561932 123288 561988
rect 123344 561932 123412 561988
rect 123468 561932 123536 561988
rect 123592 561932 123660 561988
rect 123716 561932 123784 561988
rect 123840 561932 123908 561988
rect 123964 561932 124032 561988
rect 124088 561932 124156 561988
rect 124212 561932 124280 561988
rect 124336 561932 124404 561988
rect 124460 561932 124528 561988
rect 124584 561932 124640 561988
rect 117280 561880 124640 561932
rect 128298 561978 128918 562046
rect 128298 561922 128394 561978
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 128918 561978
rect 101298 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 101918 550350
rect 101298 550226 101918 550294
rect 101298 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 101918 550226
rect 101298 550102 101918 550170
rect 101298 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 101918 550102
rect 101298 549978 101918 550046
rect 101298 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 101918 549978
rect 101298 542872 101918 549922
rect 128298 544350 128918 561922
rect 128298 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 128918 544350
rect 128298 544226 128918 544294
rect 128298 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 128918 544226
rect 104000 544063 121920 544120
rect 104000 544007 104066 544063
rect 104122 544007 104190 544063
rect 104246 544007 104314 544063
rect 104370 544007 104438 544063
rect 104494 544007 104562 544063
rect 104618 544007 104686 544063
rect 104742 544007 104810 544063
rect 104866 544007 104934 544063
rect 104990 544007 105058 544063
rect 105114 544007 105182 544063
rect 105238 544007 105306 544063
rect 105362 544007 105430 544063
rect 105486 544007 105554 544063
rect 105610 544007 105678 544063
rect 105734 544007 105802 544063
rect 105858 544007 105926 544063
rect 105982 544007 106050 544063
rect 106106 544007 106174 544063
rect 106230 544007 106298 544063
rect 106354 544007 106422 544063
rect 106478 544007 106546 544063
rect 106602 544007 106670 544063
rect 106726 544007 106794 544063
rect 106850 544007 106918 544063
rect 106974 544007 107042 544063
rect 107098 544007 107166 544063
rect 107222 544007 107290 544063
rect 107346 544007 107414 544063
rect 107470 544007 107538 544063
rect 107594 544007 107662 544063
rect 107718 544007 107786 544063
rect 107842 544007 107910 544063
rect 107966 544007 108034 544063
rect 108090 544007 108158 544063
rect 108214 544007 108282 544063
rect 108338 544007 108406 544063
rect 108462 544007 108530 544063
rect 108586 544007 108654 544063
rect 108710 544007 108778 544063
rect 108834 544007 108902 544063
rect 108958 544007 109026 544063
rect 109082 544007 109150 544063
rect 109206 544007 109274 544063
rect 109330 544007 109398 544063
rect 109454 544007 109522 544063
rect 109578 544007 109646 544063
rect 109702 544007 109770 544063
rect 109826 544007 109894 544063
rect 109950 544007 110018 544063
rect 110074 544007 110142 544063
rect 110198 544007 110266 544063
rect 110322 544007 110390 544063
rect 110446 544007 110514 544063
rect 110570 544007 110638 544063
rect 110694 544007 110762 544063
rect 110818 544007 110886 544063
rect 110942 544007 111010 544063
rect 111066 544007 111134 544063
rect 111190 544007 111258 544063
rect 111314 544007 111382 544063
rect 111438 544007 111506 544063
rect 111562 544007 111630 544063
rect 111686 544007 111754 544063
rect 111810 544007 111878 544063
rect 111934 544007 112002 544063
rect 112058 544007 112126 544063
rect 112182 544007 112250 544063
rect 112306 544007 112374 544063
rect 112430 544007 112498 544063
rect 112554 544007 112622 544063
rect 112678 544007 112746 544063
rect 112802 544007 112870 544063
rect 112926 544007 112994 544063
rect 113050 544007 113118 544063
rect 113174 544007 113242 544063
rect 113298 544007 113366 544063
rect 113422 544007 113490 544063
rect 113546 544007 113614 544063
rect 113670 544007 113738 544063
rect 113794 544007 113862 544063
rect 113918 544007 113986 544063
rect 114042 544007 114110 544063
rect 114166 544007 114234 544063
rect 114290 544007 114358 544063
rect 114414 544007 114482 544063
rect 114538 544007 114606 544063
rect 114662 544007 114730 544063
rect 114786 544007 114854 544063
rect 114910 544007 114978 544063
rect 115034 544007 115102 544063
rect 115158 544007 115226 544063
rect 115282 544007 115350 544063
rect 115406 544007 115474 544063
rect 115530 544007 115598 544063
rect 115654 544007 115722 544063
rect 115778 544007 115846 544063
rect 115902 544007 115970 544063
rect 116026 544007 116094 544063
rect 116150 544007 116218 544063
rect 116274 544007 116342 544063
rect 116398 544007 116466 544063
rect 116522 544007 116590 544063
rect 116646 544007 116714 544063
rect 116770 544007 116838 544063
rect 116894 544007 116962 544063
rect 117018 544007 117086 544063
rect 117142 544007 117210 544063
rect 117266 544007 117334 544063
rect 117390 544007 117458 544063
rect 117514 544007 117582 544063
rect 117638 544007 117706 544063
rect 117762 544007 117830 544063
rect 117886 544007 117954 544063
rect 118010 544007 118078 544063
rect 118134 544007 118202 544063
rect 118258 544007 118326 544063
rect 118382 544007 118450 544063
rect 118506 544007 118574 544063
rect 118630 544007 118698 544063
rect 118754 544007 118822 544063
rect 118878 544007 118946 544063
rect 119002 544007 119070 544063
rect 119126 544007 119194 544063
rect 119250 544007 119318 544063
rect 119374 544007 119442 544063
rect 119498 544007 119566 544063
rect 119622 544007 119690 544063
rect 119746 544007 119814 544063
rect 119870 544007 119938 544063
rect 119994 544007 120062 544063
rect 120118 544007 120186 544063
rect 120242 544007 120310 544063
rect 120366 544007 120434 544063
rect 120490 544007 120558 544063
rect 120614 544007 120682 544063
rect 120738 544007 120806 544063
rect 120862 544007 120930 544063
rect 120986 544007 121054 544063
rect 121110 544007 121178 544063
rect 121234 544007 121302 544063
rect 121358 544007 121426 544063
rect 121482 544007 121550 544063
rect 121606 544007 121674 544063
rect 121730 544007 121798 544063
rect 121854 544007 121920 544063
rect 104000 543939 121920 544007
rect 104000 543883 104066 543939
rect 104122 543883 104190 543939
rect 104246 543883 104314 543939
rect 104370 543883 104438 543939
rect 104494 543883 104562 543939
rect 104618 543883 104686 543939
rect 104742 543883 104810 543939
rect 104866 543883 104934 543939
rect 104990 543883 105058 543939
rect 105114 543883 105182 543939
rect 105238 543883 105306 543939
rect 105362 543883 105430 543939
rect 105486 543883 105554 543939
rect 105610 543883 105678 543939
rect 105734 543883 105802 543939
rect 105858 543883 105926 543939
rect 105982 543883 106050 543939
rect 106106 543883 106174 543939
rect 106230 543883 106298 543939
rect 106354 543883 106422 543939
rect 106478 543883 106546 543939
rect 106602 543883 106670 543939
rect 106726 543883 106794 543939
rect 106850 543883 106918 543939
rect 106974 543883 107042 543939
rect 107098 543883 107166 543939
rect 107222 543883 107290 543939
rect 107346 543883 107414 543939
rect 107470 543883 107538 543939
rect 107594 543883 107662 543939
rect 107718 543883 107786 543939
rect 107842 543883 107910 543939
rect 107966 543883 108034 543939
rect 108090 543883 108158 543939
rect 108214 543883 108282 543939
rect 108338 543883 108406 543939
rect 108462 543883 108530 543939
rect 108586 543883 108654 543939
rect 108710 543883 108778 543939
rect 108834 543883 108902 543939
rect 108958 543883 109026 543939
rect 109082 543883 109150 543939
rect 109206 543883 109274 543939
rect 109330 543883 109398 543939
rect 109454 543883 109522 543939
rect 109578 543883 109646 543939
rect 109702 543883 109770 543939
rect 109826 543883 109894 543939
rect 109950 543883 110018 543939
rect 110074 543883 110142 543939
rect 110198 543883 110266 543939
rect 110322 543883 110390 543939
rect 110446 543883 110514 543939
rect 110570 543883 110638 543939
rect 110694 543883 110762 543939
rect 110818 543883 110886 543939
rect 110942 543883 111010 543939
rect 111066 543883 111134 543939
rect 111190 543883 111258 543939
rect 111314 543883 111382 543939
rect 111438 543883 111506 543939
rect 111562 543883 111630 543939
rect 111686 543883 111754 543939
rect 111810 543883 111878 543939
rect 111934 543883 112002 543939
rect 112058 543883 112126 543939
rect 112182 543883 112250 543939
rect 112306 543883 112374 543939
rect 112430 543883 112498 543939
rect 112554 543883 112622 543939
rect 112678 543883 112746 543939
rect 112802 543883 112870 543939
rect 112926 543883 112994 543939
rect 113050 543883 113118 543939
rect 113174 543883 113242 543939
rect 113298 543883 113366 543939
rect 113422 543883 113490 543939
rect 113546 543883 113614 543939
rect 113670 543883 113738 543939
rect 113794 543883 113862 543939
rect 113918 543883 113986 543939
rect 114042 543883 114110 543939
rect 114166 543883 114234 543939
rect 114290 543883 114358 543939
rect 114414 543883 114482 543939
rect 114538 543883 114606 543939
rect 114662 543883 114730 543939
rect 114786 543883 114854 543939
rect 114910 543883 114978 543939
rect 115034 543883 115102 543939
rect 115158 543883 115226 543939
rect 115282 543883 115350 543939
rect 115406 543883 115474 543939
rect 115530 543883 115598 543939
rect 115654 543883 115722 543939
rect 115778 543883 115846 543939
rect 115902 543883 115970 543939
rect 116026 543883 116094 543939
rect 116150 543883 116218 543939
rect 116274 543883 116342 543939
rect 116398 543883 116466 543939
rect 116522 543883 116590 543939
rect 116646 543883 116714 543939
rect 116770 543883 116838 543939
rect 116894 543883 116962 543939
rect 117018 543883 117086 543939
rect 117142 543883 117210 543939
rect 117266 543883 117334 543939
rect 117390 543883 117458 543939
rect 117514 543883 117582 543939
rect 117638 543883 117706 543939
rect 117762 543883 117830 543939
rect 117886 543883 117954 543939
rect 118010 543883 118078 543939
rect 118134 543883 118202 543939
rect 118258 543883 118326 543939
rect 118382 543883 118450 543939
rect 118506 543883 118574 543939
rect 118630 543883 118698 543939
rect 118754 543883 118822 543939
rect 118878 543883 118946 543939
rect 119002 543883 119070 543939
rect 119126 543883 119194 543939
rect 119250 543883 119318 543939
rect 119374 543883 119442 543939
rect 119498 543883 119566 543939
rect 119622 543883 119690 543939
rect 119746 543883 119814 543939
rect 119870 543883 119938 543939
rect 119994 543883 120062 543939
rect 120118 543883 120186 543939
rect 120242 543883 120310 543939
rect 120366 543883 120434 543939
rect 120490 543883 120558 543939
rect 120614 543883 120682 543939
rect 120738 543883 120806 543939
rect 120862 543883 120930 543939
rect 120986 543883 121054 543939
rect 121110 543883 121178 543939
rect 121234 543883 121302 543939
rect 121358 543883 121426 543939
rect 121482 543883 121550 543939
rect 121606 543883 121674 543939
rect 121730 543883 121798 543939
rect 121854 543883 121920 543939
rect 104000 543826 121920 543883
rect 128298 544102 128918 544170
rect 128298 544046 128394 544102
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 128918 544102
rect 128298 543978 128918 544046
rect 128298 543922 128394 543978
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 128918 543978
rect 128298 539352 128918 543922
rect 132018 598172 132638 598268
rect 132018 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 132638 598172
rect 132018 598048 132638 598116
rect 132018 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 132638 598048
rect 132018 597924 132638 597992
rect 132018 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 132638 597924
rect 132018 597800 132638 597868
rect 132018 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 132638 597800
rect 132018 586350 132638 597744
rect 132018 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 132638 586350
rect 132018 586226 132638 586294
rect 132018 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 132638 586226
rect 132018 586102 132638 586170
rect 132018 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 132638 586102
rect 132018 585978 132638 586046
rect 132018 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 132638 585978
rect 132018 568350 132638 585922
rect 132018 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 132638 568350
rect 132018 568226 132638 568294
rect 132018 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 132638 568226
rect 132018 568102 132638 568170
rect 132018 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 132638 568102
rect 132018 567978 132638 568046
rect 132018 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 132638 567978
rect 132018 550350 132638 567922
rect 132018 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 132638 550350
rect 132018 550226 132638 550294
rect 132018 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 132638 550226
rect 132018 550102 132638 550170
rect 132018 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 132638 550102
rect 132018 549978 132638 550046
rect 132018 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 132638 549978
rect 132018 542072 132638 549922
rect 159018 597212 159638 598268
rect 159018 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 159638 597212
rect 159018 597088 159638 597156
rect 159018 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 159638 597088
rect 159018 596964 159638 597032
rect 159018 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 159638 596964
rect 159018 596840 159638 596908
rect 159018 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 159638 596840
rect 159018 580350 159638 596784
rect 159018 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 159638 580350
rect 159018 580226 159638 580294
rect 159018 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 159638 580226
rect 159018 580102 159638 580170
rect 159018 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 159638 580102
rect 159018 579978 159638 580046
rect 159018 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 159638 579978
rect 159018 562350 159638 579922
rect 159018 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 159638 562350
rect 159018 562226 159638 562294
rect 159018 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 159638 562226
rect 159018 562102 159638 562170
rect 159018 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 159638 562102
rect 159018 561978 159638 562046
rect 159018 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 159638 561978
rect 159018 544350 159638 561922
rect 159018 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 159638 544350
rect 159018 544226 159638 544294
rect 159018 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 159638 544226
rect 159018 544102 159638 544170
rect 159018 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 159638 544102
rect 159018 543978 159638 544046
rect 159018 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 159638 543978
rect 71840 532388 82880 532440
rect 71840 532332 71876 532388
rect 71932 532332 72000 532388
rect 72056 532332 72124 532388
rect 72180 532332 72248 532388
rect 72304 532332 72372 532388
rect 72428 532332 72496 532388
rect 72552 532332 72620 532388
rect 72676 532332 72744 532388
rect 72800 532332 72868 532388
rect 72924 532332 72992 532388
rect 73048 532332 73116 532388
rect 73172 532332 73240 532388
rect 73296 532332 73364 532388
rect 73420 532332 73488 532388
rect 73544 532332 73612 532388
rect 73668 532332 73736 532388
rect 73792 532332 73860 532388
rect 73916 532332 73984 532388
rect 74040 532332 74108 532388
rect 74164 532332 74232 532388
rect 74288 532332 74356 532388
rect 74412 532332 74480 532388
rect 74536 532332 74604 532388
rect 74660 532332 74728 532388
rect 74784 532332 74852 532388
rect 74908 532332 74976 532388
rect 75032 532332 75100 532388
rect 75156 532332 75224 532388
rect 75280 532332 75348 532388
rect 75404 532332 75472 532388
rect 75528 532332 75596 532388
rect 75652 532332 75720 532388
rect 75776 532332 75844 532388
rect 75900 532332 75968 532388
rect 76024 532332 76092 532388
rect 76148 532332 76216 532388
rect 76272 532332 76340 532388
rect 76396 532332 76464 532388
rect 76520 532332 76588 532388
rect 76644 532332 76712 532388
rect 76768 532332 76836 532388
rect 76892 532332 76960 532388
rect 77016 532332 77084 532388
rect 77140 532332 77208 532388
rect 77264 532332 77332 532388
rect 77388 532332 77456 532388
rect 77512 532332 77580 532388
rect 77636 532332 77704 532388
rect 77760 532332 77828 532388
rect 77884 532332 77952 532388
rect 78008 532332 78076 532388
rect 78132 532332 78200 532388
rect 78256 532332 78324 532388
rect 78380 532332 78448 532388
rect 78504 532332 78572 532388
rect 78628 532332 78696 532388
rect 78752 532332 78820 532388
rect 78876 532332 78944 532388
rect 79000 532332 79068 532388
rect 79124 532332 79192 532388
rect 79248 532332 79316 532388
rect 79372 532332 79440 532388
rect 79496 532332 79564 532388
rect 79620 532332 79688 532388
rect 79744 532332 79812 532388
rect 79868 532332 79936 532388
rect 79992 532332 80060 532388
rect 80116 532332 80184 532388
rect 80240 532332 80308 532388
rect 80364 532332 80432 532388
rect 80488 532332 80556 532388
rect 80612 532332 80680 532388
rect 80736 532332 80804 532388
rect 80860 532332 80928 532388
rect 80984 532332 81052 532388
rect 81108 532332 81176 532388
rect 81232 532332 81300 532388
rect 81356 532332 81424 532388
rect 81480 532332 81548 532388
rect 81604 532332 81672 532388
rect 81728 532332 81796 532388
rect 81852 532332 81920 532388
rect 81976 532332 82044 532388
rect 82100 532332 82168 532388
rect 82224 532332 82292 532388
rect 82348 532332 82416 532388
rect 82472 532332 82540 532388
rect 82596 532332 82664 532388
rect 82720 532332 82788 532388
rect 82844 532332 82880 532388
rect 71840 532280 82880 532332
rect 159018 526350 159638 543922
rect 159018 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 159638 526350
rect 159018 526226 159638 526294
rect 94240 526148 114400 526200
rect 94240 526092 94310 526148
rect 94366 526092 94434 526148
rect 94490 526092 94558 526148
rect 94614 526092 94682 526148
rect 94738 526092 94806 526148
rect 94862 526092 94930 526148
rect 94986 526092 95054 526148
rect 95110 526092 95178 526148
rect 95234 526092 95302 526148
rect 95358 526092 95426 526148
rect 95482 526092 95550 526148
rect 95606 526092 95674 526148
rect 95730 526092 95798 526148
rect 95854 526092 95922 526148
rect 95978 526092 96046 526148
rect 96102 526092 96170 526148
rect 96226 526092 96294 526148
rect 96350 526092 96418 526148
rect 96474 526092 96542 526148
rect 96598 526092 96666 526148
rect 96722 526092 96790 526148
rect 96846 526092 96914 526148
rect 96970 526092 97038 526148
rect 97094 526092 97162 526148
rect 97218 526092 97286 526148
rect 97342 526092 97410 526148
rect 97466 526092 97534 526148
rect 97590 526092 97658 526148
rect 97714 526092 97782 526148
rect 97838 526092 97906 526148
rect 97962 526092 98030 526148
rect 98086 526092 98154 526148
rect 98210 526092 98278 526148
rect 98334 526092 98402 526148
rect 98458 526092 98526 526148
rect 98582 526092 98650 526148
rect 98706 526092 98774 526148
rect 98830 526092 98898 526148
rect 98954 526092 99022 526148
rect 99078 526092 99146 526148
rect 99202 526092 99270 526148
rect 99326 526092 99394 526148
rect 99450 526092 99518 526148
rect 99574 526092 99642 526148
rect 99698 526092 99766 526148
rect 99822 526092 99890 526148
rect 99946 526092 100014 526148
rect 100070 526092 100138 526148
rect 100194 526092 100262 526148
rect 100318 526092 100386 526148
rect 100442 526092 100510 526148
rect 100566 526092 100634 526148
rect 100690 526092 100758 526148
rect 100814 526092 100882 526148
rect 100938 526092 101006 526148
rect 101062 526092 101130 526148
rect 101186 526092 101254 526148
rect 101310 526092 101378 526148
rect 101434 526092 101502 526148
rect 101558 526092 101626 526148
rect 101682 526092 101750 526148
rect 101806 526092 101874 526148
rect 101930 526092 101998 526148
rect 102054 526092 102122 526148
rect 102178 526092 102246 526148
rect 102302 526092 102370 526148
rect 102426 526092 102494 526148
rect 102550 526092 102618 526148
rect 102674 526092 102742 526148
rect 102798 526092 102866 526148
rect 102922 526092 102990 526148
rect 103046 526092 103114 526148
rect 103170 526092 103238 526148
rect 103294 526092 103362 526148
rect 103418 526092 103486 526148
rect 103542 526092 103610 526148
rect 103666 526092 103734 526148
rect 103790 526092 103858 526148
rect 103914 526092 103982 526148
rect 104038 526092 104106 526148
rect 104162 526092 104230 526148
rect 104286 526092 104354 526148
rect 104410 526092 104478 526148
rect 104534 526092 104602 526148
rect 104658 526092 104726 526148
rect 104782 526092 104850 526148
rect 104906 526092 104974 526148
rect 105030 526092 105098 526148
rect 105154 526092 105222 526148
rect 105278 526092 105346 526148
rect 105402 526092 105470 526148
rect 105526 526092 105594 526148
rect 105650 526092 105718 526148
rect 105774 526092 105842 526148
rect 105898 526092 105966 526148
rect 106022 526092 106090 526148
rect 106146 526092 106214 526148
rect 106270 526092 106338 526148
rect 106394 526092 106462 526148
rect 106518 526092 106586 526148
rect 106642 526092 106710 526148
rect 106766 526092 106834 526148
rect 106890 526092 106958 526148
rect 107014 526092 107082 526148
rect 107138 526092 107206 526148
rect 107262 526092 107330 526148
rect 107386 526092 107454 526148
rect 107510 526092 107578 526148
rect 107634 526092 107702 526148
rect 107758 526092 107826 526148
rect 107882 526092 107950 526148
rect 108006 526092 108074 526148
rect 108130 526092 108198 526148
rect 108254 526092 108322 526148
rect 108378 526092 108446 526148
rect 108502 526092 108570 526148
rect 108626 526092 108694 526148
rect 108750 526092 108818 526148
rect 108874 526092 108942 526148
rect 108998 526092 109066 526148
rect 109122 526092 109190 526148
rect 109246 526092 109314 526148
rect 109370 526092 109438 526148
rect 109494 526092 109562 526148
rect 109618 526092 109686 526148
rect 109742 526092 109810 526148
rect 109866 526092 109934 526148
rect 109990 526092 110058 526148
rect 110114 526092 110182 526148
rect 110238 526092 110306 526148
rect 110362 526092 110430 526148
rect 110486 526092 110554 526148
rect 110610 526092 110678 526148
rect 110734 526092 110802 526148
rect 110858 526092 110926 526148
rect 110982 526092 111050 526148
rect 111106 526092 111174 526148
rect 111230 526092 111298 526148
rect 111354 526092 111422 526148
rect 111478 526092 111546 526148
rect 111602 526092 111670 526148
rect 111726 526092 111794 526148
rect 111850 526092 111918 526148
rect 111974 526092 112042 526148
rect 112098 526092 112166 526148
rect 112222 526092 112290 526148
rect 112346 526092 112414 526148
rect 112470 526092 112538 526148
rect 112594 526092 112662 526148
rect 112718 526092 112786 526148
rect 112842 526092 112910 526148
rect 112966 526092 113034 526148
rect 113090 526092 113158 526148
rect 113214 526092 113282 526148
rect 113338 526092 113406 526148
rect 113462 526092 113530 526148
rect 113586 526092 113654 526148
rect 113710 526092 113778 526148
rect 113834 526092 113902 526148
rect 113958 526092 114026 526148
rect 114082 526092 114150 526148
rect 114206 526092 114274 526148
rect 114330 526092 114400 526148
rect 94240 526040 114400 526092
rect 159018 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 159638 526226
rect 159018 526102 159638 526170
rect 159018 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 159638 526102
rect 39858 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 40478 514350
rect 39858 514226 40478 514294
rect 39858 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 40478 514226
rect 159018 525978 159638 526046
rect 159018 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 159638 525978
rect 39858 514102 40478 514170
rect 39858 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514046 40478 514102
rect 39858 513978 40478 514046
rect 39858 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513922 40478 513978
rect 39858 496350 40478 513922
rect 60800 514130 66400 514200
rect 60800 514074 60844 514130
rect 60900 514074 60968 514130
rect 61024 514074 61092 514130
rect 61148 514074 61216 514130
rect 61272 514074 61340 514130
rect 61396 514074 61464 514130
rect 61520 514074 61588 514130
rect 61644 514074 61712 514130
rect 61768 514074 61836 514130
rect 61892 514074 61960 514130
rect 62016 514074 62084 514130
rect 62140 514074 62208 514130
rect 62264 514074 62332 514130
rect 62388 514074 62456 514130
rect 62512 514074 62580 514130
rect 62636 514074 62704 514130
rect 62760 514074 62828 514130
rect 62884 514074 62952 514130
rect 63008 514074 63076 514130
rect 63132 514074 63200 514130
rect 63256 514074 63324 514130
rect 63380 514074 63448 514130
rect 63504 514074 63572 514130
rect 63628 514074 63696 514130
rect 63752 514074 63820 514130
rect 63876 514074 63944 514130
rect 64000 514074 64068 514130
rect 64124 514074 64192 514130
rect 64248 514074 64316 514130
rect 64372 514074 64440 514130
rect 64496 514074 64564 514130
rect 64620 514074 64688 514130
rect 64744 514074 64812 514130
rect 64868 514074 64936 514130
rect 64992 514074 65060 514130
rect 65116 514074 65184 514130
rect 65240 514074 65308 514130
rect 65364 514074 65432 514130
rect 65488 514074 65556 514130
rect 65612 514074 65680 514130
rect 65736 514074 65804 514130
rect 65860 514074 65928 514130
rect 65984 514074 66052 514130
rect 66108 514074 66176 514130
rect 66232 514074 66300 514130
rect 66356 514074 66400 514130
rect 60800 514006 66400 514074
rect 60800 513950 60844 514006
rect 60900 513950 60968 514006
rect 61024 513950 61092 514006
rect 61148 513950 61216 514006
rect 61272 513950 61340 514006
rect 61396 513950 61464 514006
rect 61520 513950 61588 514006
rect 61644 513950 61712 514006
rect 61768 513950 61836 514006
rect 61892 513950 61960 514006
rect 62016 513950 62084 514006
rect 62140 513950 62208 514006
rect 62264 513950 62332 514006
rect 62388 513950 62456 514006
rect 62512 513950 62580 514006
rect 62636 513950 62704 514006
rect 62760 513950 62828 514006
rect 62884 513950 62952 514006
rect 63008 513950 63076 514006
rect 63132 513950 63200 514006
rect 63256 513950 63324 514006
rect 63380 513950 63448 514006
rect 63504 513950 63572 514006
rect 63628 513950 63696 514006
rect 63752 513950 63820 514006
rect 63876 513950 63944 514006
rect 64000 513950 64068 514006
rect 64124 513950 64192 514006
rect 64248 513950 64316 514006
rect 64372 513950 64440 514006
rect 64496 513950 64564 514006
rect 64620 513950 64688 514006
rect 64744 513950 64812 514006
rect 64868 513950 64936 514006
rect 64992 513950 65060 514006
rect 65116 513950 65184 514006
rect 65240 513950 65308 514006
rect 65364 513950 65432 514006
rect 65488 513950 65556 514006
rect 65612 513950 65680 514006
rect 65736 513950 65804 514006
rect 65860 513950 65928 514006
rect 65984 513950 66052 514006
rect 66108 513950 66176 514006
rect 66232 513950 66300 514006
rect 66356 513950 66400 514006
rect 60800 513880 66400 513950
rect 87840 508388 98400 508440
rect 87840 508332 87884 508388
rect 87940 508332 88008 508388
rect 88064 508332 88132 508388
rect 88188 508332 88256 508388
rect 88312 508332 88380 508388
rect 88436 508332 88504 508388
rect 88560 508332 88628 508388
rect 88684 508332 88752 508388
rect 88808 508332 88876 508388
rect 88932 508332 89000 508388
rect 89056 508332 89124 508388
rect 89180 508332 89248 508388
rect 89304 508332 89372 508388
rect 89428 508332 89496 508388
rect 89552 508332 89620 508388
rect 89676 508332 89744 508388
rect 89800 508332 89868 508388
rect 89924 508332 89992 508388
rect 90048 508332 90116 508388
rect 90172 508332 90240 508388
rect 90296 508332 90364 508388
rect 90420 508332 90488 508388
rect 90544 508332 90612 508388
rect 90668 508332 90736 508388
rect 90792 508332 90860 508388
rect 90916 508332 90984 508388
rect 91040 508332 91108 508388
rect 91164 508332 91232 508388
rect 91288 508332 91356 508388
rect 91412 508332 91480 508388
rect 91536 508332 91604 508388
rect 91660 508332 91728 508388
rect 91784 508332 91852 508388
rect 91908 508332 91976 508388
rect 92032 508332 92100 508388
rect 92156 508332 92224 508388
rect 92280 508332 92348 508388
rect 92404 508332 92472 508388
rect 92528 508332 92596 508388
rect 92652 508332 92720 508388
rect 92776 508332 92844 508388
rect 92900 508332 92968 508388
rect 93024 508332 93092 508388
rect 93148 508332 93216 508388
rect 93272 508332 93340 508388
rect 93396 508332 93464 508388
rect 93520 508332 93588 508388
rect 93644 508332 93712 508388
rect 93768 508332 93836 508388
rect 93892 508332 93960 508388
rect 94016 508332 94084 508388
rect 94140 508332 94208 508388
rect 94264 508332 94332 508388
rect 94388 508332 94456 508388
rect 94512 508332 94580 508388
rect 94636 508332 94704 508388
rect 94760 508332 94828 508388
rect 94884 508332 94952 508388
rect 95008 508332 95076 508388
rect 95132 508332 95200 508388
rect 95256 508332 95324 508388
rect 95380 508332 95448 508388
rect 95504 508332 95572 508388
rect 95628 508332 95696 508388
rect 95752 508332 95820 508388
rect 95876 508332 95944 508388
rect 96000 508332 96068 508388
rect 96124 508332 96192 508388
rect 96248 508332 96316 508388
rect 96372 508332 96440 508388
rect 96496 508332 96564 508388
rect 96620 508332 96688 508388
rect 96744 508332 96812 508388
rect 96868 508332 96936 508388
rect 96992 508332 97060 508388
rect 97116 508332 97184 508388
rect 97240 508332 97308 508388
rect 97364 508332 97432 508388
rect 97488 508332 97556 508388
rect 97612 508332 97680 508388
rect 97736 508332 97804 508388
rect 97860 508332 97928 508388
rect 97984 508332 98052 508388
rect 98108 508332 98176 508388
rect 98232 508332 98300 508388
rect 98356 508332 98400 508388
rect 87840 508280 98400 508332
rect 159018 508350 159638 525922
rect 159018 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 159638 508350
rect 159018 508226 159638 508294
rect 159018 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 159638 508226
rect 87680 508068 98240 508120
rect 87680 508012 87724 508068
rect 87780 508012 87848 508068
rect 87904 508012 87972 508068
rect 88028 508012 88096 508068
rect 88152 508012 88220 508068
rect 88276 508012 88344 508068
rect 88400 508012 88468 508068
rect 88524 508012 88592 508068
rect 88648 508012 88716 508068
rect 88772 508012 88840 508068
rect 88896 508012 88964 508068
rect 89020 508012 89088 508068
rect 89144 508012 89212 508068
rect 89268 508012 89336 508068
rect 89392 508012 89460 508068
rect 89516 508012 89584 508068
rect 89640 508012 89708 508068
rect 89764 508012 89832 508068
rect 89888 508012 89956 508068
rect 90012 508012 90080 508068
rect 90136 508012 90204 508068
rect 90260 508012 90328 508068
rect 90384 508012 90452 508068
rect 90508 508012 90576 508068
rect 90632 508012 90700 508068
rect 90756 508012 90824 508068
rect 90880 508012 90948 508068
rect 91004 508012 91072 508068
rect 91128 508012 91196 508068
rect 91252 508012 91320 508068
rect 91376 508012 91444 508068
rect 91500 508012 91568 508068
rect 91624 508012 91692 508068
rect 91748 508012 91816 508068
rect 91872 508012 91940 508068
rect 91996 508012 92064 508068
rect 92120 508012 92188 508068
rect 92244 508012 92312 508068
rect 92368 508012 92436 508068
rect 92492 508012 92560 508068
rect 92616 508012 92684 508068
rect 92740 508012 92808 508068
rect 92864 508012 92932 508068
rect 92988 508012 93056 508068
rect 93112 508012 93180 508068
rect 93236 508012 93304 508068
rect 93360 508012 93428 508068
rect 93484 508012 93552 508068
rect 93608 508012 93676 508068
rect 93732 508012 93800 508068
rect 93856 508012 93924 508068
rect 93980 508012 94048 508068
rect 94104 508012 94172 508068
rect 94228 508012 94296 508068
rect 94352 508012 94420 508068
rect 94476 508012 94544 508068
rect 94600 508012 94668 508068
rect 94724 508012 94792 508068
rect 94848 508012 94916 508068
rect 94972 508012 95040 508068
rect 95096 508012 95164 508068
rect 95220 508012 95288 508068
rect 95344 508012 95412 508068
rect 95468 508012 95536 508068
rect 95592 508012 95660 508068
rect 95716 508012 95784 508068
rect 95840 508012 95908 508068
rect 95964 508012 96032 508068
rect 96088 508012 96156 508068
rect 96212 508012 96280 508068
rect 96336 508012 96404 508068
rect 96460 508012 96528 508068
rect 96584 508012 96652 508068
rect 96708 508012 96776 508068
rect 96832 508012 96900 508068
rect 96956 508012 97024 508068
rect 97080 508012 97148 508068
rect 97204 508012 97272 508068
rect 97328 508012 97396 508068
rect 97452 508012 97520 508068
rect 97576 508012 97644 508068
rect 97700 508012 97768 508068
rect 97824 508012 97892 508068
rect 97948 508012 98016 508068
rect 98072 508012 98140 508068
rect 98196 508012 98240 508068
rect 87680 507960 98240 508012
rect 159018 508102 159638 508170
rect 159018 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 159638 508102
rect 159018 507978 159638 508046
rect 159018 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 159638 507978
rect 39858 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496294 40478 496350
rect 39858 496226 40478 496294
rect 61920 496388 68000 496440
rect 61920 496332 61956 496388
rect 62012 496332 62080 496388
rect 62136 496332 62204 496388
rect 62260 496332 62328 496388
rect 62384 496332 62452 496388
rect 62508 496332 62576 496388
rect 62632 496332 62700 496388
rect 62756 496332 62824 496388
rect 62880 496332 62948 496388
rect 63004 496332 63072 496388
rect 63128 496332 63196 496388
rect 63252 496332 63320 496388
rect 63376 496332 63444 496388
rect 63500 496332 63568 496388
rect 63624 496332 63692 496388
rect 63748 496332 63816 496388
rect 63872 496332 63940 496388
rect 63996 496332 64064 496388
rect 64120 496332 64188 496388
rect 64244 496332 64312 496388
rect 64368 496332 64436 496388
rect 64492 496332 64560 496388
rect 64616 496332 64684 496388
rect 64740 496332 64808 496388
rect 64864 496332 64932 496388
rect 64988 496332 65056 496388
rect 65112 496332 65180 496388
rect 65236 496332 65304 496388
rect 65360 496332 65428 496388
rect 65484 496332 65552 496388
rect 65608 496332 65676 496388
rect 65732 496332 65800 496388
rect 65856 496332 65924 496388
rect 65980 496332 66048 496388
rect 66104 496332 66172 496388
rect 66228 496332 66296 496388
rect 66352 496332 66420 496388
rect 66476 496332 66544 496388
rect 66600 496332 66668 496388
rect 66724 496332 66792 496388
rect 66848 496332 66916 496388
rect 66972 496332 67040 496388
rect 67096 496332 67164 496388
rect 67220 496332 67288 496388
rect 67344 496332 67412 496388
rect 67468 496332 67536 496388
rect 67592 496332 67660 496388
rect 67716 496332 67784 496388
rect 67840 496332 67908 496388
rect 67964 496332 68000 496388
rect 61920 496280 68000 496332
rect 39858 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 40478 496226
rect 39858 496102 40478 496170
rect 39858 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496046 40478 496102
rect 39858 495978 40478 496046
rect 39858 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495922 40478 495978
rect 39858 478350 40478 495922
rect 62080 496063 68160 496120
rect 62080 496007 62116 496063
rect 62172 496007 62240 496063
rect 62296 496007 62364 496063
rect 62420 496007 62488 496063
rect 62544 496007 62612 496063
rect 62668 496007 62736 496063
rect 62792 496007 62860 496063
rect 62916 496007 62984 496063
rect 63040 496007 63108 496063
rect 63164 496007 63232 496063
rect 63288 496007 63356 496063
rect 63412 496007 63480 496063
rect 63536 496007 63604 496063
rect 63660 496007 63728 496063
rect 63784 496007 63852 496063
rect 63908 496007 63976 496063
rect 64032 496007 64100 496063
rect 64156 496007 64224 496063
rect 64280 496007 64348 496063
rect 64404 496007 64472 496063
rect 64528 496007 64596 496063
rect 64652 496007 64720 496063
rect 64776 496007 64844 496063
rect 64900 496007 64968 496063
rect 65024 496007 65092 496063
rect 65148 496007 65216 496063
rect 65272 496007 65340 496063
rect 65396 496007 65464 496063
rect 65520 496007 65588 496063
rect 65644 496007 65712 496063
rect 65768 496007 65836 496063
rect 65892 496007 65960 496063
rect 66016 496007 66084 496063
rect 66140 496007 66208 496063
rect 66264 496007 66332 496063
rect 66388 496007 66456 496063
rect 66512 496007 66580 496063
rect 66636 496007 66704 496063
rect 66760 496007 66828 496063
rect 66884 496007 66952 496063
rect 67008 496007 67076 496063
rect 67132 496007 67200 496063
rect 67256 496007 67324 496063
rect 67380 496007 67448 496063
rect 67504 496007 67572 496063
rect 67628 496007 67696 496063
rect 67752 496007 67820 496063
rect 67876 496007 67944 496063
rect 68000 496007 68068 496063
rect 68124 496007 68160 496063
rect 62080 495939 68160 496007
rect 62080 495883 62116 495939
rect 62172 495883 62240 495939
rect 62296 495883 62364 495939
rect 62420 495883 62488 495939
rect 62544 495883 62612 495939
rect 62668 495883 62736 495939
rect 62792 495883 62860 495939
rect 62916 495883 62984 495939
rect 63040 495883 63108 495939
rect 63164 495883 63232 495939
rect 63288 495883 63356 495939
rect 63412 495883 63480 495939
rect 63536 495883 63604 495939
rect 63660 495883 63728 495939
rect 63784 495883 63852 495939
rect 63908 495883 63976 495939
rect 64032 495883 64100 495939
rect 64156 495883 64224 495939
rect 64280 495883 64348 495939
rect 64404 495883 64472 495939
rect 64528 495883 64596 495939
rect 64652 495883 64720 495939
rect 64776 495883 64844 495939
rect 64900 495883 64968 495939
rect 65024 495883 65092 495939
rect 65148 495883 65216 495939
rect 65272 495883 65340 495939
rect 65396 495883 65464 495939
rect 65520 495883 65588 495939
rect 65644 495883 65712 495939
rect 65768 495883 65836 495939
rect 65892 495883 65960 495939
rect 66016 495883 66084 495939
rect 66140 495883 66208 495939
rect 66264 495883 66332 495939
rect 66388 495883 66456 495939
rect 66512 495883 66580 495939
rect 66636 495883 66704 495939
rect 66760 495883 66828 495939
rect 66884 495883 66952 495939
rect 67008 495883 67076 495939
rect 67132 495883 67200 495939
rect 67256 495883 67324 495939
rect 67380 495883 67448 495939
rect 67504 495883 67572 495939
rect 67628 495883 67696 495939
rect 67752 495883 67820 495939
rect 67876 495883 67944 495939
rect 68000 495883 68068 495939
rect 68124 495883 68160 495939
rect 62080 495826 68160 495883
rect 82880 490413 83088 490446
rect 82880 490357 82894 490413
rect 82950 490357 83018 490413
rect 83074 490357 83088 490413
rect 82880 490289 83088 490357
rect 82880 490233 82894 490289
rect 82950 490233 83018 490289
rect 83074 490233 83088 490289
rect 82880 490200 83088 490233
rect 83128 490413 83584 490446
rect 83128 490357 83142 490413
rect 83198 490357 83266 490413
rect 83322 490357 83390 490413
rect 83446 490357 83514 490413
rect 83570 490357 83584 490413
rect 83128 490289 83584 490357
rect 83128 490233 83142 490289
rect 83198 490233 83266 490289
rect 83322 490233 83390 490289
rect 83446 490233 83514 490289
rect 83570 490233 83584 490289
rect 83128 490200 83584 490233
rect 83624 490413 84080 490446
rect 83624 490357 83638 490413
rect 83694 490357 83762 490413
rect 83818 490357 83886 490413
rect 83942 490357 84010 490413
rect 84066 490357 84080 490413
rect 83624 490289 84080 490357
rect 83624 490233 83638 490289
rect 83694 490233 83762 490289
rect 83818 490233 83886 490289
rect 83942 490233 84010 490289
rect 84066 490233 84080 490289
rect 83624 490200 84080 490233
rect 84120 490413 84576 490446
rect 84120 490357 84134 490413
rect 84190 490357 84258 490413
rect 84314 490357 84382 490413
rect 84438 490357 84506 490413
rect 84562 490357 84576 490413
rect 84120 490289 84576 490357
rect 84120 490233 84134 490289
rect 84190 490233 84258 490289
rect 84314 490233 84382 490289
rect 84438 490233 84506 490289
rect 84562 490233 84576 490289
rect 84120 490200 84576 490233
rect 84616 490413 85072 490446
rect 84616 490357 84630 490413
rect 84686 490357 84754 490413
rect 84810 490357 84878 490413
rect 84934 490357 85002 490413
rect 85058 490357 85072 490413
rect 84616 490289 85072 490357
rect 84616 490233 84630 490289
rect 84686 490233 84754 490289
rect 84810 490233 84878 490289
rect 84934 490233 85002 490289
rect 85058 490233 85072 490289
rect 84616 490200 85072 490233
rect 85112 490413 85568 490446
rect 85112 490357 85126 490413
rect 85182 490357 85250 490413
rect 85306 490357 85374 490413
rect 85430 490357 85498 490413
rect 85554 490357 85568 490413
rect 85112 490289 85568 490357
rect 85112 490233 85126 490289
rect 85182 490233 85250 490289
rect 85306 490233 85374 490289
rect 85430 490233 85498 490289
rect 85554 490233 85568 490289
rect 85112 490200 85568 490233
rect 85608 490413 86064 490446
rect 85608 490357 85622 490413
rect 85678 490357 85746 490413
rect 85802 490357 85870 490413
rect 85926 490357 85994 490413
rect 86050 490357 86064 490413
rect 85608 490289 86064 490357
rect 85608 490233 85622 490289
rect 85678 490233 85746 490289
rect 85802 490233 85870 490289
rect 85926 490233 85994 490289
rect 86050 490233 86064 490289
rect 85608 490200 86064 490233
rect 86104 490413 86560 490446
rect 86104 490357 86118 490413
rect 86174 490357 86242 490413
rect 86298 490357 86366 490413
rect 86422 490357 86490 490413
rect 86546 490357 86560 490413
rect 86104 490289 86560 490357
rect 86104 490233 86118 490289
rect 86174 490233 86242 490289
rect 86298 490233 86366 490289
rect 86422 490233 86490 490289
rect 86546 490233 86560 490289
rect 86104 490200 86560 490233
rect 128298 490350 128918 491128
rect 128298 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 128918 490350
rect 128298 490226 128918 490294
rect 128298 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 128918 490226
rect 128298 490102 128918 490170
rect 128298 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 128918 490102
rect 82720 489988 82928 490040
rect 82720 489932 82734 489988
rect 82790 489932 82858 489988
rect 82914 489932 82928 489988
rect 82720 489880 82928 489932
rect 82968 489988 83424 490040
rect 82968 489932 82982 489988
rect 83038 489932 83106 489988
rect 83162 489932 83230 489988
rect 83286 489932 83354 489988
rect 83410 489932 83424 489988
rect 82968 489880 83424 489932
rect 83464 489988 83920 490040
rect 83464 489932 83478 489988
rect 83534 489932 83602 489988
rect 83658 489932 83726 489988
rect 83782 489932 83850 489988
rect 83906 489932 83920 489988
rect 83464 489880 83920 489932
rect 83960 489988 84416 490040
rect 83960 489932 83974 489988
rect 84030 489932 84098 489988
rect 84154 489932 84222 489988
rect 84278 489932 84346 489988
rect 84402 489932 84416 489988
rect 83960 489880 84416 489932
rect 84456 489988 84912 490040
rect 84456 489932 84470 489988
rect 84526 489932 84594 489988
rect 84650 489932 84718 489988
rect 84774 489932 84842 489988
rect 84898 489932 84912 489988
rect 84456 489880 84912 489932
rect 84952 489988 85408 490040
rect 84952 489932 84966 489988
rect 85022 489932 85090 489988
rect 85146 489932 85214 489988
rect 85270 489932 85338 489988
rect 85394 489932 85408 489988
rect 84952 489880 85408 489932
rect 85448 489988 85904 490040
rect 85448 489932 85462 489988
rect 85518 489932 85586 489988
rect 85642 489932 85710 489988
rect 85766 489932 85834 489988
rect 85890 489932 85904 489988
rect 85448 489880 85904 489932
rect 85944 489988 86400 490040
rect 85944 489932 85958 489988
rect 86014 489932 86082 489988
rect 86138 489932 86206 489988
rect 86262 489932 86330 489988
rect 86386 489932 86400 489988
rect 85944 489880 86400 489932
rect 128298 489978 128918 490046
rect 128298 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 128918 489978
rect 39858 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 40478 478350
rect 39858 478226 40478 478294
rect 39858 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 40478 478226
rect 39858 478102 40478 478170
rect 39858 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 40478 478102
rect 39858 477978 40478 478046
rect 39858 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 40478 477978
rect 39858 460350 40478 477922
rect 39858 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 40478 460350
rect 39858 460226 40478 460294
rect 39858 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 40478 460226
rect 39858 460102 40478 460170
rect 39858 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 40478 460102
rect 39858 459978 40478 460046
rect 39858 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 40478 459978
rect 39858 442350 40478 459922
rect 39858 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 40478 442350
rect 39858 442226 40478 442294
rect 39858 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 40478 442226
rect 39858 442102 40478 442170
rect 39858 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 40478 442102
rect 39858 441978 40478 442046
rect 39858 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 40478 441978
rect 39858 424350 40478 441922
rect 39858 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 40478 424350
rect 39858 424226 40478 424294
rect 39858 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 40478 424226
rect 39858 424102 40478 424170
rect 39858 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 40478 424102
rect 39858 423978 40478 424046
rect 39858 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 40478 423978
rect 39858 406350 40478 423922
rect 39858 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 40478 406350
rect 39858 406226 40478 406294
rect 39858 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 40478 406226
rect 39858 406102 40478 406170
rect 39858 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 40478 406102
rect 39858 405978 40478 406046
rect 39858 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 40478 405978
rect 39858 388350 40478 405922
rect 39858 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 40478 388350
rect 39858 388226 40478 388294
rect 39858 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 40478 388226
rect 39858 388102 40478 388170
rect 39858 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 40478 388102
rect 39858 387978 40478 388046
rect 39858 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 40478 387978
rect 39858 370350 40478 387922
rect 39858 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 40478 370350
rect 39858 370226 40478 370294
rect 39858 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 40478 370226
rect 39858 370102 40478 370170
rect 39858 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 40478 370102
rect 39858 369978 40478 370046
rect 39858 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 40478 369978
rect 39858 352350 40478 369922
rect 66858 472350 67478 484408
rect 66858 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 67478 472350
rect 66858 472226 67478 472294
rect 66858 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 67478 472226
rect 66858 472102 67478 472170
rect 66858 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 67478 472102
rect 66858 471978 67478 472046
rect 66858 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 67478 471978
rect 66858 454350 67478 471922
rect 66858 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 67478 454350
rect 66858 454226 67478 454294
rect 66858 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 67478 454226
rect 66858 454102 67478 454170
rect 66858 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 67478 454102
rect 66858 453978 67478 454046
rect 66858 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 67478 453978
rect 66858 436350 67478 453922
rect 66858 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 67478 436350
rect 66858 436226 67478 436294
rect 66858 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 67478 436226
rect 66858 436102 67478 436170
rect 66858 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 67478 436102
rect 66858 435978 67478 436046
rect 66858 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 67478 435978
rect 66858 418350 67478 435922
rect 66858 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 67478 418350
rect 66858 418226 67478 418294
rect 66858 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 67478 418226
rect 66858 418102 67478 418170
rect 66858 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 67478 418102
rect 66858 417978 67478 418046
rect 66858 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 67478 417978
rect 66858 400350 67478 417922
rect 66858 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 67478 400350
rect 66858 400226 67478 400294
rect 66858 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 67478 400226
rect 66858 400102 67478 400170
rect 66858 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 67478 400102
rect 66858 399978 67478 400046
rect 66858 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 67478 399978
rect 66858 382350 67478 399922
rect 66858 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 67478 382350
rect 66858 382226 67478 382294
rect 66858 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 67478 382226
rect 66858 382102 67478 382170
rect 66858 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 67478 382102
rect 66858 381978 67478 382046
rect 66858 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 67478 381978
rect 39858 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 40478 352350
rect 39858 352226 40478 352294
rect 39858 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 40478 352226
rect 39858 352102 40478 352170
rect 39858 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 40478 352102
rect 39858 351978 40478 352046
rect 39858 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 40478 351978
rect 39858 334350 40478 351922
rect 39858 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 40478 334350
rect 39858 334226 40478 334294
rect 39858 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 40478 334226
rect 39858 334102 40478 334170
rect 39858 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 40478 334102
rect 39858 333978 40478 334046
rect 39858 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 40478 333978
rect 39858 316350 40478 333922
rect 39858 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 40478 316350
rect 39858 316226 40478 316294
rect 39858 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 40478 316226
rect 39858 316102 40478 316170
rect 39858 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 40478 316102
rect 39858 315978 40478 316046
rect 39858 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 40478 315978
rect 39858 298350 40478 315922
rect 63756 366418 63812 366428
rect 63756 304052 63812 366362
rect 63756 303986 63812 303996
rect 66858 364350 67478 381922
rect 66858 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 67478 364350
rect 66858 364226 67478 364294
rect 66858 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 67478 364226
rect 66858 364102 67478 364170
rect 66858 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 67478 364102
rect 66858 363978 67478 364046
rect 66858 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 67478 363978
rect 66858 346350 67478 363922
rect 66858 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 67478 346350
rect 66858 346226 67478 346294
rect 66858 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 67478 346226
rect 66858 346102 67478 346170
rect 66858 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 67478 346102
rect 66858 345978 67478 346046
rect 66858 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 67478 345978
rect 66858 328350 67478 345922
rect 66858 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 67478 328350
rect 66858 328226 67478 328294
rect 66858 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 67478 328226
rect 66858 328102 67478 328170
rect 66858 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 67478 328102
rect 66858 327978 67478 328046
rect 66858 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 67478 327978
rect 66858 310350 67478 327922
rect 66858 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 67478 310350
rect 66858 310226 67478 310294
rect 66858 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 67478 310226
rect 66858 310102 67478 310170
rect 66858 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 67478 310102
rect 66858 309978 67478 310046
rect 66858 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 67478 309978
rect 39858 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298294 40478 298350
rect 39858 298226 40478 298294
rect 39858 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298170 40478 298226
rect 39858 298102 40478 298170
rect 39858 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 40478 298102
rect 66858 298094 67478 309922
rect 70578 478350 71198 480728
rect 70578 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 71198 478350
rect 70578 478226 71198 478294
rect 70578 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 71198 478226
rect 77920 478308 79040 478360
rect 77920 478252 77956 478308
rect 78012 478252 78080 478308
rect 78136 478252 78204 478308
rect 78260 478252 78328 478308
rect 78384 478252 78452 478308
rect 78508 478252 78576 478308
rect 78632 478252 78700 478308
rect 78756 478252 78824 478308
rect 78880 478252 78948 478308
rect 79004 478252 79040 478308
rect 77920 478200 79040 478252
rect 70578 478102 71198 478170
rect 70578 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 71198 478102
rect 70578 477978 71198 478046
rect 70578 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 71198 477978
rect 70578 460350 71198 477922
rect 78560 477988 79040 478040
rect 78560 477932 78586 477988
rect 78642 477932 78710 477988
rect 78766 477932 78834 477988
rect 78890 477932 78958 477988
rect 79014 477932 79040 477988
rect 78560 477880 79040 477932
rect 70578 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 71198 460350
rect 70578 460226 71198 460294
rect 70578 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 71198 460226
rect 70578 460102 71198 460170
rect 70578 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 71198 460102
rect 70578 459978 71198 460046
rect 70578 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 71198 459978
rect 70578 442350 71198 459922
rect 70578 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 71198 442350
rect 70578 442226 71198 442294
rect 70578 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 71198 442226
rect 70578 442102 71198 442170
rect 70578 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 71198 442102
rect 70578 441978 71198 442046
rect 70578 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 71198 441978
rect 70578 424350 71198 441922
rect 70578 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 71198 424350
rect 70578 424226 71198 424294
rect 70578 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 71198 424226
rect 70578 424102 71198 424170
rect 70578 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 71198 424102
rect 70578 423978 71198 424046
rect 70578 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 71198 423978
rect 70578 406350 71198 423922
rect 70578 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 71198 406350
rect 70578 406226 71198 406294
rect 70578 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 71198 406226
rect 70578 406102 71198 406170
rect 70578 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 71198 406102
rect 70578 405978 71198 406046
rect 70578 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 71198 405978
rect 70578 388350 71198 405922
rect 70578 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 71198 388350
rect 70578 388226 71198 388294
rect 70578 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 71198 388226
rect 70578 388102 71198 388170
rect 70578 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 71198 388102
rect 70578 387978 71198 388046
rect 70578 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 71198 387978
rect 70578 370350 71198 387922
rect 70578 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 71198 370350
rect 70578 370226 71198 370294
rect 70578 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 71198 370226
rect 70578 370102 71198 370170
rect 70578 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 71198 370102
rect 70578 369978 71198 370046
rect 70578 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 71198 369978
rect 70578 352350 71198 369922
rect 97578 472350 98198 473048
rect 97578 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 98198 472350
rect 97578 472226 98198 472294
rect 97578 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 98198 472226
rect 97578 472102 98198 472170
rect 97578 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 98198 472102
rect 97578 471978 98198 472046
rect 97578 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 98198 471978
rect 97578 454350 98198 471922
rect 97578 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 98198 454350
rect 97578 454226 98198 454294
rect 97578 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 98198 454226
rect 97578 454102 98198 454170
rect 97578 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 98198 454102
rect 97578 453978 98198 454046
rect 97578 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 98198 453978
rect 97578 436350 98198 453922
rect 97578 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 98198 436350
rect 97578 436226 98198 436294
rect 97578 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 98198 436226
rect 97578 436102 98198 436170
rect 97578 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 98198 436102
rect 97578 435978 98198 436046
rect 97578 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 98198 435978
rect 97578 418350 98198 435922
rect 97578 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 98198 418350
rect 97578 418226 98198 418294
rect 97578 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 98198 418226
rect 97578 418102 98198 418170
rect 97578 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 98198 418102
rect 97578 417978 98198 418046
rect 97578 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 98198 417978
rect 97578 400350 98198 417922
rect 97578 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 98198 400350
rect 97578 400226 98198 400294
rect 97578 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 98198 400226
rect 97578 400102 98198 400170
rect 97578 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 98198 400102
rect 97578 399978 98198 400046
rect 97578 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 98198 399978
rect 97578 382350 98198 399922
rect 101298 460350 101918 473528
rect 101298 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 101918 460350
rect 101298 460226 101918 460294
rect 101298 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 101918 460226
rect 101298 460102 101918 460170
rect 101298 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 101918 460102
rect 101298 459978 101918 460046
rect 101298 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 101918 459978
rect 101298 442350 101918 459922
rect 101298 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 101918 442350
rect 101298 442226 101918 442294
rect 101298 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 101918 442226
rect 101298 442102 101918 442170
rect 101298 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 101918 442102
rect 101298 441978 101918 442046
rect 101298 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 101918 441978
rect 101298 424350 101918 441922
rect 101298 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 101918 424350
rect 101298 424226 101918 424294
rect 101298 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 101918 424226
rect 101298 424102 101918 424170
rect 101298 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 101918 424102
rect 101298 423978 101918 424046
rect 101298 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 101918 423978
rect 101298 406350 101918 423922
rect 101298 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 101918 406350
rect 101298 406226 101918 406294
rect 101298 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 101918 406226
rect 101298 406102 101918 406170
rect 101298 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 101918 406102
rect 101298 405978 101918 406046
rect 101298 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 101918 405978
rect 101298 388350 101918 405922
rect 101298 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 101918 388350
rect 101298 388226 101918 388294
rect 101298 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 101918 388226
rect 101298 388102 101918 388170
rect 101298 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 101918 388102
rect 101298 387978 101918 388046
rect 101298 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 101918 387978
rect 97578 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 98198 382350
rect 97578 382226 98198 382294
rect 97578 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 98198 382226
rect 97578 382102 98198 382170
rect 97578 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 98198 382102
rect 97578 381978 98198 382046
rect 97578 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 98198 381978
rect 93996 367138 94052 367148
rect 70578 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 71198 352350
rect 70578 352226 71198 352294
rect 70578 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 71198 352226
rect 70578 352102 71198 352170
rect 70578 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 71198 352102
rect 70578 351978 71198 352046
rect 70578 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 71198 351978
rect 70578 334350 71198 351922
rect 70578 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 71198 334350
rect 70578 334226 71198 334294
rect 70578 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 71198 334226
rect 70578 334102 71198 334170
rect 70578 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 71198 334102
rect 70578 333978 71198 334046
rect 70578 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 71198 333978
rect 70578 316350 71198 333922
rect 70578 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 71198 316350
rect 70578 316226 71198 316294
rect 70578 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 71198 316226
rect 70578 316102 71198 316170
rect 70578 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 71198 316102
rect 70578 315978 71198 316046
rect 70578 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 71198 315978
rect 70578 298422 71198 315922
rect 78876 365878 78932 365888
rect 78876 304052 78932 365822
rect 78876 303986 78932 303996
rect 93996 304052 94052 367082
rect 93996 303986 94052 303996
rect 97578 364350 98198 381922
rect 97578 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 98198 364350
rect 97578 364226 98198 364294
rect 97578 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 98198 364226
rect 97578 364102 98198 364170
rect 97578 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 98198 364102
rect 97578 363978 98198 364046
rect 97578 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 98198 363978
rect 97578 346350 98198 363922
rect 97578 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 98198 346350
rect 97578 346226 98198 346294
rect 97578 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 98198 346226
rect 97578 346102 98198 346170
rect 97578 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 98198 346102
rect 97578 345978 98198 346046
rect 97578 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 98198 345978
rect 97578 328350 98198 345922
rect 97578 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 98198 328350
rect 97578 328226 98198 328294
rect 97578 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 98198 328226
rect 97578 328102 98198 328170
rect 97578 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 98198 328102
rect 97578 327978 98198 328046
rect 97578 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 98198 327978
rect 97578 310350 98198 327922
rect 97578 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 98198 310350
rect 97578 310226 98198 310294
rect 97578 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 98198 310226
rect 97578 310102 98198 310170
rect 97578 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 98198 310102
rect 97578 309978 98198 310046
rect 97578 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 98198 309978
rect 70578 298366 70674 298422
rect 70730 298366 70798 298422
rect 70854 298366 70922 298422
rect 70978 298366 71046 298422
rect 71102 298366 71198 298422
rect 70578 298298 71198 298366
rect 70578 298242 70674 298298
rect 70730 298242 70798 298298
rect 70854 298242 70922 298298
rect 70978 298242 71046 298298
rect 71102 298242 71198 298298
rect 70578 298174 71198 298242
rect 70578 298118 70674 298174
rect 70730 298118 70798 298174
rect 70854 298118 70922 298174
rect 70978 298118 71046 298174
rect 71102 298118 71198 298174
rect 70578 298094 71198 298118
rect 39858 297978 40478 298046
rect 39858 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 40478 297978
rect 39858 280350 40478 297922
rect 44448 292350 44768 292384
rect 44448 292294 44518 292350
rect 44574 292294 44642 292350
rect 44698 292294 44768 292350
rect 44448 292226 44768 292294
rect 44448 292170 44518 292226
rect 44574 292170 44642 292226
rect 44698 292170 44768 292226
rect 44448 292102 44768 292170
rect 44448 292046 44518 292102
rect 44574 292046 44642 292102
rect 44698 292046 44768 292102
rect 44448 291978 44768 292046
rect 44448 291922 44518 291978
rect 44574 291922 44642 291978
rect 44698 291922 44768 291978
rect 44448 291888 44768 291922
rect 75168 292350 75488 292384
rect 75168 292294 75238 292350
rect 75294 292294 75362 292350
rect 75418 292294 75488 292350
rect 75168 292226 75488 292294
rect 75168 292170 75238 292226
rect 75294 292170 75362 292226
rect 75418 292170 75488 292226
rect 75168 292102 75488 292170
rect 75168 292046 75238 292102
rect 75294 292046 75362 292102
rect 75418 292046 75488 292102
rect 75168 291978 75488 292046
rect 75168 291922 75238 291978
rect 75294 291922 75362 291978
rect 75418 291922 75488 291978
rect 75168 291888 75488 291922
rect 97578 292350 98198 309922
rect 97578 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 98198 292350
rect 97578 292226 98198 292294
rect 97578 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 98198 292226
rect 97578 292102 98198 292170
rect 97578 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 98198 292102
rect 97578 291978 98198 292046
rect 97578 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 98198 291978
rect 39858 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 40478 280350
rect 39858 280226 40478 280294
rect 39858 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 40478 280226
rect 39858 280102 40478 280170
rect 39858 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 40478 280102
rect 39858 279978 40478 280046
rect 39858 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 40478 279978
rect 39858 262350 40478 279922
rect 59808 280350 60128 280384
rect 59808 280294 59878 280350
rect 59934 280294 60002 280350
rect 60058 280294 60128 280350
rect 59808 280226 60128 280294
rect 59808 280170 59878 280226
rect 59934 280170 60002 280226
rect 60058 280170 60128 280226
rect 59808 280102 60128 280170
rect 59808 280046 59878 280102
rect 59934 280046 60002 280102
rect 60058 280046 60128 280102
rect 59808 279978 60128 280046
rect 59808 279922 59878 279978
rect 59934 279922 60002 279978
rect 60058 279922 60128 279978
rect 59808 279888 60128 279922
rect 90528 280350 90848 280384
rect 90528 280294 90598 280350
rect 90654 280294 90722 280350
rect 90778 280294 90848 280350
rect 90528 280226 90848 280294
rect 90528 280170 90598 280226
rect 90654 280170 90722 280226
rect 90778 280170 90848 280226
rect 90528 280102 90848 280170
rect 90528 280046 90598 280102
rect 90654 280046 90722 280102
rect 90778 280046 90848 280102
rect 90528 279978 90848 280046
rect 90528 279922 90598 279978
rect 90654 279922 90722 279978
rect 90778 279922 90848 279978
rect 90528 279888 90848 279922
rect 44448 274350 44768 274384
rect 44448 274294 44518 274350
rect 44574 274294 44642 274350
rect 44698 274294 44768 274350
rect 44448 274226 44768 274294
rect 44448 274170 44518 274226
rect 44574 274170 44642 274226
rect 44698 274170 44768 274226
rect 44448 274102 44768 274170
rect 44448 274046 44518 274102
rect 44574 274046 44642 274102
rect 44698 274046 44768 274102
rect 44448 273978 44768 274046
rect 44448 273922 44518 273978
rect 44574 273922 44642 273978
rect 44698 273922 44768 273978
rect 44448 273888 44768 273922
rect 75168 274350 75488 274384
rect 75168 274294 75238 274350
rect 75294 274294 75362 274350
rect 75418 274294 75488 274350
rect 75168 274226 75488 274294
rect 75168 274170 75238 274226
rect 75294 274170 75362 274226
rect 75418 274170 75488 274226
rect 75168 274102 75488 274170
rect 75168 274046 75238 274102
rect 75294 274046 75362 274102
rect 75418 274046 75488 274102
rect 75168 273978 75488 274046
rect 75168 273922 75238 273978
rect 75294 273922 75362 273978
rect 75418 273922 75488 273978
rect 75168 273888 75488 273922
rect 97578 274350 98198 291922
rect 97578 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 98198 274350
rect 97578 274226 98198 274294
rect 97578 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 98198 274226
rect 97578 274102 98198 274170
rect 97578 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 98198 274102
rect 97578 273978 98198 274046
rect 97578 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 98198 273978
rect 39858 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 40478 262350
rect 39858 262226 40478 262294
rect 39858 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 40478 262226
rect 39858 262102 40478 262170
rect 39858 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 40478 262102
rect 39858 261978 40478 262046
rect 39858 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 40478 261978
rect 39858 244350 40478 261922
rect 59808 262350 60128 262384
rect 59808 262294 59878 262350
rect 59934 262294 60002 262350
rect 60058 262294 60128 262350
rect 59808 262226 60128 262294
rect 59808 262170 59878 262226
rect 59934 262170 60002 262226
rect 60058 262170 60128 262226
rect 59808 262102 60128 262170
rect 59808 262046 59878 262102
rect 59934 262046 60002 262102
rect 60058 262046 60128 262102
rect 59808 261978 60128 262046
rect 59808 261922 59878 261978
rect 59934 261922 60002 261978
rect 60058 261922 60128 261978
rect 59808 261888 60128 261922
rect 90528 262350 90848 262384
rect 90528 262294 90598 262350
rect 90654 262294 90722 262350
rect 90778 262294 90848 262350
rect 90528 262226 90848 262294
rect 90528 262170 90598 262226
rect 90654 262170 90722 262226
rect 90778 262170 90848 262226
rect 90528 262102 90848 262170
rect 90528 262046 90598 262102
rect 90654 262046 90722 262102
rect 90778 262046 90848 262102
rect 90528 261978 90848 262046
rect 90528 261922 90598 261978
rect 90654 261922 90722 261978
rect 90778 261922 90848 261978
rect 90528 261888 90848 261922
rect 44448 256350 44768 256384
rect 44448 256294 44518 256350
rect 44574 256294 44642 256350
rect 44698 256294 44768 256350
rect 44448 256226 44768 256294
rect 44448 256170 44518 256226
rect 44574 256170 44642 256226
rect 44698 256170 44768 256226
rect 44448 256102 44768 256170
rect 44448 256046 44518 256102
rect 44574 256046 44642 256102
rect 44698 256046 44768 256102
rect 44448 255978 44768 256046
rect 44448 255922 44518 255978
rect 44574 255922 44642 255978
rect 44698 255922 44768 255978
rect 44448 255888 44768 255922
rect 75168 256350 75488 256384
rect 75168 256294 75238 256350
rect 75294 256294 75362 256350
rect 75418 256294 75488 256350
rect 75168 256226 75488 256294
rect 75168 256170 75238 256226
rect 75294 256170 75362 256226
rect 75418 256170 75488 256226
rect 75168 256102 75488 256170
rect 75168 256046 75238 256102
rect 75294 256046 75362 256102
rect 75418 256046 75488 256102
rect 75168 255978 75488 256046
rect 75168 255922 75238 255978
rect 75294 255922 75362 255978
rect 75418 255922 75488 255978
rect 75168 255888 75488 255922
rect 97578 256350 98198 273922
rect 97578 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 98198 256350
rect 97578 256226 98198 256294
rect 97578 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 98198 256226
rect 97578 256102 98198 256170
rect 97578 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 98198 256102
rect 97578 255978 98198 256046
rect 97578 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 98198 255978
rect 39858 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 40478 244350
rect 39858 244226 40478 244294
rect 39858 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 40478 244226
rect 39858 244102 40478 244170
rect 39858 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 40478 244102
rect 39858 243978 40478 244046
rect 39858 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 40478 243978
rect 39858 226350 40478 243922
rect 46172 247078 46228 247088
rect 46172 236068 46228 247022
rect 59808 244350 60128 244384
rect 59808 244294 59878 244350
rect 59934 244294 60002 244350
rect 60058 244294 60128 244350
rect 59808 244226 60128 244294
rect 59808 244170 59878 244226
rect 59934 244170 60002 244226
rect 60058 244170 60128 244226
rect 59808 244102 60128 244170
rect 59808 244046 59878 244102
rect 59934 244046 60002 244102
rect 60058 244046 60128 244102
rect 59808 243978 60128 244046
rect 59808 243922 59878 243978
rect 59934 243922 60002 243978
rect 60058 243922 60128 243978
rect 59808 243888 60128 243922
rect 48524 240212 48580 240222
rect 46172 236002 46228 236012
rect 46956 236180 47012 236190
rect 39858 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 40478 226350
rect 39858 226226 40478 226294
rect 39858 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 40478 226226
rect 39858 226102 40478 226170
rect 39858 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 40478 226102
rect 39858 225978 40478 226046
rect 39858 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 40478 225978
rect 36138 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 36758 202350
rect 36138 202226 36758 202294
rect 36138 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 36758 202226
rect 36138 202102 36758 202170
rect 36138 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 36758 202102
rect 36138 201978 36758 202046
rect 36138 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 36758 201978
rect 36138 184350 36758 201922
rect 36138 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 36758 184350
rect 36138 184226 36758 184294
rect 36138 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 36758 184226
rect 36138 184102 36758 184170
rect 36138 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 36758 184102
rect 36138 183978 36758 184046
rect 36138 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 36758 183978
rect 36138 166350 36758 183922
rect 36138 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 36758 166350
rect 36138 166226 36758 166294
rect 36138 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 36758 166226
rect 36138 166102 36758 166170
rect 36138 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 36758 166102
rect 36138 165978 36758 166046
rect 36138 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 36758 165978
rect 36138 148350 36758 165922
rect 36138 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 36758 148350
rect 36138 148226 36758 148294
rect 36138 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 36758 148226
rect 36138 148102 36758 148170
rect 36138 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 36758 148102
rect 36138 147978 36758 148046
rect 36138 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 36758 147978
rect 36138 130350 36758 147922
rect 36138 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 36758 130350
rect 36138 130226 36758 130294
rect 36138 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 36758 130226
rect 36138 130102 36758 130170
rect 36138 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 36758 130102
rect 36138 129978 36758 130046
rect 36138 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 36758 129978
rect 36138 112350 36758 129922
rect 36138 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 36758 112350
rect 36138 112226 36758 112294
rect 36138 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 36758 112226
rect 36138 112102 36758 112170
rect 36138 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 36758 112102
rect 36138 111978 36758 112046
rect 36138 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 36758 111978
rect 36138 94350 36758 111922
rect 36138 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 36758 94350
rect 36138 94226 36758 94294
rect 36138 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 36758 94226
rect 36138 94102 36758 94170
rect 36138 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 36758 94102
rect 36138 93978 36758 94046
rect 36138 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 36758 93978
rect 36138 76350 36758 93922
rect 36138 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 36758 76350
rect 36138 76226 36758 76294
rect 36138 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 36758 76226
rect 36138 76102 36758 76170
rect 36138 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 36758 76102
rect 36138 75978 36758 76046
rect 36138 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 36758 75978
rect 36138 58350 36758 75922
rect 36138 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 36758 58350
rect 36138 58226 36758 58294
rect 36138 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 36758 58226
rect 36138 58102 36758 58170
rect 36138 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 36758 58102
rect 36138 57978 36758 58046
rect 36138 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 36758 57978
rect 36138 40350 36758 57922
rect 36138 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 36758 40350
rect 36138 40226 36758 40294
rect 36138 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 36758 40226
rect 36138 40102 36758 40170
rect 36138 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 36758 40102
rect 36138 39978 36758 40046
rect 36138 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 36758 39978
rect 36138 22350 36758 39922
rect 36138 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 36758 22350
rect 36138 22226 36758 22294
rect 36138 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 36758 22226
rect 36138 22102 36758 22170
rect 36138 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 36758 22102
rect 36138 21978 36758 22046
rect 36138 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 36758 21978
rect 36138 4350 36758 21922
rect 39676 212548 39732 212558
rect 39676 4978 39732 212492
rect 39676 4912 39732 4922
rect 39858 208350 40478 225922
rect 39858 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 40478 208350
rect 39858 208226 40478 208294
rect 39858 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 40478 208226
rect 39858 208102 40478 208170
rect 39858 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 40478 208102
rect 39858 207978 40478 208046
rect 39858 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 40478 207978
rect 39858 190350 40478 207922
rect 39858 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 40478 190350
rect 39858 190226 40478 190294
rect 39858 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 40478 190226
rect 39858 190102 40478 190170
rect 39858 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 40478 190102
rect 39858 189978 40478 190046
rect 39858 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 40478 189978
rect 39858 172350 40478 189922
rect 39858 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 40478 172350
rect 39858 172226 40478 172294
rect 39858 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 40478 172226
rect 39858 172102 40478 172170
rect 39858 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 40478 172102
rect 39858 171978 40478 172046
rect 39858 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 40478 171978
rect 39858 154350 40478 171922
rect 39858 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 40478 154350
rect 39858 154226 40478 154294
rect 39858 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 40478 154226
rect 39858 154102 40478 154170
rect 39858 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 40478 154102
rect 39858 153978 40478 154046
rect 39858 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 40478 153978
rect 39858 136350 40478 153922
rect 39858 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 40478 136350
rect 39858 136226 40478 136294
rect 39858 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 40478 136226
rect 39858 136102 40478 136170
rect 39858 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 40478 136102
rect 39858 135978 40478 136046
rect 39858 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 40478 135978
rect 39858 118350 40478 135922
rect 39858 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 40478 118350
rect 39858 118226 40478 118294
rect 39858 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 40478 118226
rect 39858 118102 40478 118170
rect 39858 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 40478 118102
rect 39858 117978 40478 118046
rect 39858 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 40478 117978
rect 39858 100350 40478 117922
rect 39858 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 40478 100350
rect 39858 100226 40478 100294
rect 39858 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 40478 100226
rect 39858 100102 40478 100170
rect 39858 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 40478 100102
rect 39858 99978 40478 100046
rect 39858 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 40478 99978
rect 39858 82350 40478 99922
rect 39858 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 40478 82350
rect 39858 82226 40478 82294
rect 39858 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 40478 82226
rect 39858 82102 40478 82170
rect 39858 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 40478 82102
rect 39858 81978 40478 82046
rect 39858 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 40478 81978
rect 39858 64350 40478 81922
rect 39858 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 40478 64350
rect 39858 64226 40478 64294
rect 39858 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 40478 64226
rect 39858 64102 40478 64170
rect 39858 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 40478 64102
rect 39858 63978 40478 64046
rect 39858 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 40478 63978
rect 39858 46350 40478 63922
rect 39858 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 40478 46350
rect 39858 46226 40478 46294
rect 39858 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 40478 46226
rect 39858 46102 40478 46170
rect 39858 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 40478 46102
rect 39858 45978 40478 46046
rect 39858 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 40478 45978
rect 39858 28350 40478 45922
rect 39858 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 40478 28350
rect 39858 28226 40478 28294
rect 39858 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 40478 28226
rect 39858 28102 40478 28170
rect 39858 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 40478 28102
rect 39858 27978 40478 28046
rect 39858 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 40478 27978
rect 39858 10350 40478 27922
rect 39858 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 40478 10350
rect 39858 10226 40478 10294
rect 39858 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 40478 10226
rect 39858 10102 40478 10170
rect 39858 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 40478 10102
rect 39858 9978 40478 10046
rect 39858 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 40478 9978
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 35084 4162 35140 4172
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 9138 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 9758 -1120
rect 9138 -1244 9758 -1176
rect 9138 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 9758 -1244
rect 9138 -1368 9758 -1300
rect 9138 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 9758 -1368
rect 9138 -1492 9758 -1424
rect 9138 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 9758 -1492
rect 9138 -1644 9758 -1548
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 39858 -1120 40478 9922
rect 41356 234478 41412 234488
rect 41356 4900 41412 234422
rect 44448 202350 44768 202384
rect 44448 202294 44518 202350
rect 44574 202294 44642 202350
rect 44698 202294 44768 202350
rect 44448 202226 44768 202294
rect 44448 202170 44518 202226
rect 44574 202170 44642 202226
rect 44698 202170 44768 202226
rect 44448 202102 44768 202170
rect 44448 202046 44518 202102
rect 44574 202046 44642 202102
rect 44698 202046 44768 202102
rect 44448 201978 44768 202046
rect 44448 201922 44518 201978
rect 44574 201922 44642 201978
rect 44698 201922 44768 201978
rect 44448 201888 44768 201922
rect 44448 184350 44768 184384
rect 44448 184294 44518 184350
rect 44574 184294 44642 184350
rect 44698 184294 44768 184350
rect 44448 184226 44768 184294
rect 44448 184170 44518 184226
rect 44574 184170 44642 184226
rect 44698 184170 44768 184226
rect 44448 184102 44768 184170
rect 44448 184046 44518 184102
rect 44574 184046 44642 184102
rect 44698 184046 44768 184102
rect 44448 183978 44768 184046
rect 44448 183922 44518 183978
rect 44574 183922 44642 183978
rect 44698 183922 44768 183978
rect 44448 183888 44768 183922
rect 44448 166350 44768 166384
rect 44448 166294 44518 166350
rect 44574 166294 44642 166350
rect 44698 166294 44768 166350
rect 44448 166226 44768 166294
rect 44448 166170 44518 166226
rect 44574 166170 44642 166226
rect 44698 166170 44768 166226
rect 44448 166102 44768 166170
rect 44448 166046 44518 166102
rect 44574 166046 44642 166102
rect 44698 166046 44768 166102
rect 44448 165978 44768 166046
rect 44448 165922 44518 165978
rect 44574 165922 44642 165978
rect 44698 165922 44768 165978
rect 44448 165888 44768 165922
rect 44448 148350 44768 148384
rect 44448 148294 44518 148350
rect 44574 148294 44642 148350
rect 44698 148294 44768 148350
rect 44448 148226 44768 148294
rect 44448 148170 44518 148226
rect 44574 148170 44642 148226
rect 44698 148170 44768 148226
rect 44448 148102 44768 148170
rect 44448 148046 44518 148102
rect 44574 148046 44642 148102
rect 44698 148046 44768 148102
rect 44448 147978 44768 148046
rect 44448 147922 44518 147978
rect 44574 147922 44642 147978
rect 44698 147922 44768 147978
rect 44448 147888 44768 147922
rect 44448 130350 44768 130384
rect 44448 130294 44518 130350
rect 44574 130294 44642 130350
rect 44698 130294 44768 130350
rect 44448 130226 44768 130294
rect 44448 130170 44518 130226
rect 44574 130170 44642 130226
rect 44698 130170 44768 130226
rect 44448 130102 44768 130170
rect 44448 130046 44518 130102
rect 44574 130046 44642 130102
rect 44698 130046 44768 130102
rect 44448 129978 44768 130046
rect 44448 129922 44518 129978
rect 44574 129922 44642 129978
rect 44698 129922 44768 129978
rect 44448 129888 44768 129922
rect 44448 112350 44768 112384
rect 44448 112294 44518 112350
rect 44574 112294 44642 112350
rect 44698 112294 44768 112350
rect 44448 112226 44768 112294
rect 44448 112170 44518 112226
rect 44574 112170 44642 112226
rect 44698 112170 44768 112226
rect 44448 112102 44768 112170
rect 44448 112046 44518 112102
rect 44574 112046 44642 112102
rect 44698 112046 44768 112102
rect 44448 111978 44768 112046
rect 44448 111922 44518 111978
rect 44574 111922 44642 111978
rect 44698 111922 44768 111978
rect 44448 111888 44768 111922
rect 44448 94350 44768 94384
rect 44448 94294 44518 94350
rect 44574 94294 44642 94350
rect 44698 94294 44768 94350
rect 44448 94226 44768 94294
rect 44448 94170 44518 94226
rect 44574 94170 44642 94226
rect 44698 94170 44768 94226
rect 44448 94102 44768 94170
rect 44448 94046 44518 94102
rect 44574 94046 44642 94102
rect 44698 94046 44768 94102
rect 44448 93978 44768 94046
rect 44448 93922 44518 93978
rect 44574 93922 44642 93978
rect 44698 93922 44768 93978
rect 44448 93888 44768 93922
rect 44448 76350 44768 76384
rect 44448 76294 44518 76350
rect 44574 76294 44642 76350
rect 44698 76294 44768 76350
rect 44448 76226 44768 76294
rect 44448 76170 44518 76226
rect 44574 76170 44642 76226
rect 44698 76170 44768 76226
rect 44448 76102 44768 76170
rect 44448 76046 44518 76102
rect 44574 76046 44642 76102
rect 44698 76046 44768 76102
rect 44448 75978 44768 76046
rect 44448 75922 44518 75978
rect 44574 75922 44642 75978
rect 44698 75922 44768 75978
rect 44448 75888 44768 75922
rect 44448 58350 44768 58384
rect 44448 58294 44518 58350
rect 44574 58294 44642 58350
rect 44698 58294 44768 58350
rect 44448 58226 44768 58294
rect 44448 58170 44518 58226
rect 44574 58170 44642 58226
rect 44698 58170 44768 58226
rect 44448 58102 44768 58170
rect 44448 58046 44518 58102
rect 44574 58046 44642 58102
rect 44698 58046 44768 58102
rect 44448 57978 44768 58046
rect 44448 57922 44518 57978
rect 44574 57922 44642 57978
rect 44698 57922 44768 57978
rect 44448 57888 44768 57922
rect 46956 49588 47012 236124
rect 46956 49522 47012 49532
rect 48524 48244 48580 240156
rect 66858 238350 67478 245074
rect 66858 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 67478 238350
rect 66858 238226 67478 238294
rect 66858 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 67478 238226
rect 66858 238102 67478 238170
rect 66858 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 67478 238102
rect 66858 237978 67478 238046
rect 66858 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 67478 237978
rect 51772 234612 51828 234622
rect 50204 234500 50260 234510
rect 48524 48178 48580 48188
rect 48636 224532 48692 224542
rect 41356 4834 41412 4844
rect 48636 4228 48692 224476
rect 49644 211764 49700 211774
rect 49532 210084 49588 210094
rect 49532 164638 49588 210028
rect 49644 206578 49700 211708
rect 49644 206512 49700 206522
rect 49532 164572 49588 164582
rect 50204 48020 50260 234444
rect 50204 47954 50260 47964
rect 50316 216020 50372 216030
rect 50316 4788 50372 215964
rect 51772 48132 51828 234556
rect 51996 224308 52052 224318
rect 51772 48066 51828 48076
rect 51884 217588 51940 217598
rect 51884 5012 51940 217532
rect 51884 4946 51940 4956
rect 50316 4722 50372 4732
rect 51996 4340 52052 224252
rect 66858 220350 67478 237922
rect 66858 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 67478 220350
rect 66858 220226 67478 220294
rect 66858 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 67478 220226
rect 66858 220102 67478 220170
rect 66858 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 67478 220102
rect 66858 219978 67478 220046
rect 66858 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 67478 219978
rect 66858 210462 67478 219922
rect 70578 244350 71198 245074
rect 70578 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 71198 244350
rect 70578 244226 71198 244294
rect 70578 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 71198 244226
rect 70578 244102 71198 244170
rect 70578 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 71198 244102
rect 70578 243978 71198 244046
rect 70578 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 71198 243978
rect 70578 226350 71198 243922
rect 90528 244350 90848 244384
rect 90528 244294 90598 244350
rect 90654 244294 90722 244350
rect 90778 244294 90848 244350
rect 90528 244226 90848 244294
rect 90528 244170 90598 244226
rect 90654 244170 90722 244226
rect 90778 244170 90848 244226
rect 90528 244102 90848 244170
rect 90528 244046 90598 244102
rect 90654 244046 90722 244102
rect 90778 244046 90848 244102
rect 90528 243978 90848 244046
rect 90528 243922 90598 243978
rect 90654 243922 90722 243978
rect 90778 243922 90848 243978
rect 90528 243888 90848 243922
rect 72940 238532 72996 238542
rect 72940 237538 72996 238476
rect 76972 238532 77028 238542
rect 76972 237718 77028 238476
rect 97578 238350 98198 255922
rect 96572 238308 96628 238318
rect 97020 238308 97076 238318
rect 96628 238252 97020 238258
rect 96572 238202 97076 238252
rect 97578 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 98198 238350
rect 97578 238226 98198 238294
rect 76972 237652 77028 237662
rect 97578 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 98198 238226
rect 97578 238102 98198 238170
rect 97578 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 98198 238102
rect 97578 237978 98198 238046
rect 97578 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 98198 237978
rect 72940 237472 72996 237482
rect 70578 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 71198 226350
rect 70578 226226 71198 226294
rect 70578 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 71198 226226
rect 70578 226102 71198 226170
rect 70578 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 71198 226102
rect 70578 225978 71198 226046
rect 70578 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 71198 225978
rect 70578 210462 71198 225922
rect 97578 220350 98198 237922
rect 99932 383460 99988 383470
rect 99932 237538 99988 383404
rect 99932 237472 99988 237482
rect 101298 370350 101918 387922
rect 128298 472350 128918 489922
rect 128298 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 128918 472350
rect 128298 472226 128918 472294
rect 128298 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 128918 472226
rect 128298 472102 128918 472170
rect 128298 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 128918 472102
rect 128298 471978 128918 472046
rect 128298 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 128918 471978
rect 128298 454350 128918 471922
rect 128298 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 128918 454350
rect 128298 454226 128918 454294
rect 128298 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 128918 454226
rect 128298 454102 128918 454170
rect 128298 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 128918 454102
rect 128298 453978 128918 454046
rect 128298 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 128918 453978
rect 128298 436350 128918 453922
rect 128298 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 128918 436350
rect 128298 436226 128918 436294
rect 128298 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 128918 436226
rect 128298 436102 128918 436170
rect 128298 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 128918 436102
rect 128298 435978 128918 436046
rect 128298 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 128918 435978
rect 128298 418350 128918 435922
rect 128298 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 128918 418350
rect 128298 418226 128918 418294
rect 128298 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 128918 418226
rect 128298 418102 128918 418170
rect 128298 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 128918 418102
rect 128298 417978 128918 418046
rect 128298 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 128918 417978
rect 128298 400350 128918 417922
rect 128298 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 128918 400350
rect 128298 400226 128918 400294
rect 128298 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 128918 400226
rect 128298 400102 128918 400170
rect 128298 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 128918 400102
rect 128298 399978 128918 400046
rect 128298 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 128918 399978
rect 101298 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 101918 370350
rect 101298 370226 101918 370294
rect 101298 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 101918 370226
rect 101298 370102 101918 370170
rect 101298 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 101918 370102
rect 101298 369978 101918 370046
rect 101298 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 101918 369978
rect 101298 352350 101918 369922
rect 101298 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 101918 352350
rect 101298 352226 101918 352294
rect 101298 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 101918 352226
rect 101298 352102 101918 352170
rect 101298 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 101918 352102
rect 101298 351978 101918 352046
rect 101298 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 101918 351978
rect 101298 334350 101918 351922
rect 101298 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 101918 334350
rect 101298 334226 101918 334294
rect 101298 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 101918 334226
rect 101298 334102 101918 334170
rect 101298 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 101918 334102
rect 101298 333978 101918 334046
rect 101298 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 101918 333978
rect 101298 316350 101918 333922
rect 101298 316294 101394 316350
rect 101450 316294 101518 316350
rect 101574 316294 101642 316350
rect 101698 316294 101766 316350
rect 101822 316294 101918 316350
rect 101298 316226 101918 316294
rect 101298 316170 101394 316226
rect 101450 316170 101518 316226
rect 101574 316170 101642 316226
rect 101698 316170 101766 316226
rect 101822 316170 101918 316226
rect 101298 316102 101918 316170
rect 101298 316046 101394 316102
rect 101450 316046 101518 316102
rect 101574 316046 101642 316102
rect 101698 316046 101766 316102
rect 101822 316046 101918 316102
rect 101298 315978 101918 316046
rect 101298 315922 101394 315978
rect 101450 315922 101518 315978
rect 101574 315922 101642 315978
rect 101698 315922 101766 315978
rect 101822 315922 101918 315978
rect 101298 298350 101918 315922
rect 101298 298294 101394 298350
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 101918 298350
rect 101298 298226 101918 298294
rect 101298 298170 101394 298226
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 101918 298226
rect 101298 298102 101918 298170
rect 101298 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 101918 298102
rect 101298 297978 101918 298046
rect 101298 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 101918 297978
rect 101298 280350 101918 297922
rect 101298 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 101918 280350
rect 101298 280226 101918 280294
rect 101298 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 101918 280226
rect 101298 280102 101918 280170
rect 101298 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 101918 280102
rect 101298 279978 101918 280046
rect 101298 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 101918 279978
rect 101298 262350 101918 279922
rect 101298 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 101918 262350
rect 101298 262226 101918 262294
rect 101298 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 101918 262226
rect 101298 262102 101918 262170
rect 101298 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 101918 262102
rect 101298 261978 101918 262046
rect 101298 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 101918 261978
rect 101298 244350 101918 261922
rect 101298 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 101918 244350
rect 101298 244226 101918 244294
rect 101298 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 101918 244226
rect 101298 244102 101918 244170
rect 101298 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 101918 244102
rect 101298 243978 101918 244046
rect 101298 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 101918 243978
rect 97578 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 98198 220350
rect 97578 220226 98198 220294
rect 97578 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 98198 220226
rect 97578 220102 98198 220170
rect 97578 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 98198 220102
rect 97578 219978 98198 220046
rect 97578 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 98198 219978
rect 97578 210462 98198 219922
rect 101298 226350 101918 243922
rect 110012 385252 110068 385262
rect 110012 237718 110068 385196
rect 128298 382350 128918 399922
rect 128298 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 128918 382350
rect 128298 382226 128918 382294
rect 128298 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 128918 382226
rect 128298 382102 128918 382170
rect 128298 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 128918 382102
rect 128298 381978 128918 382046
rect 128298 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 128918 381978
rect 128298 364350 128918 381922
rect 128298 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 128918 364350
rect 128298 364226 128918 364294
rect 128298 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 128918 364226
rect 128298 364102 128918 364170
rect 128298 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 128918 364102
rect 128298 363978 128918 364046
rect 128298 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 128918 363978
rect 128298 346350 128918 363922
rect 128298 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 128918 346350
rect 128298 346226 128918 346294
rect 128298 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 128918 346226
rect 128298 346102 128918 346170
rect 128298 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 128918 346102
rect 128298 345978 128918 346046
rect 128298 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 128918 345978
rect 128298 328350 128918 345922
rect 128298 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 128918 328350
rect 128298 328226 128918 328294
rect 128298 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 128918 328226
rect 128298 328102 128918 328170
rect 128298 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 128918 328102
rect 128298 327978 128918 328046
rect 128298 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 128918 327978
rect 128298 310350 128918 327922
rect 128298 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 128918 310350
rect 128298 310226 128918 310294
rect 128298 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 128918 310226
rect 128298 310102 128918 310170
rect 128298 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 128918 310102
rect 128298 309978 128918 310046
rect 128298 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 128918 309978
rect 128298 292350 128918 309922
rect 128298 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 128918 292350
rect 128298 292226 128918 292294
rect 128298 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 128918 292226
rect 128298 292102 128918 292170
rect 128298 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 128918 292102
rect 128298 291978 128918 292046
rect 128298 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 128918 291978
rect 121772 291844 121828 291854
rect 120092 287812 120148 287822
rect 110012 237652 110068 237662
rect 113372 286356 113428 286366
rect 101298 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 101918 226350
rect 101298 226226 101918 226294
rect 101298 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 101918 226226
rect 101298 226102 101918 226170
rect 101298 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 101918 226102
rect 101298 225978 101918 226046
rect 101298 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 101918 225978
rect 101298 210462 101918 225922
rect 113372 211092 113428 286300
rect 118412 285460 118468 285470
rect 118412 220276 118468 285404
rect 118412 220210 118468 220220
rect 120092 212772 120148 287756
rect 120092 212706 120148 212716
rect 113372 211026 113428 211036
rect 121772 210980 121828 291788
rect 121772 210914 121828 210924
rect 128298 274350 128918 291922
rect 128298 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 128918 274350
rect 128298 274226 128918 274294
rect 128298 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 128918 274226
rect 128298 274102 128918 274170
rect 128298 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 128918 274102
rect 128298 273978 128918 274046
rect 128298 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 128918 273978
rect 128298 256350 128918 273922
rect 128298 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 128918 256350
rect 128298 256226 128918 256294
rect 128298 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 128918 256226
rect 128298 256102 128918 256170
rect 128298 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 128918 256102
rect 128298 255978 128918 256046
rect 128298 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 128918 255978
rect 128298 238350 128918 255922
rect 128298 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 128918 238350
rect 128298 238226 128918 238294
rect 128298 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 128918 238226
rect 128298 238102 128918 238170
rect 128298 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 128918 238102
rect 128298 237978 128918 238046
rect 128298 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 128918 237978
rect 128298 220350 128918 237922
rect 128298 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 128918 220350
rect 128298 220226 128918 220294
rect 128298 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 128918 220226
rect 128298 220102 128918 220170
rect 128298 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 128918 220102
rect 128298 219978 128918 220046
rect 128298 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 128918 219978
rect 128298 210462 128918 219922
rect 132018 478350 132638 493368
rect 132018 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 132638 478350
rect 132018 478226 132638 478294
rect 132018 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 132638 478226
rect 132018 478102 132638 478170
rect 132018 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 132638 478102
rect 132018 477978 132638 478046
rect 132018 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 132638 477978
rect 132018 460350 132638 477922
rect 132018 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 132638 460350
rect 132018 460226 132638 460294
rect 132018 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 132638 460226
rect 132018 460102 132638 460170
rect 132018 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 132638 460102
rect 132018 459978 132638 460046
rect 132018 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 132638 459978
rect 132018 442350 132638 459922
rect 132018 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 132638 442350
rect 132018 442226 132638 442294
rect 132018 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 132638 442226
rect 132018 442102 132638 442170
rect 132018 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 132638 442102
rect 132018 441978 132638 442046
rect 132018 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 132638 441978
rect 132018 424350 132638 441922
rect 132018 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 132638 424350
rect 132018 424226 132638 424294
rect 132018 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 132638 424226
rect 132018 424102 132638 424170
rect 132018 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 132638 424102
rect 132018 423978 132638 424046
rect 132018 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 132638 423978
rect 132018 406350 132638 423922
rect 132018 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 132638 406350
rect 132018 406226 132638 406294
rect 132018 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 132638 406226
rect 132018 406102 132638 406170
rect 132018 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 132638 406102
rect 132018 405978 132638 406046
rect 132018 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 132638 405978
rect 132018 388350 132638 405922
rect 132018 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 132638 388350
rect 132018 388226 132638 388294
rect 132018 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 132638 388226
rect 132018 388102 132638 388170
rect 132018 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 132638 388102
rect 132018 387978 132638 388046
rect 132018 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 132638 387978
rect 132018 370350 132638 387922
rect 132018 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 132638 370350
rect 132018 370226 132638 370294
rect 132018 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 132638 370226
rect 132018 370102 132638 370170
rect 132018 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 132638 370102
rect 132018 369978 132638 370046
rect 132018 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 132638 369978
rect 132018 352350 132638 369922
rect 159018 490350 159638 507922
rect 159018 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 159638 490350
rect 159018 490226 159638 490294
rect 159018 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 159638 490226
rect 159018 490102 159638 490170
rect 159018 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 159638 490102
rect 159018 489978 159638 490046
rect 159018 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 159638 489978
rect 159018 472350 159638 489922
rect 159018 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 159638 472350
rect 159018 472226 159638 472294
rect 159018 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 159638 472226
rect 159018 472102 159638 472170
rect 159018 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 159638 472102
rect 159018 471978 159638 472046
rect 159018 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 159638 471978
rect 159018 454350 159638 471922
rect 159018 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 159638 454350
rect 159018 454226 159638 454294
rect 159018 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 159638 454226
rect 159018 454102 159638 454170
rect 159018 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 159638 454102
rect 159018 453978 159638 454046
rect 159018 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 159638 453978
rect 159018 436350 159638 453922
rect 159018 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 159638 436350
rect 159018 436226 159638 436294
rect 159018 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 159638 436226
rect 159018 436102 159638 436170
rect 159018 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 159638 436102
rect 159018 435978 159638 436046
rect 159018 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 159638 435978
rect 159018 418350 159638 435922
rect 159018 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 159638 418350
rect 159018 418226 159638 418294
rect 159018 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 159638 418226
rect 159018 418102 159638 418170
rect 159018 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 159638 418102
rect 159018 417978 159638 418046
rect 159018 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 159638 417978
rect 159018 400350 159638 417922
rect 159018 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 159638 400350
rect 159018 400226 159638 400294
rect 159018 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 159638 400226
rect 159018 400102 159638 400170
rect 159018 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 159638 400102
rect 159018 399978 159638 400046
rect 159018 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 159638 399978
rect 159018 382350 159638 399922
rect 159018 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 159638 382350
rect 159018 382226 159638 382294
rect 159018 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 159638 382226
rect 159018 382102 159638 382170
rect 159018 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 159638 382102
rect 159018 381978 159638 382046
rect 159018 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 159638 381978
rect 159018 364416 159638 381922
rect 159018 364360 159114 364416
rect 159170 364360 159238 364416
rect 159294 364360 159362 364416
rect 159418 364360 159486 364416
rect 159542 364360 159638 364416
rect 159018 364292 159638 364360
rect 159018 364236 159114 364292
rect 159170 364236 159238 364292
rect 159294 364236 159362 364292
rect 159418 364236 159486 364292
rect 159542 364236 159638 364292
rect 159018 364206 159638 364236
rect 162738 598172 163358 598268
rect 162738 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 163358 598172
rect 162738 598048 163358 598116
rect 162738 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 163358 598048
rect 162738 597924 163358 597992
rect 162738 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 163358 597924
rect 162738 597800 163358 597868
rect 162738 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 163358 597800
rect 162738 586350 163358 597744
rect 162738 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 163358 586350
rect 162738 586226 163358 586294
rect 162738 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 163358 586226
rect 162738 586102 163358 586170
rect 162738 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 163358 586102
rect 162738 585978 163358 586046
rect 162738 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 163358 585978
rect 162738 568350 163358 585922
rect 189738 597212 190358 598268
rect 189738 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 190358 597212
rect 189738 597088 190358 597156
rect 189738 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 190358 597088
rect 189738 596964 190358 597032
rect 189738 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 190358 596964
rect 189738 596840 190358 596908
rect 189738 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 190358 596840
rect 189738 580350 190358 596784
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 189738 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 190358 580350
rect 189738 580226 190358 580294
rect 189738 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 190358 580226
rect 189738 580102 190358 580170
rect 189738 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 190358 580102
rect 189738 579978 190358 580046
rect 189738 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 190358 579978
rect 162738 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 163358 568350
rect 162738 568226 163358 568294
rect 162738 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 163358 568226
rect 162738 568102 163358 568170
rect 162738 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 163358 568102
rect 162738 567978 163358 568046
rect 162738 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 163358 567978
rect 162738 550350 163358 567922
rect 162738 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 163358 550350
rect 162738 550226 163358 550294
rect 162738 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 163358 550226
rect 162738 550102 163358 550170
rect 162738 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 163358 550102
rect 162738 549978 163358 550046
rect 162738 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 163358 549978
rect 162738 532350 163358 549922
rect 162738 532294 162834 532350
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 163358 532350
rect 162738 532226 163358 532294
rect 162738 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 163358 532226
rect 162738 532102 163358 532170
rect 162738 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 163358 532102
rect 162738 531978 163358 532046
rect 162738 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 163358 531978
rect 162738 514350 163358 531922
rect 162738 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 163358 514350
rect 162738 514226 163358 514294
rect 162738 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 163358 514226
rect 162738 514102 163358 514170
rect 162738 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 163358 514102
rect 162738 513978 163358 514046
rect 162738 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 163358 513978
rect 162738 496350 163358 513922
rect 162738 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 163358 496350
rect 162738 496226 163358 496294
rect 162738 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 163358 496226
rect 162738 496102 163358 496170
rect 162738 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 163358 496102
rect 162738 495978 163358 496046
rect 162738 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 163358 495978
rect 162738 478350 163358 495922
rect 162738 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 163358 478350
rect 162738 478226 163358 478294
rect 162738 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 163358 478226
rect 162738 478102 163358 478170
rect 162738 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 163358 478102
rect 162738 477978 163358 478046
rect 162738 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 163358 477978
rect 162738 460350 163358 477922
rect 183036 575540 183092 575550
rect 177212 469588 177268 469598
rect 162738 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 163358 460350
rect 162738 460226 163358 460294
rect 162738 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 163358 460226
rect 162738 460102 163358 460170
rect 162738 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 163358 460102
rect 162738 459978 163358 460046
rect 162738 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 163358 459978
rect 162738 442350 163358 459922
rect 162738 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 163358 442350
rect 162738 442226 163358 442294
rect 162738 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 163358 442226
rect 162738 442102 163358 442170
rect 162738 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 163358 442102
rect 162738 441978 163358 442046
rect 162738 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 163358 441978
rect 162738 424350 163358 441922
rect 162738 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 163358 424350
rect 162738 424226 163358 424294
rect 162738 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 163358 424226
rect 162738 424102 163358 424170
rect 162738 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 163358 424102
rect 162738 423978 163358 424046
rect 162738 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 163358 423978
rect 162738 406350 163358 423922
rect 162738 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 163358 406350
rect 162738 406226 163358 406294
rect 162738 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 163358 406226
rect 162738 406102 163358 406170
rect 162738 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 163358 406102
rect 162738 405978 163358 406046
rect 162738 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 163358 405978
rect 162738 388350 163358 405922
rect 162738 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 163358 388350
rect 162738 388226 163358 388294
rect 162738 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 163358 388226
rect 162738 388102 163358 388170
rect 162738 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 163358 388102
rect 162738 387978 163358 388046
rect 162738 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 163358 387978
rect 162738 370350 163358 387922
rect 162738 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 163358 370350
rect 162738 370226 163358 370294
rect 162738 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 163358 370226
rect 162738 370102 163358 370170
rect 162738 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 163358 370102
rect 162738 369978 163358 370046
rect 162738 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 163358 369978
rect 162738 364206 163358 369922
rect 175532 466228 175588 466238
rect 132018 352294 132114 352350
rect 132170 352294 132238 352350
rect 132294 352294 132362 352350
rect 132418 352294 132486 352350
rect 132542 352294 132638 352350
rect 132018 352226 132638 352294
rect 132018 352170 132114 352226
rect 132170 352170 132238 352226
rect 132294 352170 132362 352226
rect 132418 352170 132486 352226
rect 132542 352170 132638 352226
rect 132018 352102 132638 352170
rect 132018 352046 132114 352102
rect 132170 352046 132238 352102
rect 132294 352046 132362 352102
rect 132418 352046 132486 352102
rect 132542 352046 132638 352102
rect 132018 351978 132638 352046
rect 132018 351922 132114 351978
rect 132170 351922 132238 351978
rect 132294 351922 132362 351978
rect 132418 351922 132486 351978
rect 132542 351922 132638 351978
rect 132018 334350 132638 351922
rect 149808 352350 150128 352384
rect 149808 352294 149878 352350
rect 149934 352294 150002 352350
rect 150058 352294 150128 352350
rect 149808 352226 150128 352294
rect 149808 352170 149878 352226
rect 149934 352170 150002 352226
rect 150058 352170 150128 352226
rect 149808 352102 150128 352170
rect 149808 352046 149878 352102
rect 149934 352046 150002 352102
rect 150058 352046 150128 352102
rect 149808 351978 150128 352046
rect 149808 351922 149878 351978
rect 149934 351922 150002 351978
rect 150058 351922 150128 351978
rect 149808 351888 150128 351922
rect 134448 346350 134768 346384
rect 134448 346294 134518 346350
rect 134574 346294 134642 346350
rect 134698 346294 134768 346350
rect 134448 346226 134768 346294
rect 134448 346170 134518 346226
rect 134574 346170 134642 346226
rect 134698 346170 134768 346226
rect 134448 346102 134768 346170
rect 134448 346046 134518 346102
rect 134574 346046 134642 346102
rect 134698 346046 134768 346102
rect 134448 345978 134768 346046
rect 134448 345922 134518 345978
rect 134574 345922 134642 345978
rect 134698 345922 134768 345978
rect 134448 345888 134768 345922
rect 165168 346350 165488 346384
rect 165168 346294 165238 346350
rect 165294 346294 165362 346350
rect 165418 346294 165488 346350
rect 165168 346226 165488 346294
rect 165168 346170 165238 346226
rect 165294 346170 165362 346226
rect 165418 346170 165488 346226
rect 165168 346102 165488 346170
rect 165168 346046 165238 346102
rect 165294 346046 165362 346102
rect 165418 346046 165488 346102
rect 165168 345978 165488 346046
rect 165168 345922 165238 345978
rect 165294 345922 165362 345978
rect 165418 345922 165488 345978
rect 165168 345888 165488 345922
rect 132018 334294 132114 334350
rect 132170 334294 132238 334350
rect 132294 334294 132362 334350
rect 132418 334294 132486 334350
rect 132542 334294 132638 334350
rect 132018 334226 132638 334294
rect 132018 334170 132114 334226
rect 132170 334170 132238 334226
rect 132294 334170 132362 334226
rect 132418 334170 132486 334226
rect 132542 334170 132638 334226
rect 132018 334102 132638 334170
rect 132018 334046 132114 334102
rect 132170 334046 132238 334102
rect 132294 334046 132362 334102
rect 132418 334046 132486 334102
rect 132542 334046 132638 334102
rect 132018 333978 132638 334046
rect 132018 333922 132114 333978
rect 132170 333922 132238 333978
rect 132294 333922 132362 333978
rect 132418 333922 132486 333978
rect 132542 333922 132638 333978
rect 132018 316350 132638 333922
rect 149808 334350 150128 334384
rect 149808 334294 149878 334350
rect 149934 334294 150002 334350
rect 150058 334294 150128 334350
rect 149808 334226 150128 334294
rect 149808 334170 149878 334226
rect 149934 334170 150002 334226
rect 150058 334170 150128 334226
rect 149808 334102 150128 334170
rect 149808 334046 149878 334102
rect 149934 334046 150002 334102
rect 150058 334046 150128 334102
rect 149808 333978 150128 334046
rect 149808 333922 149878 333978
rect 149934 333922 150002 333978
rect 150058 333922 150128 333978
rect 149808 333888 150128 333922
rect 134448 328350 134768 328384
rect 134448 328294 134518 328350
rect 134574 328294 134642 328350
rect 134698 328294 134768 328350
rect 134448 328226 134768 328294
rect 134448 328170 134518 328226
rect 134574 328170 134642 328226
rect 134698 328170 134768 328226
rect 134448 328102 134768 328170
rect 134448 328046 134518 328102
rect 134574 328046 134642 328102
rect 134698 328046 134768 328102
rect 134448 327978 134768 328046
rect 134448 327922 134518 327978
rect 134574 327922 134642 327978
rect 134698 327922 134768 327978
rect 134448 327888 134768 327922
rect 165168 328350 165488 328384
rect 165168 328294 165238 328350
rect 165294 328294 165362 328350
rect 165418 328294 165488 328350
rect 165168 328226 165488 328294
rect 165168 328170 165238 328226
rect 165294 328170 165362 328226
rect 165418 328170 165488 328226
rect 165168 328102 165488 328170
rect 165168 328046 165238 328102
rect 165294 328046 165362 328102
rect 165418 328046 165488 328102
rect 165168 327978 165488 328046
rect 165168 327922 165238 327978
rect 165294 327922 165362 327978
rect 165418 327922 165488 327978
rect 165168 327888 165488 327922
rect 132018 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 132638 316350
rect 132018 316226 132638 316294
rect 132018 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 132638 316226
rect 132018 316102 132638 316170
rect 132018 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 132638 316102
rect 132018 315978 132638 316046
rect 132018 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 132638 315978
rect 132018 298350 132638 315922
rect 132018 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 132638 298350
rect 132018 298226 132638 298294
rect 132018 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 132638 298226
rect 132018 298102 132638 298170
rect 132018 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 132638 298102
rect 132018 297978 132638 298046
rect 132018 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 132638 297978
rect 132018 280350 132638 297922
rect 159018 310350 159638 323954
rect 159018 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 159638 310350
rect 159018 310226 159638 310294
rect 159018 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 159638 310226
rect 159018 310102 159638 310170
rect 159018 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 159638 310102
rect 159018 309978 159638 310046
rect 159018 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 159638 309978
rect 159018 292350 159638 309922
rect 159018 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 159638 292350
rect 159018 292226 159638 292294
rect 159018 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 159638 292226
rect 159018 292102 159638 292170
rect 159018 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 159638 292102
rect 159018 291978 159638 292046
rect 159018 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 159638 291978
rect 132018 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 132638 280350
rect 132018 280226 132638 280294
rect 132018 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 132638 280226
rect 132018 280102 132638 280170
rect 132018 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 132638 280102
rect 132018 279978 132638 280046
rect 132018 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 132638 279978
rect 132018 262350 132638 279922
rect 132018 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 132638 262350
rect 132018 262226 132638 262294
rect 132018 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 132638 262226
rect 132018 262102 132638 262170
rect 132018 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 132638 262102
rect 132018 261978 132638 262046
rect 132018 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 132638 261978
rect 132018 244350 132638 261922
rect 132018 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 132638 244350
rect 132018 244226 132638 244294
rect 132018 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 132638 244226
rect 132018 244102 132638 244170
rect 132018 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 132638 244102
rect 132018 243978 132638 244046
rect 132018 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 132638 243978
rect 132018 226350 132638 243922
rect 132018 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 132638 226350
rect 132018 226226 132638 226294
rect 132018 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 132638 226226
rect 132018 226102 132638 226170
rect 132018 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 132638 226102
rect 132018 225978 132638 226046
rect 132018 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 132638 225978
rect 132018 210462 132638 225922
rect 138572 290500 138628 290510
rect 138572 217700 138628 290444
rect 159018 284908 159638 291922
rect 162738 316350 163358 323954
rect 175308 322756 175364 322766
rect 162738 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 163358 316350
rect 162738 316226 163358 316294
rect 162738 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 163358 316226
rect 162738 316102 163358 316170
rect 162738 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 163358 316102
rect 162738 315978 163358 316046
rect 162738 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 163358 315978
rect 162738 298350 163358 315922
rect 172172 322678 172228 322688
rect 168812 306628 168868 306638
rect 162738 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 163358 298350
rect 162738 298226 163358 298294
rect 162738 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 163358 298226
rect 162738 298102 163358 298170
rect 162738 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 163358 298102
rect 162738 297978 163358 298046
rect 162738 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 163358 297978
rect 162738 282254 163358 297922
rect 167244 304948 167300 304958
rect 165452 296100 165508 296110
rect 147008 280350 147328 280384
rect 147008 280294 147078 280350
rect 147134 280294 147202 280350
rect 147258 280294 147328 280350
rect 147008 280226 147328 280294
rect 147008 280170 147078 280226
rect 147134 280170 147202 280226
rect 147258 280170 147328 280226
rect 147008 280102 147328 280170
rect 147008 280046 147078 280102
rect 147134 280046 147202 280102
rect 147258 280046 147328 280102
rect 147008 279978 147328 280046
rect 147008 279922 147078 279978
rect 147134 279922 147202 279978
rect 147258 279922 147328 279978
rect 147008 279888 147328 279922
rect 152832 280350 153152 280384
rect 152832 280294 152902 280350
rect 152958 280294 153026 280350
rect 153082 280294 153152 280350
rect 152832 280226 153152 280294
rect 152832 280170 152902 280226
rect 152958 280170 153026 280226
rect 153082 280170 153152 280226
rect 152832 280102 153152 280170
rect 152832 280046 152902 280102
rect 152958 280046 153026 280102
rect 153082 280046 153152 280102
rect 152832 279978 153152 280046
rect 152832 279922 152902 279978
rect 152958 279922 153026 279978
rect 153082 279922 153152 279978
rect 152832 279888 153152 279922
rect 158656 280350 158976 280384
rect 158656 280294 158726 280350
rect 158782 280294 158850 280350
rect 158906 280294 158976 280350
rect 158656 280226 158976 280294
rect 158656 280170 158726 280226
rect 158782 280170 158850 280226
rect 158906 280170 158976 280226
rect 158656 280102 158976 280170
rect 158656 280046 158726 280102
rect 158782 280046 158850 280102
rect 158906 280046 158976 280102
rect 158656 279978 158976 280046
rect 158656 279922 158726 279978
rect 158782 279922 158850 279978
rect 158906 279922 158976 279978
rect 158656 279888 158976 279922
rect 164480 280350 164800 280384
rect 164480 280294 164550 280350
rect 164606 280294 164674 280350
rect 164730 280294 164800 280350
rect 164480 280226 164800 280294
rect 164480 280170 164550 280226
rect 164606 280170 164674 280226
rect 164730 280170 164800 280226
rect 164480 280102 164800 280170
rect 164480 280046 164550 280102
rect 164606 280046 164674 280102
rect 164730 280046 164800 280102
rect 164480 279978 164800 280046
rect 164480 279922 164550 279978
rect 164606 279922 164674 279978
rect 164730 279922 164800 279978
rect 164480 279888 164800 279922
rect 165452 279300 165508 296044
rect 165452 279234 165508 279244
rect 165676 290276 165732 290286
rect 165676 277284 165732 290220
rect 165676 277218 165732 277228
rect 167132 289156 167188 289166
rect 144096 274350 144416 274384
rect 144096 274294 144166 274350
rect 144222 274294 144290 274350
rect 144346 274294 144416 274350
rect 144096 274226 144416 274294
rect 144096 274170 144166 274226
rect 144222 274170 144290 274226
rect 144346 274170 144416 274226
rect 144096 274102 144416 274170
rect 144096 274046 144166 274102
rect 144222 274046 144290 274102
rect 144346 274046 144416 274102
rect 144096 273978 144416 274046
rect 144096 273922 144166 273978
rect 144222 273922 144290 273978
rect 144346 273922 144416 273978
rect 144096 273888 144416 273922
rect 149920 274350 150240 274384
rect 149920 274294 149990 274350
rect 150046 274294 150114 274350
rect 150170 274294 150240 274350
rect 149920 274226 150240 274294
rect 149920 274170 149990 274226
rect 150046 274170 150114 274226
rect 150170 274170 150240 274226
rect 149920 274102 150240 274170
rect 149920 274046 149990 274102
rect 150046 274046 150114 274102
rect 150170 274046 150240 274102
rect 149920 273978 150240 274046
rect 149920 273922 149990 273978
rect 150046 273922 150114 273978
rect 150170 273922 150240 273978
rect 149920 273888 150240 273922
rect 155744 274350 156064 274384
rect 155744 274294 155814 274350
rect 155870 274294 155938 274350
rect 155994 274294 156064 274350
rect 155744 274226 156064 274294
rect 155744 274170 155814 274226
rect 155870 274170 155938 274226
rect 155994 274170 156064 274226
rect 155744 274102 156064 274170
rect 155744 274046 155814 274102
rect 155870 274046 155938 274102
rect 155994 274046 156064 274102
rect 155744 273978 156064 274046
rect 155744 273922 155814 273978
rect 155870 273922 155938 273978
rect 155994 273922 156064 273978
rect 155744 273888 156064 273922
rect 161568 274350 161888 274384
rect 161568 274294 161638 274350
rect 161694 274294 161762 274350
rect 161818 274294 161888 274350
rect 161568 274226 161888 274294
rect 161568 274170 161638 274226
rect 161694 274170 161762 274226
rect 161818 274170 161888 274226
rect 161568 274102 161888 274170
rect 161568 274046 161638 274102
rect 161694 274046 161762 274102
rect 161818 274046 161888 274102
rect 161568 273978 161888 274046
rect 161568 273922 161638 273978
rect 161694 273922 161762 273978
rect 161818 273922 161888 273978
rect 161568 273888 161888 273922
rect 162738 262350 163358 265522
rect 162738 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 163358 262350
rect 162738 262226 163358 262294
rect 162738 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 163358 262226
rect 162738 262102 163358 262170
rect 162738 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 163358 262102
rect 162738 261978 163358 262046
rect 162738 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 163358 261978
rect 138572 217634 138628 217644
rect 159018 256350 159638 260964
rect 159018 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 159638 256350
rect 159018 256226 159638 256294
rect 159018 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 159638 256226
rect 159018 256102 159638 256170
rect 159018 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 159638 256102
rect 159018 255978 159638 256046
rect 159018 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 159638 255978
rect 159018 238350 159638 255922
rect 159018 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 159638 238350
rect 159018 238226 159638 238294
rect 159018 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 159638 238226
rect 159018 238102 159638 238170
rect 159018 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 159638 238102
rect 159018 237978 159638 238046
rect 159018 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 159638 237978
rect 159018 220350 159638 237922
rect 159018 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 159638 220350
rect 159018 220226 159638 220294
rect 159018 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 159638 220226
rect 159018 220102 159638 220170
rect 159018 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 159638 220102
rect 159018 219978 159638 220046
rect 159018 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 159638 219978
rect 159018 210462 159638 219922
rect 162738 244350 163358 261922
rect 162738 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 163358 244350
rect 162738 244226 163358 244294
rect 162738 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 163358 244226
rect 162738 244102 163358 244170
rect 162738 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 163358 244102
rect 162738 243978 163358 244046
rect 162738 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 163358 243978
rect 162738 226350 163358 243922
rect 162738 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 163358 226350
rect 162738 226226 163358 226294
rect 162738 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 163358 226226
rect 162738 226102 163358 226170
rect 162738 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 163358 226102
rect 162738 225978 163358 226046
rect 162738 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 163358 225978
rect 162738 210462 163358 225922
rect 167132 212660 167188 289100
rect 167244 282436 167300 304892
rect 167244 282370 167300 282380
rect 168812 281092 168868 306572
rect 168812 281026 168868 281036
rect 170492 281458 170548 281468
rect 168140 279300 168196 279310
rect 168140 278964 168196 279244
rect 168028 278068 168084 278078
rect 168028 277284 168084 278012
rect 168028 261828 168084 277228
rect 168140 263844 168196 278908
rect 170492 269892 170548 281402
rect 170492 269826 170548 269836
rect 168140 263778 168196 263788
rect 168028 261762 168084 261772
rect 172172 217700 172228 322622
rect 175308 321860 175364 322700
rect 175308 321794 175364 321804
rect 174524 321412 174580 321422
rect 174412 318724 174468 318734
rect 174300 312004 174356 312014
rect 172284 296660 172340 296670
rect 172284 283780 172340 296604
rect 172284 283714 172340 283724
rect 172172 217634 172228 217644
rect 167132 212594 167188 212604
rect 174300 210532 174356 311948
rect 174412 212772 174468 318668
rect 174524 212884 174580 321356
rect 174524 212818 174580 212828
rect 174636 320068 174692 320078
rect 174412 212706 174468 212716
rect 174300 210466 174356 210476
rect 174636 209636 174692 320012
rect 175532 277060 175588 466172
rect 175532 276994 175588 277004
rect 175644 281428 175700 281438
rect 175644 268772 175700 281372
rect 177212 274372 177268 469532
rect 180572 467908 180628 467918
rect 177324 431956 177380 431966
rect 177324 278404 177380 431900
rect 178892 358708 178948 358718
rect 178108 340138 178164 340148
rect 178108 339556 178164 340082
rect 178108 320180 178164 339500
rect 178892 326116 178948 358652
rect 178892 326050 178948 326060
rect 178108 320114 178164 320124
rect 177324 278338 177380 278348
rect 177884 317380 177940 317390
rect 177212 274306 177268 274316
rect 175644 268706 175700 268716
rect 177884 219716 177940 317324
rect 179676 316036 179732 316046
rect 177884 219650 177940 219660
rect 177996 313348 178052 313358
rect 177996 211092 178052 313292
rect 179676 212996 179732 315980
rect 180572 275716 180628 467852
rect 182476 377860 182532 377870
rect 182252 377188 182308 377198
rect 180684 373828 180740 373838
rect 180684 352996 180740 373772
rect 180684 352930 180740 352940
rect 181356 325444 181412 325454
rect 180572 275650 180628 275660
rect 181244 306628 181300 306638
rect 181244 219828 181300 306572
rect 181244 219762 181300 219772
rect 179676 212930 179732 212940
rect 177996 211026 178052 211036
rect 174636 209570 174692 209580
rect 181356 209412 181412 325388
rect 182252 279748 182308 377132
rect 182476 363076 182532 377804
rect 182476 363010 182532 363020
rect 182924 299908 182980 299918
rect 182252 279682 182308 279692
rect 182364 285684 182420 285694
rect 182364 281988 182420 285628
rect 182364 239876 182420 281932
rect 182476 283668 182532 283678
rect 182476 272132 182532 283612
rect 182476 272066 182532 272076
rect 182364 239810 182420 239820
rect 182924 214788 182980 299852
rect 183036 260932 183092 575484
rect 184716 567924 184772 567934
rect 184492 522116 184548 522126
rect 183932 500612 183988 500622
rect 183932 285684 183988 500556
rect 184492 378838 184548 522060
rect 184492 378772 184548 378782
rect 184604 401604 184660 401614
rect 184156 375172 184212 375182
rect 184044 372484 184100 372494
rect 184044 350420 184100 372428
rect 184156 356356 184212 375116
rect 184156 356290 184212 356300
rect 184044 350354 184100 350364
rect 183932 285618 183988 285628
rect 184380 314692 184436 314702
rect 183036 260866 183092 260876
rect 184380 239316 184436 314636
rect 184380 239250 184436 239260
rect 184492 305284 184548 305294
rect 182924 214722 182980 214732
rect 184492 213220 184548 305228
rect 184604 254212 184660 401548
rect 184716 259588 184772 567868
rect 189738 562350 190358 579922
rect 189738 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 190358 562350
rect 189738 562226 190358 562294
rect 189738 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 190358 562226
rect 189738 562102 190358 562170
rect 189738 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 190358 562102
rect 189738 561978 190358 562046
rect 189738 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 190358 561978
rect 189738 544350 190358 561922
rect 189738 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 190358 544350
rect 189738 544226 190358 544294
rect 189738 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 190358 544226
rect 189738 544102 190358 544170
rect 189738 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 190358 544102
rect 189738 543978 190358 544046
rect 189738 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 190358 543978
rect 186396 529284 186452 529294
rect 185388 428932 185444 428942
rect 185388 278068 185444 428876
rect 186172 404038 186228 404048
rect 185948 402418 186004 402428
rect 185612 371140 185668 371150
rect 185388 277284 185444 278012
rect 185388 277218 185444 277228
rect 185500 364420 185556 364430
rect 184716 259522 184772 259532
rect 184604 254146 184660 254156
rect 184492 213154 184548 213164
rect 185500 211078 185556 364364
rect 185612 358708 185668 371084
rect 185612 358642 185668 358652
rect 185836 310660 185892 310670
rect 185724 307972 185780 307982
rect 185724 211204 185780 307916
rect 185724 211138 185780 211148
rect 185500 211012 185556 211022
rect 185836 209748 185892 310604
rect 185948 256900 186004 402362
rect 185948 256834 186004 256844
rect 186060 402388 186116 402398
rect 186060 255556 186116 402332
rect 186172 258244 186228 403982
rect 186396 383908 186452 529228
rect 189738 526350 190358 543922
rect 189738 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 190358 526350
rect 189738 526226 190358 526294
rect 189738 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 190358 526226
rect 189738 526102 190358 526170
rect 189738 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 190358 526102
rect 189738 525978 190358 526046
rect 189738 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 190358 525978
rect 189738 508350 190358 525922
rect 189738 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 190358 508350
rect 189738 508226 190358 508294
rect 189738 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 190358 508226
rect 189738 508102 190358 508170
rect 189738 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 190358 508102
rect 189738 507978 190358 508046
rect 189738 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 190358 507978
rect 189738 490350 190358 507922
rect 189738 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 190358 490350
rect 189738 490226 190358 490294
rect 189738 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 190358 490226
rect 189738 490102 190358 490170
rect 189738 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 190358 490102
rect 189738 489978 190358 490046
rect 189738 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 190358 489978
rect 187516 486276 187572 486286
rect 186396 383842 186452 383852
rect 187292 436100 187348 436110
rect 186956 302596 187012 302606
rect 186844 301252 186900 301262
rect 186508 282212 186564 282222
rect 186172 258178 186228 258188
rect 186284 280420 186340 280430
rect 186284 279076 186340 280364
rect 186060 255490 186116 255500
rect 186284 239764 186340 279020
rect 186508 278908 186564 282156
rect 186396 278852 186564 278908
rect 186396 268858 186452 278852
rect 186396 265860 186452 268802
rect 186396 265794 186452 265804
rect 186284 239698 186340 239708
rect 186844 218148 186900 301196
rect 186844 218082 186900 218092
rect 186956 218036 187012 302540
rect 187068 298564 187124 298574
rect 187068 241332 187124 298508
rect 187292 290668 187348 436044
rect 187404 376516 187460 376526
rect 187404 359716 187460 376460
rect 187404 359650 187460 359660
rect 187404 322756 187460 322766
rect 187404 322678 187460 322700
rect 187404 322612 187460 322622
rect 187516 296548 187572 486220
rect 187964 479108 188020 479118
rect 187852 457604 187908 457614
rect 187740 303940 187796 303950
rect 187516 296482 187572 296492
rect 187628 297220 187684 297230
rect 187180 290612 187348 290668
rect 187404 295876 187460 295886
rect 187180 287398 187236 290612
rect 187292 289828 187348 289838
rect 187292 289018 187348 289772
rect 187292 288952 187348 288962
rect 187180 287342 187348 287398
rect 187180 287218 187236 287228
rect 187180 285684 187236 287162
rect 187180 285618 187236 285628
rect 187180 280532 187236 280542
rect 187180 252868 187236 280476
rect 187292 280420 187348 287342
rect 187292 280354 187348 280364
rect 187180 252802 187236 252812
rect 187292 277284 187348 277294
rect 187068 241266 187124 241276
rect 187292 239652 187348 277228
rect 187404 241220 187460 295820
rect 187404 241154 187460 241164
rect 187516 294532 187572 294542
rect 187292 239586 187348 239596
rect 186956 217970 187012 217980
rect 187516 216468 187572 294476
rect 187628 216580 187684 297164
rect 187740 221172 187796 303884
rect 187852 281458 187908 457548
rect 187964 295652 188020 479052
rect 187964 295586 188020 295596
rect 189738 472350 190358 489922
rect 189738 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 190358 472350
rect 189738 472226 190358 472294
rect 189738 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 190358 472226
rect 189738 472102 190358 472170
rect 189738 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 190358 472102
rect 189738 471978 190358 472046
rect 189738 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 190358 471978
rect 189738 454350 190358 471922
rect 189738 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 190358 454350
rect 189738 454226 190358 454294
rect 189738 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 190358 454226
rect 189738 454102 190358 454170
rect 189738 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 190358 454102
rect 189738 453978 190358 454046
rect 189738 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 190358 453978
rect 189738 436350 190358 453922
rect 189738 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 190358 436350
rect 189738 436226 190358 436294
rect 189738 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 190358 436226
rect 189738 436102 190358 436170
rect 189738 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 190358 436102
rect 189738 435978 190358 436046
rect 189738 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 190358 435978
rect 189738 418350 190358 435922
rect 193116 591108 193172 591118
rect 190652 421876 190708 421896
rect 190652 421792 190708 421802
rect 192332 421858 192388 421868
rect 189738 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 190358 418350
rect 189738 418226 190358 418294
rect 189738 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 190358 418226
rect 189738 418102 190358 418170
rect 189738 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 190358 418102
rect 189738 417978 190358 418046
rect 189738 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 190358 417978
rect 189738 400350 190358 417922
rect 189738 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 190358 400350
rect 189738 400226 190358 400294
rect 189738 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 190358 400226
rect 189738 400102 190358 400170
rect 189738 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 190358 400102
rect 189738 399978 190358 400046
rect 189738 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 190358 399978
rect 189738 382350 190358 399922
rect 189738 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 190358 382350
rect 189738 382226 190358 382294
rect 189738 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 190358 382226
rect 189738 382102 190358 382170
rect 189738 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 190358 382102
rect 189738 381978 190358 382046
rect 189738 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 190358 381978
rect 189738 364350 190358 381922
rect 192332 379204 192388 421802
rect 193116 407764 193172 591052
rect 193340 590884 193396 590894
rect 193340 409108 193396 590828
rect 193458 586350 194078 597744
rect 220458 597212 221078 598268
rect 220458 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 221078 597212
rect 220458 597088 221078 597156
rect 220458 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 221078 597088
rect 220458 596964 221078 597032
rect 220458 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 221078 596964
rect 220458 596840 221078 596908
rect 220458 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 221078 596840
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 193458 568670 194078 585922
rect 194236 590660 194292 590670
rect 193340 409042 193396 409052
rect 193116 407698 193172 407708
rect 192332 379138 192388 379148
rect 193458 406350 194078 410034
rect 193458 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 194078 406350
rect 193458 406226 194078 406294
rect 193458 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 194078 406226
rect 193458 406102 194078 406170
rect 193458 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 194078 406102
rect 193458 405978 194078 406046
rect 193458 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 194078 405978
rect 193458 388350 194078 405922
rect 194236 405860 194292 590604
rect 220458 580350 221078 596784
rect 220458 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 221078 580350
rect 220458 580226 221078 580294
rect 220458 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 221078 580226
rect 220458 580102 221078 580170
rect 220458 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 221078 580102
rect 220458 579978 221078 580046
rect 220458 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 221078 579978
rect 220458 568670 221078 579922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 568670 224798 585922
rect 251178 597212 251798 598268
rect 251178 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 251798 597212
rect 251178 597088 251798 597156
rect 251178 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 251798 597088
rect 251178 596964 251798 597032
rect 251178 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 251798 596964
rect 251178 596840 251798 596908
rect 251178 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 251798 596840
rect 251178 580350 251798 596784
rect 251178 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 251798 580350
rect 251178 580226 251798 580294
rect 251178 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 251798 580226
rect 251178 580102 251798 580170
rect 251178 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 251798 580102
rect 251178 579978 251798 580046
rect 251178 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 251798 579978
rect 251178 568670 251798 579922
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 568670 255518 585922
rect 281898 597212 282518 598268
rect 281898 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 282518 597212
rect 281898 597088 282518 597156
rect 281898 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 282518 597088
rect 281898 596964 282518 597032
rect 281898 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 282518 596964
rect 281898 596840 282518 596908
rect 281898 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 282518 596840
rect 281898 580350 282518 596784
rect 281898 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 282518 580350
rect 281898 580226 282518 580294
rect 281898 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 282518 580226
rect 281898 580102 282518 580170
rect 281898 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 282518 580102
rect 281898 579978 282518 580046
rect 281898 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 282518 579978
rect 281898 568670 282518 579922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 568670 286238 585922
rect 312618 597212 313238 598268
rect 312618 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 313238 597212
rect 312618 597088 313238 597156
rect 312618 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 313238 597088
rect 312618 596964 313238 597032
rect 312618 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 313238 596964
rect 312618 596840 313238 596908
rect 312618 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 313238 596840
rect 312618 580350 313238 596784
rect 312618 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 313238 580350
rect 312618 580226 313238 580294
rect 312618 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 313238 580226
rect 312618 580102 313238 580170
rect 312618 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 313238 580102
rect 312618 579978 313238 580046
rect 312618 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 313238 579978
rect 312618 568670 313238 579922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 316338 568670 316958 585922
rect 343338 597212 343958 598268
rect 343338 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 343958 597212
rect 343338 597088 343958 597156
rect 343338 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 343958 597088
rect 343338 596964 343958 597032
rect 343338 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 343958 596964
rect 343338 596840 343958 596908
rect 343338 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 343958 596840
rect 343338 580350 343958 596784
rect 343338 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 343958 580350
rect 343338 580226 343958 580294
rect 343338 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 343958 580226
rect 343338 580102 343958 580170
rect 343338 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 343958 580102
rect 343338 579978 343958 580046
rect 343338 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 343958 579978
rect 343338 568670 343958 579922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 568670 347678 585922
rect 374058 597212 374678 598268
rect 374058 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 374678 597212
rect 374058 597088 374678 597156
rect 374058 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 374678 597088
rect 374058 596964 374678 597032
rect 374058 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 374678 596964
rect 374058 596840 374678 596908
rect 374058 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 374678 596840
rect 374058 580350 374678 596784
rect 374058 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 374678 580350
rect 374058 580226 374678 580294
rect 374058 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 374678 580226
rect 374058 580102 374678 580170
rect 374058 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 374678 580102
rect 374058 579978 374678 580046
rect 374058 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 374678 579978
rect 374058 568670 374678 579922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 568670 378398 585922
rect 404778 597212 405398 598268
rect 404778 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 405398 597212
rect 404778 597088 405398 597156
rect 404778 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 405398 597088
rect 404778 596964 405398 597032
rect 404778 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 405398 596964
rect 404778 596840 405398 596908
rect 404778 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 405398 596840
rect 404778 580350 405398 596784
rect 404778 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 405398 580350
rect 404778 580226 405398 580294
rect 404778 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 405398 580226
rect 404778 580102 405398 580170
rect 404778 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 405398 580102
rect 404778 579978 405398 580046
rect 404778 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 405398 579978
rect 404778 568670 405398 579922
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 568670 409118 585922
rect 435498 597212 436118 598268
rect 435498 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 436118 597212
rect 435498 597088 436118 597156
rect 435498 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 436118 597088
rect 435498 596964 436118 597032
rect 435498 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 436118 596964
rect 435498 596840 436118 596908
rect 435498 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 436118 596840
rect 435498 580350 436118 596784
rect 435498 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 436118 580350
rect 435498 580226 436118 580294
rect 435498 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 436118 580226
rect 435498 580102 436118 580170
rect 435498 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 436118 580102
rect 435498 579978 436118 580046
rect 435498 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 436118 579978
rect 435498 568670 436118 579922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 568670 439838 585922
rect 466218 597212 466838 598268
rect 466218 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 466838 597212
rect 466218 597088 466838 597156
rect 466218 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 466838 597088
rect 466218 596964 466838 597032
rect 466218 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 466838 596964
rect 466218 596840 466838 596908
rect 466218 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 466838 596840
rect 466218 580350 466838 596784
rect 466218 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 466838 580350
rect 466218 580226 466838 580294
rect 466218 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 466838 580226
rect 466218 580102 466838 580170
rect 466218 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 466838 580102
rect 466218 579978 466838 580046
rect 466218 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 466838 579978
rect 466218 568670 466838 579922
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 568670 470558 585922
rect 496938 597212 497558 598268
rect 496938 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 497558 597212
rect 496938 597088 497558 597156
rect 496938 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 497558 597088
rect 496938 596964 497558 597032
rect 496938 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 497558 596964
rect 496938 596840 497558 596908
rect 496938 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 497558 596840
rect 496938 580350 497558 596784
rect 496938 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 497558 580350
rect 496938 580226 497558 580294
rect 496938 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 497558 580226
rect 496938 580102 497558 580170
rect 496938 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 497558 580102
rect 496938 579978 497558 580046
rect 496938 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 497558 579978
rect 496938 568670 497558 579922
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 527658 597212 528278 598268
rect 527658 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 528278 597212
rect 527658 597088 528278 597156
rect 527658 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 528278 597088
rect 527658 596964 528278 597032
rect 527658 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 528278 596964
rect 527658 596840 528278 596908
rect 527658 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 528278 596840
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 568670 501278 585922
rect 511308 590660 511364 590670
rect 194448 562350 194768 562384
rect 194448 562294 194518 562350
rect 194574 562294 194642 562350
rect 194698 562294 194768 562350
rect 194448 562226 194768 562294
rect 194448 562170 194518 562226
rect 194574 562170 194642 562226
rect 194698 562170 194768 562226
rect 194448 562102 194768 562170
rect 194448 562046 194518 562102
rect 194574 562046 194642 562102
rect 194698 562046 194768 562102
rect 194448 561978 194768 562046
rect 194448 561922 194518 561978
rect 194574 561922 194642 561978
rect 194698 561922 194768 561978
rect 194448 561888 194768 561922
rect 225168 562350 225488 562384
rect 225168 562294 225238 562350
rect 225294 562294 225362 562350
rect 225418 562294 225488 562350
rect 225168 562226 225488 562294
rect 225168 562170 225238 562226
rect 225294 562170 225362 562226
rect 225418 562170 225488 562226
rect 225168 562102 225488 562170
rect 225168 562046 225238 562102
rect 225294 562046 225362 562102
rect 225418 562046 225488 562102
rect 225168 561978 225488 562046
rect 225168 561922 225238 561978
rect 225294 561922 225362 561978
rect 225418 561922 225488 561978
rect 225168 561888 225488 561922
rect 255888 562350 256208 562384
rect 255888 562294 255958 562350
rect 256014 562294 256082 562350
rect 256138 562294 256208 562350
rect 255888 562226 256208 562294
rect 255888 562170 255958 562226
rect 256014 562170 256082 562226
rect 256138 562170 256208 562226
rect 255888 562102 256208 562170
rect 255888 562046 255958 562102
rect 256014 562046 256082 562102
rect 256138 562046 256208 562102
rect 255888 561978 256208 562046
rect 255888 561922 255958 561978
rect 256014 561922 256082 561978
rect 256138 561922 256208 561978
rect 255888 561888 256208 561922
rect 286608 562350 286928 562384
rect 286608 562294 286678 562350
rect 286734 562294 286802 562350
rect 286858 562294 286928 562350
rect 286608 562226 286928 562294
rect 286608 562170 286678 562226
rect 286734 562170 286802 562226
rect 286858 562170 286928 562226
rect 286608 562102 286928 562170
rect 286608 562046 286678 562102
rect 286734 562046 286802 562102
rect 286858 562046 286928 562102
rect 286608 561978 286928 562046
rect 286608 561922 286678 561978
rect 286734 561922 286802 561978
rect 286858 561922 286928 561978
rect 286608 561888 286928 561922
rect 317328 562350 317648 562384
rect 317328 562294 317398 562350
rect 317454 562294 317522 562350
rect 317578 562294 317648 562350
rect 317328 562226 317648 562294
rect 317328 562170 317398 562226
rect 317454 562170 317522 562226
rect 317578 562170 317648 562226
rect 317328 562102 317648 562170
rect 317328 562046 317398 562102
rect 317454 562046 317522 562102
rect 317578 562046 317648 562102
rect 317328 561978 317648 562046
rect 317328 561922 317398 561978
rect 317454 561922 317522 561978
rect 317578 561922 317648 561978
rect 317328 561888 317648 561922
rect 348048 562350 348368 562384
rect 348048 562294 348118 562350
rect 348174 562294 348242 562350
rect 348298 562294 348368 562350
rect 348048 562226 348368 562294
rect 348048 562170 348118 562226
rect 348174 562170 348242 562226
rect 348298 562170 348368 562226
rect 348048 562102 348368 562170
rect 348048 562046 348118 562102
rect 348174 562046 348242 562102
rect 348298 562046 348368 562102
rect 348048 561978 348368 562046
rect 348048 561922 348118 561978
rect 348174 561922 348242 561978
rect 348298 561922 348368 561978
rect 348048 561888 348368 561922
rect 378768 562350 379088 562384
rect 378768 562294 378838 562350
rect 378894 562294 378962 562350
rect 379018 562294 379088 562350
rect 378768 562226 379088 562294
rect 378768 562170 378838 562226
rect 378894 562170 378962 562226
rect 379018 562170 379088 562226
rect 378768 562102 379088 562170
rect 378768 562046 378838 562102
rect 378894 562046 378962 562102
rect 379018 562046 379088 562102
rect 378768 561978 379088 562046
rect 378768 561922 378838 561978
rect 378894 561922 378962 561978
rect 379018 561922 379088 561978
rect 378768 561888 379088 561922
rect 409488 562350 409808 562384
rect 409488 562294 409558 562350
rect 409614 562294 409682 562350
rect 409738 562294 409808 562350
rect 409488 562226 409808 562294
rect 409488 562170 409558 562226
rect 409614 562170 409682 562226
rect 409738 562170 409808 562226
rect 409488 562102 409808 562170
rect 409488 562046 409558 562102
rect 409614 562046 409682 562102
rect 409738 562046 409808 562102
rect 409488 561978 409808 562046
rect 409488 561922 409558 561978
rect 409614 561922 409682 561978
rect 409738 561922 409808 561978
rect 409488 561888 409808 561922
rect 440208 562350 440528 562384
rect 440208 562294 440278 562350
rect 440334 562294 440402 562350
rect 440458 562294 440528 562350
rect 440208 562226 440528 562294
rect 440208 562170 440278 562226
rect 440334 562170 440402 562226
rect 440458 562170 440528 562226
rect 440208 562102 440528 562170
rect 440208 562046 440278 562102
rect 440334 562046 440402 562102
rect 440458 562046 440528 562102
rect 440208 561978 440528 562046
rect 440208 561922 440278 561978
rect 440334 561922 440402 561978
rect 440458 561922 440528 561978
rect 440208 561888 440528 561922
rect 470928 562350 471248 562384
rect 470928 562294 470998 562350
rect 471054 562294 471122 562350
rect 471178 562294 471248 562350
rect 470928 562226 471248 562294
rect 470928 562170 470998 562226
rect 471054 562170 471122 562226
rect 471178 562170 471248 562226
rect 470928 562102 471248 562170
rect 470928 562046 470998 562102
rect 471054 562046 471122 562102
rect 471178 562046 471248 562102
rect 470928 561978 471248 562046
rect 470928 561922 470998 561978
rect 471054 561922 471122 561978
rect 471178 561922 471248 561978
rect 470928 561888 471248 561922
rect 501648 562350 501968 562384
rect 501648 562294 501718 562350
rect 501774 562294 501842 562350
rect 501898 562294 501968 562350
rect 501648 562226 501968 562294
rect 501648 562170 501718 562226
rect 501774 562170 501842 562226
rect 501898 562170 501968 562226
rect 501648 562102 501968 562170
rect 501648 562046 501718 562102
rect 501774 562046 501842 562102
rect 501898 562046 501968 562102
rect 501648 561978 501968 562046
rect 501648 561922 501718 561978
rect 501774 561922 501842 561978
rect 501898 561922 501968 561978
rect 501648 561888 501968 561922
rect 209808 550350 210128 550384
rect 209808 550294 209878 550350
rect 209934 550294 210002 550350
rect 210058 550294 210128 550350
rect 209808 550226 210128 550294
rect 209808 550170 209878 550226
rect 209934 550170 210002 550226
rect 210058 550170 210128 550226
rect 209808 550102 210128 550170
rect 209808 550046 209878 550102
rect 209934 550046 210002 550102
rect 210058 550046 210128 550102
rect 209808 549978 210128 550046
rect 209808 549922 209878 549978
rect 209934 549922 210002 549978
rect 210058 549922 210128 549978
rect 209808 549888 210128 549922
rect 240528 550350 240848 550384
rect 240528 550294 240598 550350
rect 240654 550294 240722 550350
rect 240778 550294 240848 550350
rect 240528 550226 240848 550294
rect 240528 550170 240598 550226
rect 240654 550170 240722 550226
rect 240778 550170 240848 550226
rect 240528 550102 240848 550170
rect 240528 550046 240598 550102
rect 240654 550046 240722 550102
rect 240778 550046 240848 550102
rect 240528 549978 240848 550046
rect 240528 549922 240598 549978
rect 240654 549922 240722 549978
rect 240778 549922 240848 549978
rect 240528 549888 240848 549922
rect 271248 550350 271568 550384
rect 271248 550294 271318 550350
rect 271374 550294 271442 550350
rect 271498 550294 271568 550350
rect 271248 550226 271568 550294
rect 271248 550170 271318 550226
rect 271374 550170 271442 550226
rect 271498 550170 271568 550226
rect 271248 550102 271568 550170
rect 271248 550046 271318 550102
rect 271374 550046 271442 550102
rect 271498 550046 271568 550102
rect 271248 549978 271568 550046
rect 271248 549922 271318 549978
rect 271374 549922 271442 549978
rect 271498 549922 271568 549978
rect 271248 549888 271568 549922
rect 301968 550350 302288 550384
rect 301968 550294 302038 550350
rect 302094 550294 302162 550350
rect 302218 550294 302288 550350
rect 301968 550226 302288 550294
rect 301968 550170 302038 550226
rect 302094 550170 302162 550226
rect 302218 550170 302288 550226
rect 301968 550102 302288 550170
rect 301968 550046 302038 550102
rect 302094 550046 302162 550102
rect 302218 550046 302288 550102
rect 301968 549978 302288 550046
rect 301968 549922 302038 549978
rect 302094 549922 302162 549978
rect 302218 549922 302288 549978
rect 301968 549888 302288 549922
rect 332688 550350 333008 550384
rect 332688 550294 332758 550350
rect 332814 550294 332882 550350
rect 332938 550294 333008 550350
rect 332688 550226 333008 550294
rect 332688 550170 332758 550226
rect 332814 550170 332882 550226
rect 332938 550170 333008 550226
rect 332688 550102 333008 550170
rect 332688 550046 332758 550102
rect 332814 550046 332882 550102
rect 332938 550046 333008 550102
rect 332688 549978 333008 550046
rect 332688 549922 332758 549978
rect 332814 549922 332882 549978
rect 332938 549922 333008 549978
rect 332688 549888 333008 549922
rect 363408 550350 363728 550384
rect 363408 550294 363478 550350
rect 363534 550294 363602 550350
rect 363658 550294 363728 550350
rect 363408 550226 363728 550294
rect 363408 550170 363478 550226
rect 363534 550170 363602 550226
rect 363658 550170 363728 550226
rect 363408 550102 363728 550170
rect 363408 550046 363478 550102
rect 363534 550046 363602 550102
rect 363658 550046 363728 550102
rect 363408 549978 363728 550046
rect 363408 549922 363478 549978
rect 363534 549922 363602 549978
rect 363658 549922 363728 549978
rect 363408 549888 363728 549922
rect 394128 550350 394448 550384
rect 394128 550294 394198 550350
rect 394254 550294 394322 550350
rect 394378 550294 394448 550350
rect 394128 550226 394448 550294
rect 394128 550170 394198 550226
rect 394254 550170 394322 550226
rect 394378 550170 394448 550226
rect 394128 550102 394448 550170
rect 394128 550046 394198 550102
rect 394254 550046 394322 550102
rect 394378 550046 394448 550102
rect 394128 549978 394448 550046
rect 394128 549922 394198 549978
rect 394254 549922 394322 549978
rect 394378 549922 394448 549978
rect 394128 549888 394448 549922
rect 424848 550350 425168 550384
rect 424848 550294 424918 550350
rect 424974 550294 425042 550350
rect 425098 550294 425168 550350
rect 424848 550226 425168 550294
rect 424848 550170 424918 550226
rect 424974 550170 425042 550226
rect 425098 550170 425168 550226
rect 424848 550102 425168 550170
rect 424848 550046 424918 550102
rect 424974 550046 425042 550102
rect 425098 550046 425168 550102
rect 424848 549978 425168 550046
rect 424848 549922 424918 549978
rect 424974 549922 425042 549978
rect 425098 549922 425168 549978
rect 424848 549888 425168 549922
rect 455568 550350 455888 550384
rect 455568 550294 455638 550350
rect 455694 550294 455762 550350
rect 455818 550294 455888 550350
rect 455568 550226 455888 550294
rect 455568 550170 455638 550226
rect 455694 550170 455762 550226
rect 455818 550170 455888 550226
rect 455568 550102 455888 550170
rect 455568 550046 455638 550102
rect 455694 550046 455762 550102
rect 455818 550046 455888 550102
rect 455568 549978 455888 550046
rect 455568 549922 455638 549978
rect 455694 549922 455762 549978
rect 455818 549922 455888 549978
rect 455568 549888 455888 549922
rect 486288 550350 486608 550384
rect 486288 550294 486358 550350
rect 486414 550294 486482 550350
rect 486538 550294 486608 550350
rect 486288 550226 486608 550294
rect 486288 550170 486358 550226
rect 486414 550170 486482 550226
rect 486538 550170 486608 550226
rect 486288 550102 486608 550170
rect 486288 550046 486358 550102
rect 486414 550046 486482 550102
rect 486538 550046 486608 550102
rect 486288 549978 486608 550046
rect 486288 549922 486358 549978
rect 486414 549922 486482 549978
rect 486538 549922 486608 549978
rect 486288 549888 486608 549922
rect 194448 544350 194768 544384
rect 194448 544294 194518 544350
rect 194574 544294 194642 544350
rect 194698 544294 194768 544350
rect 194448 544226 194768 544294
rect 194448 544170 194518 544226
rect 194574 544170 194642 544226
rect 194698 544170 194768 544226
rect 194448 544102 194768 544170
rect 194448 544046 194518 544102
rect 194574 544046 194642 544102
rect 194698 544046 194768 544102
rect 194448 543978 194768 544046
rect 194448 543922 194518 543978
rect 194574 543922 194642 543978
rect 194698 543922 194768 543978
rect 194448 543888 194768 543922
rect 225168 544350 225488 544384
rect 225168 544294 225238 544350
rect 225294 544294 225362 544350
rect 225418 544294 225488 544350
rect 225168 544226 225488 544294
rect 225168 544170 225238 544226
rect 225294 544170 225362 544226
rect 225418 544170 225488 544226
rect 225168 544102 225488 544170
rect 225168 544046 225238 544102
rect 225294 544046 225362 544102
rect 225418 544046 225488 544102
rect 225168 543978 225488 544046
rect 225168 543922 225238 543978
rect 225294 543922 225362 543978
rect 225418 543922 225488 543978
rect 225168 543888 225488 543922
rect 255888 544350 256208 544384
rect 255888 544294 255958 544350
rect 256014 544294 256082 544350
rect 256138 544294 256208 544350
rect 255888 544226 256208 544294
rect 255888 544170 255958 544226
rect 256014 544170 256082 544226
rect 256138 544170 256208 544226
rect 255888 544102 256208 544170
rect 255888 544046 255958 544102
rect 256014 544046 256082 544102
rect 256138 544046 256208 544102
rect 255888 543978 256208 544046
rect 255888 543922 255958 543978
rect 256014 543922 256082 543978
rect 256138 543922 256208 543978
rect 255888 543888 256208 543922
rect 286608 544350 286928 544384
rect 286608 544294 286678 544350
rect 286734 544294 286802 544350
rect 286858 544294 286928 544350
rect 286608 544226 286928 544294
rect 286608 544170 286678 544226
rect 286734 544170 286802 544226
rect 286858 544170 286928 544226
rect 286608 544102 286928 544170
rect 286608 544046 286678 544102
rect 286734 544046 286802 544102
rect 286858 544046 286928 544102
rect 286608 543978 286928 544046
rect 286608 543922 286678 543978
rect 286734 543922 286802 543978
rect 286858 543922 286928 543978
rect 286608 543888 286928 543922
rect 317328 544350 317648 544384
rect 317328 544294 317398 544350
rect 317454 544294 317522 544350
rect 317578 544294 317648 544350
rect 317328 544226 317648 544294
rect 317328 544170 317398 544226
rect 317454 544170 317522 544226
rect 317578 544170 317648 544226
rect 317328 544102 317648 544170
rect 317328 544046 317398 544102
rect 317454 544046 317522 544102
rect 317578 544046 317648 544102
rect 317328 543978 317648 544046
rect 317328 543922 317398 543978
rect 317454 543922 317522 543978
rect 317578 543922 317648 543978
rect 317328 543888 317648 543922
rect 348048 544350 348368 544384
rect 348048 544294 348118 544350
rect 348174 544294 348242 544350
rect 348298 544294 348368 544350
rect 348048 544226 348368 544294
rect 348048 544170 348118 544226
rect 348174 544170 348242 544226
rect 348298 544170 348368 544226
rect 348048 544102 348368 544170
rect 348048 544046 348118 544102
rect 348174 544046 348242 544102
rect 348298 544046 348368 544102
rect 348048 543978 348368 544046
rect 348048 543922 348118 543978
rect 348174 543922 348242 543978
rect 348298 543922 348368 543978
rect 348048 543888 348368 543922
rect 378768 544350 379088 544384
rect 378768 544294 378838 544350
rect 378894 544294 378962 544350
rect 379018 544294 379088 544350
rect 378768 544226 379088 544294
rect 378768 544170 378838 544226
rect 378894 544170 378962 544226
rect 379018 544170 379088 544226
rect 378768 544102 379088 544170
rect 378768 544046 378838 544102
rect 378894 544046 378962 544102
rect 379018 544046 379088 544102
rect 378768 543978 379088 544046
rect 378768 543922 378838 543978
rect 378894 543922 378962 543978
rect 379018 543922 379088 543978
rect 378768 543888 379088 543922
rect 409488 544350 409808 544384
rect 409488 544294 409558 544350
rect 409614 544294 409682 544350
rect 409738 544294 409808 544350
rect 409488 544226 409808 544294
rect 409488 544170 409558 544226
rect 409614 544170 409682 544226
rect 409738 544170 409808 544226
rect 409488 544102 409808 544170
rect 409488 544046 409558 544102
rect 409614 544046 409682 544102
rect 409738 544046 409808 544102
rect 409488 543978 409808 544046
rect 409488 543922 409558 543978
rect 409614 543922 409682 543978
rect 409738 543922 409808 543978
rect 409488 543888 409808 543922
rect 440208 544350 440528 544384
rect 440208 544294 440278 544350
rect 440334 544294 440402 544350
rect 440458 544294 440528 544350
rect 440208 544226 440528 544294
rect 440208 544170 440278 544226
rect 440334 544170 440402 544226
rect 440458 544170 440528 544226
rect 440208 544102 440528 544170
rect 440208 544046 440278 544102
rect 440334 544046 440402 544102
rect 440458 544046 440528 544102
rect 440208 543978 440528 544046
rect 440208 543922 440278 543978
rect 440334 543922 440402 543978
rect 440458 543922 440528 543978
rect 440208 543888 440528 543922
rect 470928 544350 471248 544384
rect 470928 544294 470998 544350
rect 471054 544294 471122 544350
rect 471178 544294 471248 544350
rect 470928 544226 471248 544294
rect 470928 544170 470998 544226
rect 471054 544170 471122 544226
rect 471178 544170 471248 544226
rect 470928 544102 471248 544170
rect 470928 544046 470998 544102
rect 471054 544046 471122 544102
rect 471178 544046 471248 544102
rect 470928 543978 471248 544046
rect 470928 543922 470998 543978
rect 471054 543922 471122 543978
rect 471178 543922 471248 543978
rect 470928 543888 471248 543922
rect 501648 544350 501968 544384
rect 501648 544294 501718 544350
rect 501774 544294 501842 544350
rect 501898 544294 501968 544350
rect 501648 544226 501968 544294
rect 501648 544170 501718 544226
rect 501774 544170 501842 544226
rect 501898 544170 501968 544226
rect 501648 544102 501968 544170
rect 501648 544046 501718 544102
rect 501774 544046 501842 544102
rect 501898 544046 501968 544102
rect 501648 543978 501968 544046
rect 501648 543922 501718 543978
rect 501774 543922 501842 543978
rect 501898 543922 501968 543978
rect 501648 543888 501968 543922
rect 209808 532350 210128 532384
rect 209808 532294 209878 532350
rect 209934 532294 210002 532350
rect 210058 532294 210128 532350
rect 209808 532226 210128 532294
rect 209808 532170 209878 532226
rect 209934 532170 210002 532226
rect 210058 532170 210128 532226
rect 209808 532102 210128 532170
rect 209808 532046 209878 532102
rect 209934 532046 210002 532102
rect 210058 532046 210128 532102
rect 209808 531978 210128 532046
rect 209808 531922 209878 531978
rect 209934 531922 210002 531978
rect 210058 531922 210128 531978
rect 209808 531888 210128 531922
rect 240528 532350 240848 532384
rect 240528 532294 240598 532350
rect 240654 532294 240722 532350
rect 240778 532294 240848 532350
rect 240528 532226 240848 532294
rect 240528 532170 240598 532226
rect 240654 532170 240722 532226
rect 240778 532170 240848 532226
rect 240528 532102 240848 532170
rect 240528 532046 240598 532102
rect 240654 532046 240722 532102
rect 240778 532046 240848 532102
rect 240528 531978 240848 532046
rect 240528 531922 240598 531978
rect 240654 531922 240722 531978
rect 240778 531922 240848 531978
rect 240528 531888 240848 531922
rect 271248 532350 271568 532384
rect 271248 532294 271318 532350
rect 271374 532294 271442 532350
rect 271498 532294 271568 532350
rect 271248 532226 271568 532294
rect 271248 532170 271318 532226
rect 271374 532170 271442 532226
rect 271498 532170 271568 532226
rect 271248 532102 271568 532170
rect 271248 532046 271318 532102
rect 271374 532046 271442 532102
rect 271498 532046 271568 532102
rect 271248 531978 271568 532046
rect 271248 531922 271318 531978
rect 271374 531922 271442 531978
rect 271498 531922 271568 531978
rect 271248 531888 271568 531922
rect 301968 532350 302288 532384
rect 301968 532294 302038 532350
rect 302094 532294 302162 532350
rect 302218 532294 302288 532350
rect 301968 532226 302288 532294
rect 301968 532170 302038 532226
rect 302094 532170 302162 532226
rect 302218 532170 302288 532226
rect 301968 532102 302288 532170
rect 301968 532046 302038 532102
rect 302094 532046 302162 532102
rect 302218 532046 302288 532102
rect 301968 531978 302288 532046
rect 301968 531922 302038 531978
rect 302094 531922 302162 531978
rect 302218 531922 302288 531978
rect 301968 531888 302288 531922
rect 332688 532350 333008 532384
rect 332688 532294 332758 532350
rect 332814 532294 332882 532350
rect 332938 532294 333008 532350
rect 332688 532226 333008 532294
rect 332688 532170 332758 532226
rect 332814 532170 332882 532226
rect 332938 532170 333008 532226
rect 332688 532102 333008 532170
rect 332688 532046 332758 532102
rect 332814 532046 332882 532102
rect 332938 532046 333008 532102
rect 332688 531978 333008 532046
rect 332688 531922 332758 531978
rect 332814 531922 332882 531978
rect 332938 531922 333008 531978
rect 332688 531888 333008 531922
rect 363408 532350 363728 532384
rect 363408 532294 363478 532350
rect 363534 532294 363602 532350
rect 363658 532294 363728 532350
rect 363408 532226 363728 532294
rect 363408 532170 363478 532226
rect 363534 532170 363602 532226
rect 363658 532170 363728 532226
rect 363408 532102 363728 532170
rect 363408 532046 363478 532102
rect 363534 532046 363602 532102
rect 363658 532046 363728 532102
rect 363408 531978 363728 532046
rect 363408 531922 363478 531978
rect 363534 531922 363602 531978
rect 363658 531922 363728 531978
rect 363408 531888 363728 531922
rect 394128 532350 394448 532384
rect 394128 532294 394198 532350
rect 394254 532294 394322 532350
rect 394378 532294 394448 532350
rect 394128 532226 394448 532294
rect 394128 532170 394198 532226
rect 394254 532170 394322 532226
rect 394378 532170 394448 532226
rect 394128 532102 394448 532170
rect 394128 532046 394198 532102
rect 394254 532046 394322 532102
rect 394378 532046 394448 532102
rect 394128 531978 394448 532046
rect 394128 531922 394198 531978
rect 394254 531922 394322 531978
rect 394378 531922 394448 531978
rect 394128 531888 394448 531922
rect 424848 532350 425168 532384
rect 424848 532294 424918 532350
rect 424974 532294 425042 532350
rect 425098 532294 425168 532350
rect 424848 532226 425168 532294
rect 424848 532170 424918 532226
rect 424974 532170 425042 532226
rect 425098 532170 425168 532226
rect 424848 532102 425168 532170
rect 424848 532046 424918 532102
rect 424974 532046 425042 532102
rect 425098 532046 425168 532102
rect 424848 531978 425168 532046
rect 424848 531922 424918 531978
rect 424974 531922 425042 531978
rect 425098 531922 425168 531978
rect 424848 531888 425168 531922
rect 455568 532350 455888 532384
rect 455568 532294 455638 532350
rect 455694 532294 455762 532350
rect 455818 532294 455888 532350
rect 455568 532226 455888 532294
rect 455568 532170 455638 532226
rect 455694 532170 455762 532226
rect 455818 532170 455888 532226
rect 455568 532102 455888 532170
rect 455568 532046 455638 532102
rect 455694 532046 455762 532102
rect 455818 532046 455888 532102
rect 455568 531978 455888 532046
rect 455568 531922 455638 531978
rect 455694 531922 455762 531978
rect 455818 531922 455888 531978
rect 455568 531888 455888 531922
rect 486288 532350 486608 532384
rect 486288 532294 486358 532350
rect 486414 532294 486482 532350
rect 486538 532294 486608 532350
rect 486288 532226 486608 532294
rect 486288 532170 486358 532226
rect 486414 532170 486482 532226
rect 486538 532170 486608 532226
rect 486288 532102 486608 532170
rect 486288 532046 486358 532102
rect 486414 532046 486482 532102
rect 486538 532046 486608 532102
rect 486288 531978 486608 532046
rect 486288 531922 486358 531978
rect 486414 531922 486482 531978
rect 486538 531922 486608 531978
rect 486288 531888 486608 531922
rect 194448 526350 194768 526384
rect 194448 526294 194518 526350
rect 194574 526294 194642 526350
rect 194698 526294 194768 526350
rect 194448 526226 194768 526294
rect 194448 526170 194518 526226
rect 194574 526170 194642 526226
rect 194698 526170 194768 526226
rect 194448 526102 194768 526170
rect 194448 526046 194518 526102
rect 194574 526046 194642 526102
rect 194698 526046 194768 526102
rect 194448 525978 194768 526046
rect 194448 525922 194518 525978
rect 194574 525922 194642 525978
rect 194698 525922 194768 525978
rect 194448 525888 194768 525922
rect 225168 526350 225488 526384
rect 225168 526294 225238 526350
rect 225294 526294 225362 526350
rect 225418 526294 225488 526350
rect 225168 526226 225488 526294
rect 225168 526170 225238 526226
rect 225294 526170 225362 526226
rect 225418 526170 225488 526226
rect 225168 526102 225488 526170
rect 225168 526046 225238 526102
rect 225294 526046 225362 526102
rect 225418 526046 225488 526102
rect 225168 525978 225488 526046
rect 225168 525922 225238 525978
rect 225294 525922 225362 525978
rect 225418 525922 225488 525978
rect 225168 525888 225488 525922
rect 255888 526350 256208 526384
rect 255888 526294 255958 526350
rect 256014 526294 256082 526350
rect 256138 526294 256208 526350
rect 255888 526226 256208 526294
rect 255888 526170 255958 526226
rect 256014 526170 256082 526226
rect 256138 526170 256208 526226
rect 255888 526102 256208 526170
rect 255888 526046 255958 526102
rect 256014 526046 256082 526102
rect 256138 526046 256208 526102
rect 255888 525978 256208 526046
rect 255888 525922 255958 525978
rect 256014 525922 256082 525978
rect 256138 525922 256208 525978
rect 255888 525888 256208 525922
rect 286608 526350 286928 526384
rect 286608 526294 286678 526350
rect 286734 526294 286802 526350
rect 286858 526294 286928 526350
rect 286608 526226 286928 526294
rect 286608 526170 286678 526226
rect 286734 526170 286802 526226
rect 286858 526170 286928 526226
rect 286608 526102 286928 526170
rect 286608 526046 286678 526102
rect 286734 526046 286802 526102
rect 286858 526046 286928 526102
rect 286608 525978 286928 526046
rect 286608 525922 286678 525978
rect 286734 525922 286802 525978
rect 286858 525922 286928 525978
rect 286608 525888 286928 525922
rect 317328 526350 317648 526384
rect 317328 526294 317398 526350
rect 317454 526294 317522 526350
rect 317578 526294 317648 526350
rect 317328 526226 317648 526294
rect 317328 526170 317398 526226
rect 317454 526170 317522 526226
rect 317578 526170 317648 526226
rect 317328 526102 317648 526170
rect 317328 526046 317398 526102
rect 317454 526046 317522 526102
rect 317578 526046 317648 526102
rect 317328 525978 317648 526046
rect 317328 525922 317398 525978
rect 317454 525922 317522 525978
rect 317578 525922 317648 525978
rect 317328 525888 317648 525922
rect 348048 526350 348368 526384
rect 348048 526294 348118 526350
rect 348174 526294 348242 526350
rect 348298 526294 348368 526350
rect 348048 526226 348368 526294
rect 348048 526170 348118 526226
rect 348174 526170 348242 526226
rect 348298 526170 348368 526226
rect 348048 526102 348368 526170
rect 348048 526046 348118 526102
rect 348174 526046 348242 526102
rect 348298 526046 348368 526102
rect 348048 525978 348368 526046
rect 348048 525922 348118 525978
rect 348174 525922 348242 525978
rect 348298 525922 348368 525978
rect 348048 525888 348368 525922
rect 378768 526350 379088 526384
rect 378768 526294 378838 526350
rect 378894 526294 378962 526350
rect 379018 526294 379088 526350
rect 378768 526226 379088 526294
rect 378768 526170 378838 526226
rect 378894 526170 378962 526226
rect 379018 526170 379088 526226
rect 378768 526102 379088 526170
rect 378768 526046 378838 526102
rect 378894 526046 378962 526102
rect 379018 526046 379088 526102
rect 378768 525978 379088 526046
rect 378768 525922 378838 525978
rect 378894 525922 378962 525978
rect 379018 525922 379088 525978
rect 378768 525888 379088 525922
rect 409488 526350 409808 526384
rect 409488 526294 409558 526350
rect 409614 526294 409682 526350
rect 409738 526294 409808 526350
rect 409488 526226 409808 526294
rect 409488 526170 409558 526226
rect 409614 526170 409682 526226
rect 409738 526170 409808 526226
rect 409488 526102 409808 526170
rect 409488 526046 409558 526102
rect 409614 526046 409682 526102
rect 409738 526046 409808 526102
rect 409488 525978 409808 526046
rect 409488 525922 409558 525978
rect 409614 525922 409682 525978
rect 409738 525922 409808 525978
rect 409488 525888 409808 525922
rect 440208 526350 440528 526384
rect 440208 526294 440278 526350
rect 440334 526294 440402 526350
rect 440458 526294 440528 526350
rect 440208 526226 440528 526294
rect 440208 526170 440278 526226
rect 440334 526170 440402 526226
rect 440458 526170 440528 526226
rect 440208 526102 440528 526170
rect 440208 526046 440278 526102
rect 440334 526046 440402 526102
rect 440458 526046 440528 526102
rect 440208 525978 440528 526046
rect 440208 525922 440278 525978
rect 440334 525922 440402 525978
rect 440458 525922 440528 525978
rect 440208 525888 440528 525922
rect 470928 526350 471248 526384
rect 470928 526294 470998 526350
rect 471054 526294 471122 526350
rect 471178 526294 471248 526350
rect 470928 526226 471248 526294
rect 470928 526170 470998 526226
rect 471054 526170 471122 526226
rect 471178 526170 471248 526226
rect 470928 526102 471248 526170
rect 470928 526046 470998 526102
rect 471054 526046 471122 526102
rect 471178 526046 471248 526102
rect 470928 525978 471248 526046
rect 470928 525922 470998 525978
rect 471054 525922 471122 525978
rect 471178 525922 471248 525978
rect 470928 525888 471248 525922
rect 501648 526350 501968 526384
rect 501648 526294 501718 526350
rect 501774 526294 501842 526350
rect 501898 526294 501968 526350
rect 501648 526226 501968 526294
rect 501648 526170 501718 526226
rect 501774 526170 501842 526226
rect 501898 526170 501968 526226
rect 501648 526102 501968 526170
rect 501648 526046 501718 526102
rect 501774 526046 501842 526102
rect 501898 526046 501968 526102
rect 501648 525978 501968 526046
rect 501648 525922 501718 525978
rect 501774 525922 501842 525978
rect 501898 525922 501968 525978
rect 501648 525888 501968 525922
rect 209808 514350 210128 514384
rect 209808 514294 209878 514350
rect 209934 514294 210002 514350
rect 210058 514294 210128 514350
rect 209808 514226 210128 514294
rect 209808 514170 209878 514226
rect 209934 514170 210002 514226
rect 210058 514170 210128 514226
rect 209808 514102 210128 514170
rect 209808 514046 209878 514102
rect 209934 514046 210002 514102
rect 210058 514046 210128 514102
rect 209808 513978 210128 514046
rect 209808 513922 209878 513978
rect 209934 513922 210002 513978
rect 210058 513922 210128 513978
rect 209808 513888 210128 513922
rect 240528 514350 240848 514384
rect 240528 514294 240598 514350
rect 240654 514294 240722 514350
rect 240778 514294 240848 514350
rect 240528 514226 240848 514294
rect 240528 514170 240598 514226
rect 240654 514170 240722 514226
rect 240778 514170 240848 514226
rect 240528 514102 240848 514170
rect 240528 514046 240598 514102
rect 240654 514046 240722 514102
rect 240778 514046 240848 514102
rect 240528 513978 240848 514046
rect 240528 513922 240598 513978
rect 240654 513922 240722 513978
rect 240778 513922 240848 513978
rect 240528 513888 240848 513922
rect 271248 514350 271568 514384
rect 271248 514294 271318 514350
rect 271374 514294 271442 514350
rect 271498 514294 271568 514350
rect 271248 514226 271568 514294
rect 271248 514170 271318 514226
rect 271374 514170 271442 514226
rect 271498 514170 271568 514226
rect 271248 514102 271568 514170
rect 271248 514046 271318 514102
rect 271374 514046 271442 514102
rect 271498 514046 271568 514102
rect 271248 513978 271568 514046
rect 271248 513922 271318 513978
rect 271374 513922 271442 513978
rect 271498 513922 271568 513978
rect 271248 513888 271568 513922
rect 301968 514350 302288 514384
rect 301968 514294 302038 514350
rect 302094 514294 302162 514350
rect 302218 514294 302288 514350
rect 301968 514226 302288 514294
rect 301968 514170 302038 514226
rect 302094 514170 302162 514226
rect 302218 514170 302288 514226
rect 301968 514102 302288 514170
rect 301968 514046 302038 514102
rect 302094 514046 302162 514102
rect 302218 514046 302288 514102
rect 301968 513978 302288 514046
rect 301968 513922 302038 513978
rect 302094 513922 302162 513978
rect 302218 513922 302288 513978
rect 301968 513888 302288 513922
rect 332688 514350 333008 514384
rect 332688 514294 332758 514350
rect 332814 514294 332882 514350
rect 332938 514294 333008 514350
rect 332688 514226 333008 514294
rect 332688 514170 332758 514226
rect 332814 514170 332882 514226
rect 332938 514170 333008 514226
rect 332688 514102 333008 514170
rect 332688 514046 332758 514102
rect 332814 514046 332882 514102
rect 332938 514046 333008 514102
rect 332688 513978 333008 514046
rect 332688 513922 332758 513978
rect 332814 513922 332882 513978
rect 332938 513922 333008 513978
rect 332688 513888 333008 513922
rect 363408 514350 363728 514384
rect 363408 514294 363478 514350
rect 363534 514294 363602 514350
rect 363658 514294 363728 514350
rect 363408 514226 363728 514294
rect 363408 514170 363478 514226
rect 363534 514170 363602 514226
rect 363658 514170 363728 514226
rect 363408 514102 363728 514170
rect 363408 514046 363478 514102
rect 363534 514046 363602 514102
rect 363658 514046 363728 514102
rect 363408 513978 363728 514046
rect 363408 513922 363478 513978
rect 363534 513922 363602 513978
rect 363658 513922 363728 513978
rect 363408 513888 363728 513922
rect 394128 514350 394448 514384
rect 394128 514294 394198 514350
rect 394254 514294 394322 514350
rect 394378 514294 394448 514350
rect 394128 514226 394448 514294
rect 394128 514170 394198 514226
rect 394254 514170 394322 514226
rect 394378 514170 394448 514226
rect 394128 514102 394448 514170
rect 394128 514046 394198 514102
rect 394254 514046 394322 514102
rect 394378 514046 394448 514102
rect 394128 513978 394448 514046
rect 394128 513922 394198 513978
rect 394254 513922 394322 513978
rect 394378 513922 394448 513978
rect 394128 513888 394448 513922
rect 424848 514350 425168 514384
rect 424848 514294 424918 514350
rect 424974 514294 425042 514350
rect 425098 514294 425168 514350
rect 424848 514226 425168 514294
rect 424848 514170 424918 514226
rect 424974 514170 425042 514226
rect 425098 514170 425168 514226
rect 424848 514102 425168 514170
rect 424848 514046 424918 514102
rect 424974 514046 425042 514102
rect 425098 514046 425168 514102
rect 424848 513978 425168 514046
rect 424848 513922 424918 513978
rect 424974 513922 425042 513978
rect 425098 513922 425168 513978
rect 424848 513888 425168 513922
rect 455568 514350 455888 514384
rect 455568 514294 455638 514350
rect 455694 514294 455762 514350
rect 455818 514294 455888 514350
rect 455568 514226 455888 514294
rect 455568 514170 455638 514226
rect 455694 514170 455762 514226
rect 455818 514170 455888 514226
rect 455568 514102 455888 514170
rect 455568 514046 455638 514102
rect 455694 514046 455762 514102
rect 455818 514046 455888 514102
rect 455568 513978 455888 514046
rect 455568 513922 455638 513978
rect 455694 513922 455762 513978
rect 455818 513922 455888 513978
rect 455568 513888 455888 513922
rect 486288 514350 486608 514384
rect 486288 514294 486358 514350
rect 486414 514294 486482 514350
rect 486538 514294 486608 514350
rect 486288 514226 486608 514294
rect 486288 514170 486358 514226
rect 486414 514170 486482 514226
rect 486538 514170 486608 514226
rect 486288 514102 486608 514170
rect 486288 514046 486358 514102
rect 486414 514046 486482 514102
rect 486538 514046 486608 514102
rect 486288 513978 486608 514046
rect 486288 513922 486358 513978
rect 486414 513922 486482 513978
rect 486538 513922 486608 513978
rect 486288 513888 486608 513922
rect 194448 508350 194768 508384
rect 194448 508294 194518 508350
rect 194574 508294 194642 508350
rect 194698 508294 194768 508350
rect 194448 508226 194768 508294
rect 194448 508170 194518 508226
rect 194574 508170 194642 508226
rect 194698 508170 194768 508226
rect 194448 508102 194768 508170
rect 194448 508046 194518 508102
rect 194574 508046 194642 508102
rect 194698 508046 194768 508102
rect 194448 507978 194768 508046
rect 194448 507922 194518 507978
rect 194574 507922 194642 507978
rect 194698 507922 194768 507978
rect 194448 507888 194768 507922
rect 225168 508350 225488 508384
rect 225168 508294 225238 508350
rect 225294 508294 225362 508350
rect 225418 508294 225488 508350
rect 225168 508226 225488 508294
rect 225168 508170 225238 508226
rect 225294 508170 225362 508226
rect 225418 508170 225488 508226
rect 225168 508102 225488 508170
rect 225168 508046 225238 508102
rect 225294 508046 225362 508102
rect 225418 508046 225488 508102
rect 225168 507978 225488 508046
rect 225168 507922 225238 507978
rect 225294 507922 225362 507978
rect 225418 507922 225488 507978
rect 225168 507888 225488 507922
rect 255888 508350 256208 508384
rect 255888 508294 255958 508350
rect 256014 508294 256082 508350
rect 256138 508294 256208 508350
rect 255888 508226 256208 508294
rect 255888 508170 255958 508226
rect 256014 508170 256082 508226
rect 256138 508170 256208 508226
rect 255888 508102 256208 508170
rect 255888 508046 255958 508102
rect 256014 508046 256082 508102
rect 256138 508046 256208 508102
rect 255888 507978 256208 508046
rect 255888 507922 255958 507978
rect 256014 507922 256082 507978
rect 256138 507922 256208 507978
rect 255888 507888 256208 507922
rect 286608 508350 286928 508384
rect 286608 508294 286678 508350
rect 286734 508294 286802 508350
rect 286858 508294 286928 508350
rect 286608 508226 286928 508294
rect 286608 508170 286678 508226
rect 286734 508170 286802 508226
rect 286858 508170 286928 508226
rect 286608 508102 286928 508170
rect 286608 508046 286678 508102
rect 286734 508046 286802 508102
rect 286858 508046 286928 508102
rect 286608 507978 286928 508046
rect 286608 507922 286678 507978
rect 286734 507922 286802 507978
rect 286858 507922 286928 507978
rect 286608 507888 286928 507922
rect 317328 508350 317648 508384
rect 317328 508294 317398 508350
rect 317454 508294 317522 508350
rect 317578 508294 317648 508350
rect 317328 508226 317648 508294
rect 317328 508170 317398 508226
rect 317454 508170 317522 508226
rect 317578 508170 317648 508226
rect 317328 508102 317648 508170
rect 317328 508046 317398 508102
rect 317454 508046 317522 508102
rect 317578 508046 317648 508102
rect 317328 507978 317648 508046
rect 317328 507922 317398 507978
rect 317454 507922 317522 507978
rect 317578 507922 317648 507978
rect 317328 507888 317648 507922
rect 348048 508350 348368 508384
rect 348048 508294 348118 508350
rect 348174 508294 348242 508350
rect 348298 508294 348368 508350
rect 348048 508226 348368 508294
rect 348048 508170 348118 508226
rect 348174 508170 348242 508226
rect 348298 508170 348368 508226
rect 348048 508102 348368 508170
rect 348048 508046 348118 508102
rect 348174 508046 348242 508102
rect 348298 508046 348368 508102
rect 348048 507978 348368 508046
rect 348048 507922 348118 507978
rect 348174 507922 348242 507978
rect 348298 507922 348368 507978
rect 348048 507888 348368 507922
rect 378768 508350 379088 508384
rect 378768 508294 378838 508350
rect 378894 508294 378962 508350
rect 379018 508294 379088 508350
rect 378768 508226 379088 508294
rect 378768 508170 378838 508226
rect 378894 508170 378962 508226
rect 379018 508170 379088 508226
rect 378768 508102 379088 508170
rect 378768 508046 378838 508102
rect 378894 508046 378962 508102
rect 379018 508046 379088 508102
rect 378768 507978 379088 508046
rect 378768 507922 378838 507978
rect 378894 507922 378962 507978
rect 379018 507922 379088 507978
rect 378768 507888 379088 507922
rect 409488 508350 409808 508384
rect 409488 508294 409558 508350
rect 409614 508294 409682 508350
rect 409738 508294 409808 508350
rect 409488 508226 409808 508294
rect 409488 508170 409558 508226
rect 409614 508170 409682 508226
rect 409738 508170 409808 508226
rect 409488 508102 409808 508170
rect 409488 508046 409558 508102
rect 409614 508046 409682 508102
rect 409738 508046 409808 508102
rect 409488 507978 409808 508046
rect 409488 507922 409558 507978
rect 409614 507922 409682 507978
rect 409738 507922 409808 507978
rect 409488 507888 409808 507922
rect 440208 508350 440528 508384
rect 440208 508294 440278 508350
rect 440334 508294 440402 508350
rect 440458 508294 440528 508350
rect 440208 508226 440528 508294
rect 440208 508170 440278 508226
rect 440334 508170 440402 508226
rect 440458 508170 440528 508226
rect 440208 508102 440528 508170
rect 440208 508046 440278 508102
rect 440334 508046 440402 508102
rect 440458 508046 440528 508102
rect 440208 507978 440528 508046
rect 440208 507922 440278 507978
rect 440334 507922 440402 507978
rect 440458 507922 440528 507978
rect 440208 507888 440528 507922
rect 470928 508350 471248 508384
rect 470928 508294 470998 508350
rect 471054 508294 471122 508350
rect 471178 508294 471248 508350
rect 470928 508226 471248 508294
rect 470928 508170 470998 508226
rect 471054 508170 471122 508226
rect 471178 508170 471248 508226
rect 470928 508102 471248 508170
rect 470928 508046 470998 508102
rect 471054 508046 471122 508102
rect 471178 508046 471248 508102
rect 470928 507978 471248 508046
rect 470928 507922 470998 507978
rect 471054 507922 471122 507978
rect 471178 507922 471248 507978
rect 470928 507888 471248 507922
rect 501648 508350 501968 508384
rect 501648 508294 501718 508350
rect 501774 508294 501842 508350
rect 501898 508294 501968 508350
rect 501648 508226 501968 508294
rect 501648 508170 501718 508226
rect 501774 508170 501842 508226
rect 501898 508170 501968 508226
rect 501648 508102 501968 508170
rect 501648 508046 501718 508102
rect 501774 508046 501842 508102
rect 501898 508046 501968 508102
rect 501648 507978 501968 508046
rect 501648 507922 501718 507978
rect 501774 507922 501842 507978
rect 501898 507922 501968 507978
rect 501648 507888 501968 507922
rect 209808 496350 210128 496384
rect 209808 496294 209878 496350
rect 209934 496294 210002 496350
rect 210058 496294 210128 496350
rect 209808 496226 210128 496294
rect 209808 496170 209878 496226
rect 209934 496170 210002 496226
rect 210058 496170 210128 496226
rect 209808 496102 210128 496170
rect 209808 496046 209878 496102
rect 209934 496046 210002 496102
rect 210058 496046 210128 496102
rect 209808 495978 210128 496046
rect 209808 495922 209878 495978
rect 209934 495922 210002 495978
rect 210058 495922 210128 495978
rect 209808 495888 210128 495922
rect 240528 496350 240848 496384
rect 240528 496294 240598 496350
rect 240654 496294 240722 496350
rect 240778 496294 240848 496350
rect 240528 496226 240848 496294
rect 240528 496170 240598 496226
rect 240654 496170 240722 496226
rect 240778 496170 240848 496226
rect 240528 496102 240848 496170
rect 240528 496046 240598 496102
rect 240654 496046 240722 496102
rect 240778 496046 240848 496102
rect 240528 495978 240848 496046
rect 240528 495922 240598 495978
rect 240654 495922 240722 495978
rect 240778 495922 240848 495978
rect 240528 495888 240848 495922
rect 271248 496350 271568 496384
rect 271248 496294 271318 496350
rect 271374 496294 271442 496350
rect 271498 496294 271568 496350
rect 271248 496226 271568 496294
rect 271248 496170 271318 496226
rect 271374 496170 271442 496226
rect 271498 496170 271568 496226
rect 271248 496102 271568 496170
rect 271248 496046 271318 496102
rect 271374 496046 271442 496102
rect 271498 496046 271568 496102
rect 271248 495978 271568 496046
rect 271248 495922 271318 495978
rect 271374 495922 271442 495978
rect 271498 495922 271568 495978
rect 271248 495888 271568 495922
rect 301968 496350 302288 496384
rect 301968 496294 302038 496350
rect 302094 496294 302162 496350
rect 302218 496294 302288 496350
rect 301968 496226 302288 496294
rect 301968 496170 302038 496226
rect 302094 496170 302162 496226
rect 302218 496170 302288 496226
rect 301968 496102 302288 496170
rect 301968 496046 302038 496102
rect 302094 496046 302162 496102
rect 302218 496046 302288 496102
rect 301968 495978 302288 496046
rect 301968 495922 302038 495978
rect 302094 495922 302162 495978
rect 302218 495922 302288 495978
rect 301968 495888 302288 495922
rect 332688 496350 333008 496384
rect 332688 496294 332758 496350
rect 332814 496294 332882 496350
rect 332938 496294 333008 496350
rect 332688 496226 333008 496294
rect 332688 496170 332758 496226
rect 332814 496170 332882 496226
rect 332938 496170 333008 496226
rect 332688 496102 333008 496170
rect 332688 496046 332758 496102
rect 332814 496046 332882 496102
rect 332938 496046 333008 496102
rect 332688 495978 333008 496046
rect 332688 495922 332758 495978
rect 332814 495922 332882 495978
rect 332938 495922 333008 495978
rect 332688 495888 333008 495922
rect 363408 496350 363728 496384
rect 363408 496294 363478 496350
rect 363534 496294 363602 496350
rect 363658 496294 363728 496350
rect 363408 496226 363728 496294
rect 363408 496170 363478 496226
rect 363534 496170 363602 496226
rect 363658 496170 363728 496226
rect 363408 496102 363728 496170
rect 363408 496046 363478 496102
rect 363534 496046 363602 496102
rect 363658 496046 363728 496102
rect 363408 495978 363728 496046
rect 363408 495922 363478 495978
rect 363534 495922 363602 495978
rect 363658 495922 363728 495978
rect 363408 495888 363728 495922
rect 394128 496350 394448 496384
rect 394128 496294 394198 496350
rect 394254 496294 394322 496350
rect 394378 496294 394448 496350
rect 394128 496226 394448 496294
rect 394128 496170 394198 496226
rect 394254 496170 394322 496226
rect 394378 496170 394448 496226
rect 394128 496102 394448 496170
rect 394128 496046 394198 496102
rect 394254 496046 394322 496102
rect 394378 496046 394448 496102
rect 394128 495978 394448 496046
rect 394128 495922 394198 495978
rect 394254 495922 394322 495978
rect 394378 495922 394448 495978
rect 394128 495888 394448 495922
rect 424848 496350 425168 496384
rect 424848 496294 424918 496350
rect 424974 496294 425042 496350
rect 425098 496294 425168 496350
rect 424848 496226 425168 496294
rect 424848 496170 424918 496226
rect 424974 496170 425042 496226
rect 425098 496170 425168 496226
rect 424848 496102 425168 496170
rect 424848 496046 424918 496102
rect 424974 496046 425042 496102
rect 425098 496046 425168 496102
rect 424848 495978 425168 496046
rect 424848 495922 424918 495978
rect 424974 495922 425042 495978
rect 425098 495922 425168 495978
rect 424848 495888 425168 495922
rect 455568 496350 455888 496384
rect 455568 496294 455638 496350
rect 455694 496294 455762 496350
rect 455818 496294 455888 496350
rect 455568 496226 455888 496294
rect 455568 496170 455638 496226
rect 455694 496170 455762 496226
rect 455818 496170 455888 496226
rect 455568 496102 455888 496170
rect 455568 496046 455638 496102
rect 455694 496046 455762 496102
rect 455818 496046 455888 496102
rect 455568 495978 455888 496046
rect 455568 495922 455638 495978
rect 455694 495922 455762 495978
rect 455818 495922 455888 495978
rect 455568 495888 455888 495922
rect 486288 496350 486608 496384
rect 486288 496294 486358 496350
rect 486414 496294 486482 496350
rect 486538 496294 486608 496350
rect 486288 496226 486608 496294
rect 486288 496170 486358 496226
rect 486414 496170 486482 496226
rect 486538 496170 486608 496226
rect 486288 496102 486608 496170
rect 486288 496046 486358 496102
rect 486414 496046 486482 496102
rect 486538 496046 486608 496102
rect 486288 495978 486608 496046
rect 486288 495922 486358 495978
rect 486414 495922 486482 495978
rect 486538 495922 486608 495978
rect 486288 495888 486608 495922
rect 194448 490350 194768 490384
rect 194448 490294 194518 490350
rect 194574 490294 194642 490350
rect 194698 490294 194768 490350
rect 194448 490226 194768 490294
rect 194448 490170 194518 490226
rect 194574 490170 194642 490226
rect 194698 490170 194768 490226
rect 194448 490102 194768 490170
rect 194448 490046 194518 490102
rect 194574 490046 194642 490102
rect 194698 490046 194768 490102
rect 194448 489978 194768 490046
rect 194448 489922 194518 489978
rect 194574 489922 194642 489978
rect 194698 489922 194768 489978
rect 194448 489888 194768 489922
rect 225168 490350 225488 490384
rect 225168 490294 225238 490350
rect 225294 490294 225362 490350
rect 225418 490294 225488 490350
rect 225168 490226 225488 490294
rect 225168 490170 225238 490226
rect 225294 490170 225362 490226
rect 225418 490170 225488 490226
rect 225168 490102 225488 490170
rect 225168 490046 225238 490102
rect 225294 490046 225362 490102
rect 225418 490046 225488 490102
rect 225168 489978 225488 490046
rect 225168 489922 225238 489978
rect 225294 489922 225362 489978
rect 225418 489922 225488 489978
rect 225168 489888 225488 489922
rect 255888 490350 256208 490384
rect 255888 490294 255958 490350
rect 256014 490294 256082 490350
rect 256138 490294 256208 490350
rect 255888 490226 256208 490294
rect 255888 490170 255958 490226
rect 256014 490170 256082 490226
rect 256138 490170 256208 490226
rect 255888 490102 256208 490170
rect 255888 490046 255958 490102
rect 256014 490046 256082 490102
rect 256138 490046 256208 490102
rect 255888 489978 256208 490046
rect 255888 489922 255958 489978
rect 256014 489922 256082 489978
rect 256138 489922 256208 489978
rect 255888 489888 256208 489922
rect 286608 490350 286928 490384
rect 286608 490294 286678 490350
rect 286734 490294 286802 490350
rect 286858 490294 286928 490350
rect 286608 490226 286928 490294
rect 286608 490170 286678 490226
rect 286734 490170 286802 490226
rect 286858 490170 286928 490226
rect 286608 490102 286928 490170
rect 286608 490046 286678 490102
rect 286734 490046 286802 490102
rect 286858 490046 286928 490102
rect 286608 489978 286928 490046
rect 286608 489922 286678 489978
rect 286734 489922 286802 489978
rect 286858 489922 286928 489978
rect 286608 489888 286928 489922
rect 317328 490350 317648 490384
rect 317328 490294 317398 490350
rect 317454 490294 317522 490350
rect 317578 490294 317648 490350
rect 317328 490226 317648 490294
rect 317328 490170 317398 490226
rect 317454 490170 317522 490226
rect 317578 490170 317648 490226
rect 317328 490102 317648 490170
rect 317328 490046 317398 490102
rect 317454 490046 317522 490102
rect 317578 490046 317648 490102
rect 317328 489978 317648 490046
rect 317328 489922 317398 489978
rect 317454 489922 317522 489978
rect 317578 489922 317648 489978
rect 317328 489888 317648 489922
rect 348048 490350 348368 490384
rect 348048 490294 348118 490350
rect 348174 490294 348242 490350
rect 348298 490294 348368 490350
rect 348048 490226 348368 490294
rect 348048 490170 348118 490226
rect 348174 490170 348242 490226
rect 348298 490170 348368 490226
rect 348048 490102 348368 490170
rect 348048 490046 348118 490102
rect 348174 490046 348242 490102
rect 348298 490046 348368 490102
rect 348048 489978 348368 490046
rect 348048 489922 348118 489978
rect 348174 489922 348242 489978
rect 348298 489922 348368 489978
rect 348048 489888 348368 489922
rect 378768 490350 379088 490384
rect 378768 490294 378838 490350
rect 378894 490294 378962 490350
rect 379018 490294 379088 490350
rect 378768 490226 379088 490294
rect 378768 490170 378838 490226
rect 378894 490170 378962 490226
rect 379018 490170 379088 490226
rect 378768 490102 379088 490170
rect 378768 490046 378838 490102
rect 378894 490046 378962 490102
rect 379018 490046 379088 490102
rect 378768 489978 379088 490046
rect 378768 489922 378838 489978
rect 378894 489922 378962 489978
rect 379018 489922 379088 489978
rect 378768 489888 379088 489922
rect 409488 490350 409808 490384
rect 409488 490294 409558 490350
rect 409614 490294 409682 490350
rect 409738 490294 409808 490350
rect 409488 490226 409808 490294
rect 409488 490170 409558 490226
rect 409614 490170 409682 490226
rect 409738 490170 409808 490226
rect 409488 490102 409808 490170
rect 409488 490046 409558 490102
rect 409614 490046 409682 490102
rect 409738 490046 409808 490102
rect 409488 489978 409808 490046
rect 409488 489922 409558 489978
rect 409614 489922 409682 489978
rect 409738 489922 409808 489978
rect 409488 489888 409808 489922
rect 440208 490350 440528 490384
rect 440208 490294 440278 490350
rect 440334 490294 440402 490350
rect 440458 490294 440528 490350
rect 440208 490226 440528 490294
rect 440208 490170 440278 490226
rect 440334 490170 440402 490226
rect 440458 490170 440528 490226
rect 440208 490102 440528 490170
rect 440208 490046 440278 490102
rect 440334 490046 440402 490102
rect 440458 490046 440528 490102
rect 440208 489978 440528 490046
rect 440208 489922 440278 489978
rect 440334 489922 440402 489978
rect 440458 489922 440528 489978
rect 440208 489888 440528 489922
rect 470928 490350 471248 490384
rect 470928 490294 470998 490350
rect 471054 490294 471122 490350
rect 471178 490294 471248 490350
rect 470928 490226 471248 490294
rect 470928 490170 470998 490226
rect 471054 490170 471122 490226
rect 471178 490170 471248 490226
rect 470928 490102 471248 490170
rect 470928 490046 470998 490102
rect 471054 490046 471122 490102
rect 471178 490046 471248 490102
rect 470928 489978 471248 490046
rect 470928 489922 470998 489978
rect 471054 489922 471122 489978
rect 471178 489922 471248 489978
rect 470928 489888 471248 489922
rect 501648 490350 501968 490384
rect 501648 490294 501718 490350
rect 501774 490294 501842 490350
rect 501898 490294 501968 490350
rect 501648 490226 501968 490294
rect 501648 490170 501718 490226
rect 501774 490170 501842 490226
rect 501898 490170 501968 490226
rect 501648 490102 501968 490170
rect 501648 490046 501718 490102
rect 501774 490046 501842 490102
rect 501898 490046 501968 490102
rect 501648 489978 501968 490046
rect 501648 489922 501718 489978
rect 501774 489922 501842 489978
rect 501898 489922 501968 489978
rect 501648 489888 501968 489922
rect 209808 478350 210128 478384
rect 209808 478294 209878 478350
rect 209934 478294 210002 478350
rect 210058 478294 210128 478350
rect 209808 478226 210128 478294
rect 209808 478170 209878 478226
rect 209934 478170 210002 478226
rect 210058 478170 210128 478226
rect 209808 478102 210128 478170
rect 209808 478046 209878 478102
rect 209934 478046 210002 478102
rect 210058 478046 210128 478102
rect 209808 477978 210128 478046
rect 209808 477922 209878 477978
rect 209934 477922 210002 477978
rect 210058 477922 210128 477978
rect 209808 477888 210128 477922
rect 240528 478350 240848 478384
rect 240528 478294 240598 478350
rect 240654 478294 240722 478350
rect 240778 478294 240848 478350
rect 240528 478226 240848 478294
rect 240528 478170 240598 478226
rect 240654 478170 240722 478226
rect 240778 478170 240848 478226
rect 240528 478102 240848 478170
rect 240528 478046 240598 478102
rect 240654 478046 240722 478102
rect 240778 478046 240848 478102
rect 240528 477978 240848 478046
rect 240528 477922 240598 477978
rect 240654 477922 240722 477978
rect 240778 477922 240848 477978
rect 240528 477888 240848 477922
rect 271248 478350 271568 478384
rect 271248 478294 271318 478350
rect 271374 478294 271442 478350
rect 271498 478294 271568 478350
rect 271248 478226 271568 478294
rect 271248 478170 271318 478226
rect 271374 478170 271442 478226
rect 271498 478170 271568 478226
rect 271248 478102 271568 478170
rect 271248 478046 271318 478102
rect 271374 478046 271442 478102
rect 271498 478046 271568 478102
rect 271248 477978 271568 478046
rect 271248 477922 271318 477978
rect 271374 477922 271442 477978
rect 271498 477922 271568 477978
rect 271248 477888 271568 477922
rect 301968 478350 302288 478384
rect 301968 478294 302038 478350
rect 302094 478294 302162 478350
rect 302218 478294 302288 478350
rect 301968 478226 302288 478294
rect 301968 478170 302038 478226
rect 302094 478170 302162 478226
rect 302218 478170 302288 478226
rect 301968 478102 302288 478170
rect 301968 478046 302038 478102
rect 302094 478046 302162 478102
rect 302218 478046 302288 478102
rect 301968 477978 302288 478046
rect 301968 477922 302038 477978
rect 302094 477922 302162 477978
rect 302218 477922 302288 477978
rect 301968 477888 302288 477922
rect 332688 478350 333008 478384
rect 332688 478294 332758 478350
rect 332814 478294 332882 478350
rect 332938 478294 333008 478350
rect 332688 478226 333008 478294
rect 332688 478170 332758 478226
rect 332814 478170 332882 478226
rect 332938 478170 333008 478226
rect 332688 478102 333008 478170
rect 332688 478046 332758 478102
rect 332814 478046 332882 478102
rect 332938 478046 333008 478102
rect 332688 477978 333008 478046
rect 332688 477922 332758 477978
rect 332814 477922 332882 477978
rect 332938 477922 333008 477978
rect 332688 477888 333008 477922
rect 363408 478350 363728 478384
rect 363408 478294 363478 478350
rect 363534 478294 363602 478350
rect 363658 478294 363728 478350
rect 363408 478226 363728 478294
rect 363408 478170 363478 478226
rect 363534 478170 363602 478226
rect 363658 478170 363728 478226
rect 363408 478102 363728 478170
rect 363408 478046 363478 478102
rect 363534 478046 363602 478102
rect 363658 478046 363728 478102
rect 363408 477978 363728 478046
rect 363408 477922 363478 477978
rect 363534 477922 363602 477978
rect 363658 477922 363728 477978
rect 363408 477888 363728 477922
rect 394128 478350 394448 478384
rect 394128 478294 394198 478350
rect 394254 478294 394322 478350
rect 394378 478294 394448 478350
rect 394128 478226 394448 478294
rect 394128 478170 394198 478226
rect 394254 478170 394322 478226
rect 394378 478170 394448 478226
rect 394128 478102 394448 478170
rect 394128 478046 394198 478102
rect 394254 478046 394322 478102
rect 394378 478046 394448 478102
rect 394128 477978 394448 478046
rect 394128 477922 394198 477978
rect 394254 477922 394322 477978
rect 394378 477922 394448 477978
rect 394128 477888 394448 477922
rect 424848 478350 425168 478384
rect 424848 478294 424918 478350
rect 424974 478294 425042 478350
rect 425098 478294 425168 478350
rect 424848 478226 425168 478294
rect 424848 478170 424918 478226
rect 424974 478170 425042 478226
rect 425098 478170 425168 478226
rect 424848 478102 425168 478170
rect 424848 478046 424918 478102
rect 424974 478046 425042 478102
rect 425098 478046 425168 478102
rect 424848 477978 425168 478046
rect 424848 477922 424918 477978
rect 424974 477922 425042 477978
rect 425098 477922 425168 477978
rect 424848 477888 425168 477922
rect 455568 478350 455888 478384
rect 455568 478294 455638 478350
rect 455694 478294 455762 478350
rect 455818 478294 455888 478350
rect 455568 478226 455888 478294
rect 455568 478170 455638 478226
rect 455694 478170 455762 478226
rect 455818 478170 455888 478226
rect 455568 478102 455888 478170
rect 455568 478046 455638 478102
rect 455694 478046 455762 478102
rect 455818 478046 455888 478102
rect 455568 477978 455888 478046
rect 455568 477922 455638 477978
rect 455694 477922 455762 477978
rect 455818 477922 455888 477978
rect 455568 477888 455888 477922
rect 486288 478350 486608 478384
rect 486288 478294 486358 478350
rect 486414 478294 486482 478350
rect 486538 478294 486608 478350
rect 486288 478226 486608 478294
rect 486288 478170 486358 478226
rect 486414 478170 486482 478226
rect 486538 478170 486608 478226
rect 486288 478102 486608 478170
rect 486288 478046 486358 478102
rect 486414 478046 486482 478102
rect 486538 478046 486608 478102
rect 486288 477978 486608 478046
rect 486288 477922 486358 477978
rect 486414 477922 486482 477978
rect 486538 477922 486608 477978
rect 486288 477888 486608 477922
rect 194448 472350 194768 472384
rect 194448 472294 194518 472350
rect 194574 472294 194642 472350
rect 194698 472294 194768 472350
rect 194448 472226 194768 472294
rect 194448 472170 194518 472226
rect 194574 472170 194642 472226
rect 194698 472170 194768 472226
rect 194448 472102 194768 472170
rect 194448 472046 194518 472102
rect 194574 472046 194642 472102
rect 194698 472046 194768 472102
rect 194448 471978 194768 472046
rect 194448 471922 194518 471978
rect 194574 471922 194642 471978
rect 194698 471922 194768 471978
rect 194448 471888 194768 471922
rect 225168 472350 225488 472384
rect 225168 472294 225238 472350
rect 225294 472294 225362 472350
rect 225418 472294 225488 472350
rect 225168 472226 225488 472294
rect 225168 472170 225238 472226
rect 225294 472170 225362 472226
rect 225418 472170 225488 472226
rect 225168 472102 225488 472170
rect 225168 472046 225238 472102
rect 225294 472046 225362 472102
rect 225418 472046 225488 472102
rect 225168 471978 225488 472046
rect 225168 471922 225238 471978
rect 225294 471922 225362 471978
rect 225418 471922 225488 471978
rect 225168 471888 225488 471922
rect 255888 472350 256208 472384
rect 255888 472294 255958 472350
rect 256014 472294 256082 472350
rect 256138 472294 256208 472350
rect 255888 472226 256208 472294
rect 255888 472170 255958 472226
rect 256014 472170 256082 472226
rect 256138 472170 256208 472226
rect 255888 472102 256208 472170
rect 255888 472046 255958 472102
rect 256014 472046 256082 472102
rect 256138 472046 256208 472102
rect 255888 471978 256208 472046
rect 255888 471922 255958 471978
rect 256014 471922 256082 471978
rect 256138 471922 256208 471978
rect 255888 471888 256208 471922
rect 286608 472350 286928 472384
rect 286608 472294 286678 472350
rect 286734 472294 286802 472350
rect 286858 472294 286928 472350
rect 286608 472226 286928 472294
rect 286608 472170 286678 472226
rect 286734 472170 286802 472226
rect 286858 472170 286928 472226
rect 286608 472102 286928 472170
rect 286608 472046 286678 472102
rect 286734 472046 286802 472102
rect 286858 472046 286928 472102
rect 286608 471978 286928 472046
rect 286608 471922 286678 471978
rect 286734 471922 286802 471978
rect 286858 471922 286928 471978
rect 286608 471888 286928 471922
rect 317328 472350 317648 472384
rect 317328 472294 317398 472350
rect 317454 472294 317522 472350
rect 317578 472294 317648 472350
rect 317328 472226 317648 472294
rect 317328 472170 317398 472226
rect 317454 472170 317522 472226
rect 317578 472170 317648 472226
rect 317328 472102 317648 472170
rect 317328 472046 317398 472102
rect 317454 472046 317522 472102
rect 317578 472046 317648 472102
rect 317328 471978 317648 472046
rect 317328 471922 317398 471978
rect 317454 471922 317522 471978
rect 317578 471922 317648 471978
rect 317328 471888 317648 471922
rect 348048 472350 348368 472384
rect 348048 472294 348118 472350
rect 348174 472294 348242 472350
rect 348298 472294 348368 472350
rect 348048 472226 348368 472294
rect 348048 472170 348118 472226
rect 348174 472170 348242 472226
rect 348298 472170 348368 472226
rect 348048 472102 348368 472170
rect 348048 472046 348118 472102
rect 348174 472046 348242 472102
rect 348298 472046 348368 472102
rect 348048 471978 348368 472046
rect 348048 471922 348118 471978
rect 348174 471922 348242 471978
rect 348298 471922 348368 471978
rect 348048 471888 348368 471922
rect 378768 472350 379088 472384
rect 378768 472294 378838 472350
rect 378894 472294 378962 472350
rect 379018 472294 379088 472350
rect 378768 472226 379088 472294
rect 378768 472170 378838 472226
rect 378894 472170 378962 472226
rect 379018 472170 379088 472226
rect 378768 472102 379088 472170
rect 378768 472046 378838 472102
rect 378894 472046 378962 472102
rect 379018 472046 379088 472102
rect 378768 471978 379088 472046
rect 378768 471922 378838 471978
rect 378894 471922 378962 471978
rect 379018 471922 379088 471978
rect 378768 471888 379088 471922
rect 409488 472350 409808 472384
rect 409488 472294 409558 472350
rect 409614 472294 409682 472350
rect 409738 472294 409808 472350
rect 409488 472226 409808 472294
rect 409488 472170 409558 472226
rect 409614 472170 409682 472226
rect 409738 472170 409808 472226
rect 409488 472102 409808 472170
rect 409488 472046 409558 472102
rect 409614 472046 409682 472102
rect 409738 472046 409808 472102
rect 409488 471978 409808 472046
rect 409488 471922 409558 471978
rect 409614 471922 409682 471978
rect 409738 471922 409808 471978
rect 409488 471888 409808 471922
rect 440208 472350 440528 472384
rect 440208 472294 440278 472350
rect 440334 472294 440402 472350
rect 440458 472294 440528 472350
rect 440208 472226 440528 472294
rect 440208 472170 440278 472226
rect 440334 472170 440402 472226
rect 440458 472170 440528 472226
rect 440208 472102 440528 472170
rect 440208 472046 440278 472102
rect 440334 472046 440402 472102
rect 440458 472046 440528 472102
rect 440208 471978 440528 472046
rect 440208 471922 440278 471978
rect 440334 471922 440402 471978
rect 440458 471922 440528 471978
rect 440208 471888 440528 471922
rect 470928 472350 471248 472384
rect 470928 472294 470998 472350
rect 471054 472294 471122 472350
rect 471178 472294 471248 472350
rect 470928 472226 471248 472294
rect 470928 472170 470998 472226
rect 471054 472170 471122 472226
rect 471178 472170 471248 472226
rect 470928 472102 471248 472170
rect 470928 472046 470998 472102
rect 471054 472046 471122 472102
rect 471178 472046 471248 472102
rect 470928 471978 471248 472046
rect 470928 471922 470998 471978
rect 471054 471922 471122 471978
rect 471178 471922 471248 471978
rect 470928 471888 471248 471922
rect 501648 472350 501968 472384
rect 501648 472294 501718 472350
rect 501774 472294 501842 472350
rect 501898 472294 501968 472350
rect 501648 472226 501968 472294
rect 501648 472170 501718 472226
rect 501774 472170 501842 472226
rect 501898 472170 501968 472226
rect 501648 472102 501968 472170
rect 501648 472046 501718 472102
rect 501774 472046 501842 472102
rect 501898 472046 501968 472102
rect 501648 471978 501968 472046
rect 501648 471922 501718 471978
rect 501774 471922 501842 471978
rect 501898 471922 501968 471978
rect 501648 471888 501968 471922
rect 209808 460350 210128 460384
rect 209808 460294 209878 460350
rect 209934 460294 210002 460350
rect 210058 460294 210128 460350
rect 209808 460226 210128 460294
rect 209808 460170 209878 460226
rect 209934 460170 210002 460226
rect 210058 460170 210128 460226
rect 209808 460102 210128 460170
rect 209808 460046 209878 460102
rect 209934 460046 210002 460102
rect 210058 460046 210128 460102
rect 209808 459978 210128 460046
rect 209808 459922 209878 459978
rect 209934 459922 210002 459978
rect 210058 459922 210128 459978
rect 209808 459888 210128 459922
rect 240528 460350 240848 460384
rect 240528 460294 240598 460350
rect 240654 460294 240722 460350
rect 240778 460294 240848 460350
rect 240528 460226 240848 460294
rect 240528 460170 240598 460226
rect 240654 460170 240722 460226
rect 240778 460170 240848 460226
rect 240528 460102 240848 460170
rect 240528 460046 240598 460102
rect 240654 460046 240722 460102
rect 240778 460046 240848 460102
rect 240528 459978 240848 460046
rect 240528 459922 240598 459978
rect 240654 459922 240722 459978
rect 240778 459922 240848 459978
rect 240528 459888 240848 459922
rect 271248 460350 271568 460384
rect 271248 460294 271318 460350
rect 271374 460294 271442 460350
rect 271498 460294 271568 460350
rect 271248 460226 271568 460294
rect 271248 460170 271318 460226
rect 271374 460170 271442 460226
rect 271498 460170 271568 460226
rect 271248 460102 271568 460170
rect 271248 460046 271318 460102
rect 271374 460046 271442 460102
rect 271498 460046 271568 460102
rect 271248 459978 271568 460046
rect 271248 459922 271318 459978
rect 271374 459922 271442 459978
rect 271498 459922 271568 459978
rect 271248 459888 271568 459922
rect 301968 460350 302288 460384
rect 301968 460294 302038 460350
rect 302094 460294 302162 460350
rect 302218 460294 302288 460350
rect 301968 460226 302288 460294
rect 301968 460170 302038 460226
rect 302094 460170 302162 460226
rect 302218 460170 302288 460226
rect 301968 460102 302288 460170
rect 301968 460046 302038 460102
rect 302094 460046 302162 460102
rect 302218 460046 302288 460102
rect 301968 459978 302288 460046
rect 301968 459922 302038 459978
rect 302094 459922 302162 459978
rect 302218 459922 302288 459978
rect 301968 459888 302288 459922
rect 332688 460350 333008 460384
rect 332688 460294 332758 460350
rect 332814 460294 332882 460350
rect 332938 460294 333008 460350
rect 332688 460226 333008 460294
rect 332688 460170 332758 460226
rect 332814 460170 332882 460226
rect 332938 460170 333008 460226
rect 332688 460102 333008 460170
rect 332688 460046 332758 460102
rect 332814 460046 332882 460102
rect 332938 460046 333008 460102
rect 332688 459978 333008 460046
rect 332688 459922 332758 459978
rect 332814 459922 332882 459978
rect 332938 459922 333008 459978
rect 332688 459888 333008 459922
rect 363408 460350 363728 460384
rect 363408 460294 363478 460350
rect 363534 460294 363602 460350
rect 363658 460294 363728 460350
rect 363408 460226 363728 460294
rect 363408 460170 363478 460226
rect 363534 460170 363602 460226
rect 363658 460170 363728 460226
rect 363408 460102 363728 460170
rect 363408 460046 363478 460102
rect 363534 460046 363602 460102
rect 363658 460046 363728 460102
rect 363408 459978 363728 460046
rect 363408 459922 363478 459978
rect 363534 459922 363602 459978
rect 363658 459922 363728 459978
rect 363408 459888 363728 459922
rect 394128 460350 394448 460384
rect 394128 460294 394198 460350
rect 394254 460294 394322 460350
rect 394378 460294 394448 460350
rect 394128 460226 394448 460294
rect 394128 460170 394198 460226
rect 394254 460170 394322 460226
rect 394378 460170 394448 460226
rect 394128 460102 394448 460170
rect 394128 460046 394198 460102
rect 394254 460046 394322 460102
rect 394378 460046 394448 460102
rect 394128 459978 394448 460046
rect 394128 459922 394198 459978
rect 394254 459922 394322 459978
rect 394378 459922 394448 459978
rect 394128 459888 394448 459922
rect 424848 460350 425168 460384
rect 424848 460294 424918 460350
rect 424974 460294 425042 460350
rect 425098 460294 425168 460350
rect 424848 460226 425168 460294
rect 424848 460170 424918 460226
rect 424974 460170 425042 460226
rect 425098 460170 425168 460226
rect 424848 460102 425168 460170
rect 424848 460046 424918 460102
rect 424974 460046 425042 460102
rect 425098 460046 425168 460102
rect 424848 459978 425168 460046
rect 424848 459922 424918 459978
rect 424974 459922 425042 459978
rect 425098 459922 425168 459978
rect 424848 459888 425168 459922
rect 455568 460350 455888 460384
rect 455568 460294 455638 460350
rect 455694 460294 455762 460350
rect 455818 460294 455888 460350
rect 455568 460226 455888 460294
rect 455568 460170 455638 460226
rect 455694 460170 455762 460226
rect 455818 460170 455888 460226
rect 455568 460102 455888 460170
rect 455568 460046 455638 460102
rect 455694 460046 455762 460102
rect 455818 460046 455888 460102
rect 455568 459978 455888 460046
rect 455568 459922 455638 459978
rect 455694 459922 455762 459978
rect 455818 459922 455888 459978
rect 455568 459888 455888 459922
rect 486288 460350 486608 460384
rect 486288 460294 486358 460350
rect 486414 460294 486482 460350
rect 486538 460294 486608 460350
rect 486288 460226 486608 460294
rect 486288 460170 486358 460226
rect 486414 460170 486482 460226
rect 486538 460170 486608 460226
rect 486288 460102 486608 460170
rect 486288 460046 486358 460102
rect 486414 460046 486482 460102
rect 486538 460046 486608 460102
rect 486288 459978 486608 460046
rect 486288 459922 486358 459978
rect 486414 459922 486482 459978
rect 486538 459922 486608 459978
rect 486288 459888 486608 459922
rect 194448 454350 194768 454384
rect 194448 454294 194518 454350
rect 194574 454294 194642 454350
rect 194698 454294 194768 454350
rect 194448 454226 194768 454294
rect 194448 454170 194518 454226
rect 194574 454170 194642 454226
rect 194698 454170 194768 454226
rect 194448 454102 194768 454170
rect 194448 454046 194518 454102
rect 194574 454046 194642 454102
rect 194698 454046 194768 454102
rect 194448 453978 194768 454046
rect 194448 453922 194518 453978
rect 194574 453922 194642 453978
rect 194698 453922 194768 453978
rect 194448 453888 194768 453922
rect 225168 454350 225488 454384
rect 225168 454294 225238 454350
rect 225294 454294 225362 454350
rect 225418 454294 225488 454350
rect 225168 454226 225488 454294
rect 225168 454170 225238 454226
rect 225294 454170 225362 454226
rect 225418 454170 225488 454226
rect 225168 454102 225488 454170
rect 225168 454046 225238 454102
rect 225294 454046 225362 454102
rect 225418 454046 225488 454102
rect 225168 453978 225488 454046
rect 225168 453922 225238 453978
rect 225294 453922 225362 453978
rect 225418 453922 225488 453978
rect 225168 453888 225488 453922
rect 255888 454350 256208 454384
rect 255888 454294 255958 454350
rect 256014 454294 256082 454350
rect 256138 454294 256208 454350
rect 255888 454226 256208 454294
rect 255888 454170 255958 454226
rect 256014 454170 256082 454226
rect 256138 454170 256208 454226
rect 255888 454102 256208 454170
rect 255888 454046 255958 454102
rect 256014 454046 256082 454102
rect 256138 454046 256208 454102
rect 255888 453978 256208 454046
rect 255888 453922 255958 453978
rect 256014 453922 256082 453978
rect 256138 453922 256208 453978
rect 255888 453888 256208 453922
rect 286608 454350 286928 454384
rect 286608 454294 286678 454350
rect 286734 454294 286802 454350
rect 286858 454294 286928 454350
rect 286608 454226 286928 454294
rect 286608 454170 286678 454226
rect 286734 454170 286802 454226
rect 286858 454170 286928 454226
rect 286608 454102 286928 454170
rect 286608 454046 286678 454102
rect 286734 454046 286802 454102
rect 286858 454046 286928 454102
rect 286608 453978 286928 454046
rect 286608 453922 286678 453978
rect 286734 453922 286802 453978
rect 286858 453922 286928 453978
rect 286608 453888 286928 453922
rect 317328 454350 317648 454384
rect 317328 454294 317398 454350
rect 317454 454294 317522 454350
rect 317578 454294 317648 454350
rect 317328 454226 317648 454294
rect 317328 454170 317398 454226
rect 317454 454170 317522 454226
rect 317578 454170 317648 454226
rect 317328 454102 317648 454170
rect 317328 454046 317398 454102
rect 317454 454046 317522 454102
rect 317578 454046 317648 454102
rect 317328 453978 317648 454046
rect 317328 453922 317398 453978
rect 317454 453922 317522 453978
rect 317578 453922 317648 453978
rect 317328 453888 317648 453922
rect 348048 454350 348368 454384
rect 348048 454294 348118 454350
rect 348174 454294 348242 454350
rect 348298 454294 348368 454350
rect 348048 454226 348368 454294
rect 348048 454170 348118 454226
rect 348174 454170 348242 454226
rect 348298 454170 348368 454226
rect 348048 454102 348368 454170
rect 348048 454046 348118 454102
rect 348174 454046 348242 454102
rect 348298 454046 348368 454102
rect 348048 453978 348368 454046
rect 348048 453922 348118 453978
rect 348174 453922 348242 453978
rect 348298 453922 348368 453978
rect 348048 453888 348368 453922
rect 378768 454350 379088 454384
rect 378768 454294 378838 454350
rect 378894 454294 378962 454350
rect 379018 454294 379088 454350
rect 378768 454226 379088 454294
rect 378768 454170 378838 454226
rect 378894 454170 378962 454226
rect 379018 454170 379088 454226
rect 378768 454102 379088 454170
rect 378768 454046 378838 454102
rect 378894 454046 378962 454102
rect 379018 454046 379088 454102
rect 378768 453978 379088 454046
rect 378768 453922 378838 453978
rect 378894 453922 378962 453978
rect 379018 453922 379088 453978
rect 378768 453888 379088 453922
rect 409488 454350 409808 454384
rect 409488 454294 409558 454350
rect 409614 454294 409682 454350
rect 409738 454294 409808 454350
rect 409488 454226 409808 454294
rect 409488 454170 409558 454226
rect 409614 454170 409682 454226
rect 409738 454170 409808 454226
rect 409488 454102 409808 454170
rect 409488 454046 409558 454102
rect 409614 454046 409682 454102
rect 409738 454046 409808 454102
rect 409488 453978 409808 454046
rect 409488 453922 409558 453978
rect 409614 453922 409682 453978
rect 409738 453922 409808 453978
rect 409488 453888 409808 453922
rect 440208 454350 440528 454384
rect 440208 454294 440278 454350
rect 440334 454294 440402 454350
rect 440458 454294 440528 454350
rect 440208 454226 440528 454294
rect 440208 454170 440278 454226
rect 440334 454170 440402 454226
rect 440458 454170 440528 454226
rect 440208 454102 440528 454170
rect 440208 454046 440278 454102
rect 440334 454046 440402 454102
rect 440458 454046 440528 454102
rect 440208 453978 440528 454046
rect 440208 453922 440278 453978
rect 440334 453922 440402 453978
rect 440458 453922 440528 453978
rect 440208 453888 440528 453922
rect 470928 454350 471248 454384
rect 470928 454294 470998 454350
rect 471054 454294 471122 454350
rect 471178 454294 471248 454350
rect 470928 454226 471248 454294
rect 470928 454170 470998 454226
rect 471054 454170 471122 454226
rect 471178 454170 471248 454226
rect 470928 454102 471248 454170
rect 470928 454046 470998 454102
rect 471054 454046 471122 454102
rect 471178 454046 471248 454102
rect 470928 453978 471248 454046
rect 470928 453922 470998 453978
rect 471054 453922 471122 453978
rect 471178 453922 471248 453978
rect 470928 453888 471248 453922
rect 501648 454350 501968 454384
rect 501648 454294 501718 454350
rect 501774 454294 501842 454350
rect 501898 454294 501968 454350
rect 501648 454226 501968 454294
rect 501648 454170 501718 454226
rect 501774 454170 501842 454226
rect 501898 454170 501968 454226
rect 501648 454102 501968 454170
rect 501648 454046 501718 454102
rect 501774 454046 501842 454102
rect 501898 454046 501968 454102
rect 501648 453978 501968 454046
rect 501648 453922 501718 453978
rect 501774 453922 501842 453978
rect 501898 453922 501968 453978
rect 501648 453888 501968 453922
rect 209808 442350 210128 442384
rect 209808 442294 209878 442350
rect 209934 442294 210002 442350
rect 210058 442294 210128 442350
rect 209808 442226 210128 442294
rect 209808 442170 209878 442226
rect 209934 442170 210002 442226
rect 210058 442170 210128 442226
rect 209808 442102 210128 442170
rect 209808 442046 209878 442102
rect 209934 442046 210002 442102
rect 210058 442046 210128 442102
rect 209808 441978 210128 442046
rect 209808 441922 209878 441978
rect 209934 441922 210002 441978
rect 210058 441922 210128 441978
rect 209808 441888 210128 441922
rect 240528 442350 240848 442384
rect 240528 442294 240598 442350
rect 240654 442294 240722 442350
rect 240778 442294 240848 442350
rect 240528 442226 240848 442294
rect 240528 442170 240598 442226
rect 240654 442170 240722 442226
rect 240778 442170 240848 442226
rect 240528 442102 240848 442170
rect 240528 442046 240598 442102
rect 240654 442046 240722 442102
rect 240778 442046 240848 442102
rect 240528 441978 240848 442046
rect 240528 441922 240598 441978
rect 240654 441922 240722 441978
rect 240778 441922 240848 441978
rect 240528 441888 240848 441922
rect 271248 442350 271568 442384
rect 271248 442294 271318 442350
rect 271374 442294 271442 442350
rect 271498 442294 271568 442350
rect 271248 442226 271568 442294
rect 271248 442170 271318 442226
rect 271374 442170 271442 442226
rect 271498 442170 271568 442226
rect 271248 442102 271568 442170
rect 271248 442046 271318 442102
rect 271374 442046 271442 442102
rect 271498 442046 271568 442102
rect 271248 441978 271568 442046
rect 271248 441922 271318 441978
rect 271374 441922 271442 441978
rect 271498 441922 271568 441978
rect 271248 441888 271568 441922
rect 301968 442350 302288 442384
rect 301968 442294 302038 442350
rect 302094 442294 302162 442350
rect 302218 442294 302288 442350
rect 301968 442226 302288 442294
rect 301968 442170 302038 442226
rect 302094 442170 302162 442226
rect 302218 442170 302288 442226
rect 301968 442102 302288 442170
rect 301968 442046 302038 442102
rect 302094 442046 302162 442102
rect 302218 442046 302288 442102
rect 301968 441978 302288 442046
rect 301968 441922 302038 441978
rect 302094 441922 302162 441978
rect 302218 441922 302288 441978
rect 301968 441888 302288 441922
rect 332688 442350 333008 442384
rect 332688 442294 332758 442350
rect 332814 442294 332882 442350
rect 332938 442294 333008 442350
rect 332688 442226 333008 442294
rect 332688 442170 332758 442226
rect 332814 442170 332882 442226
rect 332938 442170 333008 442226
rect 332688 442102 333008 442170
rect 332688 442046 332758 442102
rect 332814 442046 332882 442102
rect 332938 442046 333008 442102
rect 332688 441978 333008 442046
rect 332688 441922 332758 441978
rect 332814 441922 332882 441978
rect 332938 441922 333008 441978
rect 332688 441888 333008 441922
rect 363408 442350 363728 442384
rect 363408 442294 363478 442350
rect 363534 442294 363602 442350
rect 363658 442294 363728 442350
rect 363408 442226 363728 442294
rect 363408 442170 363478 442226
rect 363534 442170 363602 442226
rect 363658 442170 363728 442226
rect 363408 442102 363728 442170
rect 363408 442046 363478 442102
rect 363534 442046 363602 442102
rect 363658 442046 363728 442102
rect 363408 441978 363728 442046
rect 363408 441922 363478 441978
rect 363534 441922 363602 441978
rect 363658 441922 363728 441978
rect 363408 441888 363728 441922
rect 394128 442350 394448 442384
rect 394128 442294 394198 442350
rect 394254 442294 394322 442350
rect 394378 442294 394448 442350
rect 394128 442226 394448 442294
rect 394128 442170 394198 442226
rect 394254 442170 394322 442226
rect 394378 442170 394448 442226
rect 394128 442102 394448 442170
rect 394128 442046 394198 442102
rect 394254 442046 394322 442102
rect 394378 442046 394448 442102
rect 394128 441978 394448 442046
rect 394128 441922 394198 441978
rect 394254 441922 394322 441978
rect 394378 441922 394448 441978
rect 394128 441888 394448 441922
rect 424848 442350 425168 442384
rect 424848 442294 424918 442350
rect 424974 442294 425042 442350
rect 425098 442294 425168 442350
rect 424848 442226 425168 442294
rect 424848 442170 424918 442226
rect 424974 442170 425042 442226
rect 425098 442170 425168 442226
rect 424848 442102 425168 442170
rect 424848 442046 424918 442102
rect 424974 442046 425042 442102
rect 425098 442046 425168 442102
rect 424848 441978 425168 442046
rect 424848 441922 424918 441978
rect 424974 441922 425042 441978
rect 425098 441922 425168 441978
rect 424848 441888 425168 441922
rect 455568 442350 455888 442384
rect 455568 442294 455638 442350
rect 455694 442294 455762 442350
rect 455818 442294 455888 442350
rect 455568 442226 455888 442294
rect 455568 442170 455638 442226
rect 455694 442170 455762 442226
rect 455818 442170 455888 442226
rect 455568 442102 455888 442170
rect 455568 442046 455638 442102
rect 455694 442046 455762 442102
rect 455818 442046 455888 442102
rect 455568 441978 455888 442046
rect 455568 441922 455638 441978
rect 455694 441922 455762 441978
rect 455818 441922 455888 441978
rect 455568 441888 455888 441922
rect 486288 442350 486608 442384
rect 486288 442294 486358 442350
rect 486414 442294 486482 442350
rect 486538 442294 486608 442350
rect 486288 442226 486608 442294
rect 486288 442170 486358 442226
rect 486414 442170 486482 442226
rect 486538 442170 486608 442226
rect 486288 442102 486608 442170
rect 486288 442046 486358 442102
rect 486414 442046 486482 442102
rect 486538 442046 486608 442102
rect 486288 441978 486608 442046
rect 486288 441922 486358 441978
rect 486414 441922 486482 441978
rect 486538 441922 486608 441978
rect 486288 441888 486608 441922
rect 194448 436350 194768 436384
rect 194448 436294 194518 436350
rect 194574 436294 194642 436350
rect 194698 436294 194768 436350
rect 194448 436226 194768 436294
rect 194448 436170 194518 436226
rect 194574 436170 194642 436226
rect 194698 436170 194768 436226
rect 194448 436102 194768 436170
rect 194448 436046 194518 436102
rect 194574 436046 194642 436102
rect 194698 436046 194768 436102
rect 194448 435978 194768 436046
rect 194448 435922 194518 435978
rect 194574 435922 194642 435978
rect 194698 435922 194768 435978
rect 194448 435888 194768 435922
rect 225168 436350 225488 436384
rect 225168 436294 225238 436350
rect 225294 436294 225362 436350
rect 225418 436294 225488 436350
rect 225168 436226 225488 436294
rect 225168 436170 225238 436226
rect 225294 436170 225362 436226
rect 225418 436170 225488 436226
rect 225168 436102 225488 436170
rect 225168 436046 225238 436102
rect 225294 436046 225362 436102
rect 225418 436046 225488 436102
rect 225168 435978 225488 436046
rect 225168 435922 225238 435978
rect 225294 435922 225362 435978
rect 225418 435922 225488 435978
rect 225168 435888 225488 435922
rect 255888 436350 256208 436384
rect 255888 436294 255958 436350
rect 256014 436294 256082 436350
rect 256138 436294 256208 436350
rect 255888 436226 256208 436294
rect 255888 436170 255958 436226
rect 256014 436170 256082 436226
rect 256138 436170 256208 436226
rect 255888 436102 256208 436170
rect 255888 436046 255958 436102
rect 256014 436046 256082 436102
rect 256138 436046 256208 436102
rect 255888 435978 256208 436046
rect 255888 435922 255958 435978
rect 256014 435922 256082 435978
rect 256138 435922 256208 435978
rect 255888 435888 256208 435922
rect 286608 436350 286928 436384
rect 286608 436294 286678 436350
rect 286734 436294 286802 436350
rect 286858 436294 286928 436350
rect 286608 436226 286928 436294
rect 286608 436170 286678 436226
rect 286734 436170 286802 436226
rect 286858 436170 286928 436226
rect 286608 436102 286928 436170
rect 286608 436046 286678 436102
rect 286734 436046 286802 436102
rect 286858 436046 286928 436102
rect 286608 435978 286928 436046
rect 286608 435922 286678 435978
rect 286734 435922 286802 435978
rect 286858 435922 286928 435978
rect 286608 435888 286928 435922
rect 317328 436350 317648 436384
rect 317328 436294 317398 436350
rect 317454 436294 317522 436350
rect 317578 436294 317648 436350
rect 317328 436226 317648 436294
rect 317328 436170 317398 436226
rect 317454 436170 317522 436226
rect 317578 436170 317648 436226
rect 317328 436102 317648 436170
rect 317328 436046 317398 436102
rect 317454 436046 317522 436102
rect 317578 436046 317648 436102
rect 317328 435978 317648 436046
rect 317328 435922 317398 435978
rect 317454 435922 317522 435978
rect 317578 435922 317648 435978
rect 317328 435888 317648 435922
rect 348048 436350 348368 436384
rect 348048 436294 348118 436350
rect 348174 436294 348242 436350
rect 348298 436294 348368 436350
rect 348048 436226 348368 436294
rect 348048 436170 348118 436226
rect 348174 436170 348242 436226
rect 348298 436170 348368 436226
rect 348048 436102 348368 436170
rect 348048 436046 348118 436102
rect 348174 436046 348242 436102
rect 348298 436046 348368 436102
rect 348048 435978 348368 436046
rect 348048 435922 348118 435978
rect 348174 435922 348242 435978
rect 348298 435922 348368 435978
rect 348048 435888 348368 435922
rect 378768 436350 379088 436384
rect 378768 436294 378838 436350
rect 378894 436294 378962 436350
rect 379018 436294 379088 436350
rect 378768 436226 379088 436294
rect 378768 436170 378838 436226
rect 378894 436170 378962 436226
rect 379018 436170 379088 436226
rect 378768 436102 379088 436170
rect 378768 436046 378838 436102
rect 378894 436046 378962 436102
rect 379018 436046 379088 436102
rect 378768 435978 379088 436046
rect 378768 435922 378838 435978
rect 378894 435922 378962 435978
rect 379018 435922 379088 435978
rect 378768 435888 379088 435922
rect 409488 436350 409808 436384
rect 409488 436294 409558 436350
rect 409614 436294 409682 436350
rect 409738 436294 409808 436350
rect 409488 436226 409808 436294
rect 409488 436170 409558 436226
rect 409614 436170 409682 436226
rect 409738 436170 409808 436226
rect 409488 436102 409808 436170
rect 409488 436046 409558 436102
rect 409614 436046 409682 436102
rect 409738 436046 409808 436102
rect 409488 435978 409808 436046
rect 409488 435922 409558 435978
rect 409614 435922 409682 435978
rect 409738 435922 409808 435978
rect 409488 435888 409808 435922
rect 440208 436350 440528 436384
rect 440208 436294 440278 436350
rect 440334 436294 440402 436350
rect 440458 436294 440528 436350
rect 440208 436226 440528 436294
rect 440208 436170 440278 436226
rect 440334 436170 440402 436226
rect 440458 436170 440528 436226
rect 440208 436102 440528 436170
rect 440208 436046 440278 436102
rect 440334 436046 440402 436102
rect 440458 436046 440528 436102
rect 440208 435978 440528 436046
rect 440208 435922 440278 435978
rect 440334 435922 440402 435978
rect 440458 435922 440528 435978
rect 440208 435888 440528 435922
rect 470928 436350 471248 436384
rect 470928 436294 470998 436350
rect 471054 436294 471122 436350
rect 471178 436294 471248 436350
rect 470928 436226 471248 436294
rect 470928 436170 470998 436226
rect 471054 436170 471122 436226
rect 471178 436170 471248 436226
rect 470928 436102 471248 436170
rect 470928 436046 470998 436102
rect 471054 436046 471122 436102
rect 471178 436046 471248 436102
rect 470928 435978 471248 436046
rect 470928 435922 470998 435978
rect 471054 435922 471122 435978
rect 471178 435922 471248 435978
rect 470928 435888 471248 435922
rect 501648 436350 501968 436384
rect 501648 436294 501718 436350
rect 501774 436294 501842 436350
rect 501898 436294 501968 436350
rect 501648 436226 501968 436294
rect 501648 436170 501718 436226
rect 501774 436170 501842 436226
rect 501898 436170 501968 436226
rect 501648 436102 501968 436170
rect 501648 436046 501718 436102
rect 501774 436046 501842 436102
rect 501898 436046 501968 436102
rect 501648 435978 501968 436046
rect 501648 435922 501718 435978
rect 501774 435922 501842 435978
rect 501898 435922 501968 435978
rect 501648 435888 501968 435922
rect 209808 424350 210128 424384
rect 209808 424294 209878 424350
rect 209934 424294 210002 424350
rect 210058 424294 210128 424350
rect 209808 424226 210128 424294
rect 209808 424170 209878 424226
rect 209934 424170 210002 424226
rect 210058 424170 210128 424226
rect 209808 424102 210128 424170
rect 209808 424046 209878 424102
rect 209934 424046 210002 424102
rect 210058 424046 210128 424102
rect 209808 423978 210128 424046
rect 209808 423922 209878 423978
rect 209934 423922 210002 423978
rect 210058 423922 210128 423978
rect 209808 423888 210128 423922
rect 240528 424350 240848 424384
rect 240528 424294 240598 424350
rect 240654 424294 240722 424350
rect 240778 424294 240848 424350
rect 240528 424226 240848 424294
rect 240528 424170 240598 424226
rect 240654 424170 240722 424226
rect 240778 424170 240848 424226
rect 240528 424102 240848 424170
rect 240528 424046 240598 424102
rect 240654 424046 240722 424102
rect 240778 424046 240848 424102
rect 240528 423978 240848 424046
rect 240528 423922 240598 423978
rect 240654 423922 240722 423978
rect 240778 423922 240848 423978
rect 240528 423888 240848 423922
rect 271248 424350 271568 424384
rect 271248 424294 271318 424350
rect 271374 424294 271442 424350
rect 271498 424294 271568 424350
rect 271248 424226 271568 424294
rect 271248 424170 271318 424226
rect 271374 424170 271442 424226
rect 271498 424170 271568 424226
rect 271248 424102 271568 424170
rect 271248 424046 271318 424102
rect 271374 424046 271442 424102
rect 271498 424046 271568 424102
rect 271248 423978 271568 424046
rect 271248 423922 271318 423978
rect 271374 423922 271442 423978
rect 271498 423922 271568 423978
rect 271248 423888 271568 423922
rect 301968 424350 302288 424384
rect 301968 424294 302038 424350
rect 302094 424294 302162 424350
rect 302218 424294 302288 424350
rect 301968 424226 302288 424294
rect 301968 424170 302038 424226
rect 302094 424170 302162 424226
rect 302218 424170 302288 424226
rect 301968 424102 302288 424170
rect 301968 424046 302038 424102
rect 302094 424046 302162 424102
rect 302218 424046 302288 424102
rect 301968 423978 302288 424046
rect 301968 423922 302038 423978
rect 302094 423922 302162 423978
rect 302218 423922 302288 423978
rect 301968 423888 302288 423922
rect 332688 424350 333008 424384
rect 332688 424294 332758 424350
rect 332814 424294 332882 424350
rect 332938 424294 333008 424350
rect 332688 424226 333008 424294
rect 332688 424170 332758 424226
rect 332814 424170 332882 424226
rect 332938 424170 333008 424226
rect 332688 424102 333008 424170
rect 332688 424046 332758 424102
rect 332814 424046 332882 424102
rect 332938 424046 333008 424102
rect 332688 423978 333008 424046
rect 332688 423922 332758 423978
rect 332814 423922 332882 423978
rect 332938 423922 333008 423978
rect 332688 423888 333008 423922
rect 363408 424350 363728 424384
rect 363408 424294 363478 424350
rect 363534 424294 363602 424350
rect 363658 424294 363728 424350
rect 363408 424226 363728 424294
rect 363408 424170 363478 424226
rect 363534 424170 363602 424226
rect 363658 424170 363728 424226
rect 363408 424102 363728 424170
rect 363408 424046 363478 424102
rect 363534 424046 363602 424102
rect 363658 424046 363728 424102
rect 363408 423978 363728 424046
rect 363408 423922 363478 423978
rect 363534 423922 363602 423978
rect 363658 423922 363728 423978
rect 363408 423888 363728 423922
rect 394128 424350 394448 424384
rect 394128 424294 394198 424350
rect 394254 424294 394322 424350
rect 394378 424294 394448 424350
rect 394128 424226 394448 424294
rect 394128 424170 394198 424226
rect 394254 424170 394322 424226
rect 394378 424170 394448 424226
rect 394128 424102 394448 424170
rect 394128 424046 394198 424102
rect 394254 424046 394322 424102
rect 394378 424046 394448 424102
rect 394128 423978 394448 424046
rect 394128 423922 394198 423978
rect 394254 423922 394322 423978
rect 394378 423922 394448 423978
rect 394128 423888 394448 423922
rect 424848 424350 425168 424384
rect 424848 424294 424918 424350
rect 424974 424294 425042 424350
rect 425098 424294 425168 424350
rect 424848 424226 425168 424294
rect 424848 424170 424918 424226
rect 424974 424170 425042 424226
rect 425098 424170 425168 424226
rect 424848 424102 425168 424170
rect 424848 424046 424918 424102
rect 424974 424046 425042 424102
rect 425098 424046 425168 424102
rect 424848 423978 425168 424046
rect 424848 423922 424918 423978
rect 424974 423922 425042 423978
rect 425098 423922 425168 423978
rect 424848 423888 425168 423922
rect 455568 424350 455888 424384
rect 455568 424294 455638 424350
rect 455694 424294 455762 424350
rect 455818 424294 455888 424350
rect 455568 424226 455888 424294
rect 455568 424170 455638 424226
rect 455694 424170 455762 424226
rect 455818 424170 455888 424226
rect 455568 424102 455888 424170
rect 455568 424046 455638 424102
rect 455694 424046 455762 424102
rect 455818 424046 455888 424102
rect 455568 423978 455888 424046
rect 455568 423922 455638 423978
rect 455694 423922 455762 423978
rect 455818 423922 455888 423978
rect 455568 423888 455888 423922
rect 486288 424350 486608 424384
rect 486288 424294 486358 424350
rect 486414 424294 486482 424350
rect 486538 424294 486608 424350
rect 486288 424226 486608 424294
rect 486288 424170 486358 424226
rect 486414 424170 486482 424226
rect 486538 424170 486608 424226
rect 486288 424102 486608 424170
rect 486288 424046 486358 424102
rect 486414 424046 486482 424102
rect 486538 424046 486608 424102
rect 486288 423978 486608 424046
rect 486288 423922 486358 423978
rect 486414 423922 486482 423978
rect 486538 423922 486608 423978
rect 486288 423888 486608 423922
rect 194448 418350 194768 418384
rect 194448 418294 194518 418350
rect 194574 418294 194642 418350
rect 194698 418294 194768 418350
rect 194448 418226 194768 418294
rect 194448 418170 194518 418226
rect 194574 418170 194642 418226
rect 194698 418170 194768 418226
rect 194448 418102 194768 418170
rect 194448 418046 194518 418102
rect 194574 418046 194642 418102
rect 194698 418046 194768 418102
rect 194448 417978 194768 418046
rect 194448 417922 194518 417978
rect 194574 417922 194642 417978
rect 194698 417922 194768 417978
rect 194448 417888 194768 417922
rect 225168 418350 225488 418384
rect 225168 418294 225238 418350
rect 225294 418294 225362 418350
rect 225418 418294 225488 418350
rect 225168 418226 225488 418294
rect 225168 418170 225238 418226
rect 225294 418170 225362 418226
rect 225418 418170 225488 418226
rect 225168 418102 225488 418170
rect 225168 418046 225238 418102
rect 225294 418046 225362 418102
rect 225418 418046 225488 418102
rect 225168 417978 225488 418046
rect 225168 417922 225238 417978
rect 225294 417922 225362 417978
rect 225418 417922 225488 417978
rect 225168 417888 225488 417922
rect 255888 418350 256208 418384
rect 255888 418294 255958 418350
rect 256014 418294 256082 418350
rect 256138 418294 256208 418350
rect 255888 418226 256208 418294
rect 255888 418170 255958 418226
rect 256014 418170 256082 418226
rect 256138 418170 256208 418226
rect 255888 418102 256208 418170
rect 255888 418046 255958 418102
rect 256014 418046 256082 418102
rect 256138 418046 256208 418102
rect 255888 417978 256208 418046
rect 255888 417922 255958 417978
rect 256014 417922 256082 417978
rect 256138 417922 256208 417978
rect 255888 417888 256208 417922
rect 286608 418350 286928 418384
rect 286608 418294 286678 418350
rect 286734 418294 286802 418350
rect 286858 418294 286928 418350
rect 286608 418226 286928 418294
rect 286608 418170 286678 418226
rect 286734 418170 286802 418226
rect 286858 418170 286928 418226
rect 286608 418102 286928 418170
rect 286608 418046 286678 418102
rect 286734 418046 286802 418102
rect 286858 418046 286928 418102
rect 286608 417978 286928 418046
rect 286608 417922 286678 417978
rect 286734 417922 286802 417978
rect 286858 417922 286928 417978
rect 286608 417888 286928 417922
rect 317328 418350 317648 418384
rect 317328 418294 317398 418350
rect 317454 418294 317522 418350
rect 317578 418294 317648 418350
rect 317328 418226 317648 418294
rect 317328 418170 317398 418226
rect 317454 418170 317522 418226
rect 317578 418170 317648 418226
rect 317328 418102 317648 418170
rect 317328 418046 317398 418102
rect 317454 418046 317522 418102
rect 317578 418046 317648 418102
rect 317328 417978 317648 418046
rect 317328 417922 317398 417978
rect 317454 417922 317522 417978
rect 317578 417922 317648 417978
rect 317328 417888 317648 417922
rect 348048 418350 348368 418384
rect 348048 418294 348118 418350
rect 348174 418294 348242 418350
rect 348298 418294 348368 418350
rect 348048 418226 348368 418294
rect 348048 418170 348118 418226
rect 348174 418170 348242 418226
rect 348298 418170 348368 418226
rect 348048 418102 348368 418170
rect 348048 418046 348118 418102
rect 348174 418046 348242 418102
rect 348298 418046 348368 418102
rect 348048 417978 348368 418046
rect 348048 417922 348118 417978
rect 348174 417922 348242 417978
rect 348298 417922 348368 417978
rect 348048 417888 348368 417922
rect 378768 418350 379088 418384
rect 378768 418294 378838 418350
rect 378894 418294 378962 418350
rect 379018 418294 379088 418350
rect 378768 418226 379088 418294
rect 378768 418170 378838 418226
rect 378894 418170 378962 418226
rect 379018 418170 379088 418226
rect 378768 418102 379088 418170
rect 378768 418046 378838 418102
rect 378894 418046 378962 418102
rect 379018 418046 379088 418102
rect 378768 417978 379088 418046
rect 378768 417922 378838 417978
rect 378894 417922 378962 417978
rect 379018 417922 379088 417978
rect 378768 417888 379088 417922
rect 409488 418350 409808 418384
rect 409488 418294 409558 418350
rect 409614 418294 409682 418350
rect 409738 418294 409808 418350
rect 409488 418226 409808 418294
rect 409488 418170 409558 418226
rect 409614 418170 409682 418226
rect 409738 418170 409808 418226
rect 409488 418102 409808 418170
rect 409488 418046 409558 418102
rect 409614 418046 409682 418102
rect 409738 418046 409808 418102
rect 409488 417978 409808 418046
rect 409488 417922 409558 417978
rect 409614 417922 409682 417978
rect 409738 417922 409808 417978
rect 409488 417888 409808 417922
rect 440208 418350 440528 418384
rect 440208 418294 440278 418350
rect 440334 418294 440402 418350
rect 440458 418294 440528 418350
rect 440208 418226 440528 418294
rect 440208 418170 440278 418226
rect 440334 418170 440402 418226
rect 440458 418170 440528 418226
rect 440208 418102 440528 418170
rect 440208 418046 440278 418102
rect 440334 418046 440402 418102
rect 440458 418046 440528 418102
rect 440208 417978 440528 418046
rect 440208 417922 440278 417978
rect 440334 417922 440402 417978
rect 440458 417922 440528 417978
rect 440208 417888 440528 417922
rect 470928 418350 471248 418384
rect 470928 418294 470998 418350
rect 471054 418294 471122 418350
rect 471178 418294 471248 418350
rect 470928 418226 471248 418294
rect 470928 418170 470998 418226
rect 471054 418170 471122 418226
rect 471178 418170 471248 418226
rect 470928 418102 471248 418170
rect 470928 418046 470998 418102
rect 471054 418046 471122 418102
rect 471178 418046 471248 418102
rect 470928 417978 471248 418046
rect 470928 417922 470998 417978
rect 471054 417922 471122 417978
rect 471178 417922 471248 417978
rect 470928 417888 471248 417922
rect 501648 418350 501968 418384
rect 501648 418294 501718 418350
rect 501774 418294 501842 418350
rect 501898 418294 501968 418350
rect 501648 418226 501968 418294
rect 501648 418170 501718 418226
rect 501774 418170 501842 418226
rect 501898 418170 501968 418226
rect 501648 418102 501968 418170
rect 501648 418046 501718 418102
rect 501774 418046 501842 418102
rect 501898 418046 501968 418102
rect 501648 417978 501968 418046
rect 501648 417922 501718 417978
rect 501774 417922 501842 417978
rect 501898 417922 501968 417978
rect 501648 417888 501968 417922
rect 357196 411058 357252 411068
rect 334236 410878 334292 410888
rect 324156 410698 324212 410708
rect 194236 405794 194292 405804
rect 209916 404578 209972 404588
rect 208236 404398 208292 404408
rect 206556 404218 206612 404228
rect 193458 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 194078 388350
rect 193458 388226 194078 388294
rect 193458 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 194078 388226
rect 193458 388102 194078 388170
rect 193458 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 194078 388102
rect 193458 387978 194078 388046
rect 193458 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 194078 387978
rect 189738 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 190358 364350
rect 189738 364226 190358 364294
rect 189738 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 190358 364226
rect 189738 364102 190358 364170
rect 189738 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 190358 364102
rect 189738 363978 190358 364046
rect 189738 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 190358 363978
rect 189738 346350 190358 363922
rect 189738 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 190358 346350
rect 189738 346226 190358 346294
rect 189738 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 190358 346226
rect 189738 346102 190358 346170
rect 189738 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 190358 346102
rect 189738 345978 190358 346046
rect 189738 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 190358 345978
rect 189738 328350 190358 345922
rect 189738 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 190358 328350
rect 189738 328226 190358 328294
rect 189738 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 190358 328226
rect 189738 328102 190358 328170
rect 189738 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 190358 328102
rect 189738 327978 190358 328046
rect 189738 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 190358 327978
rect 189738 310350 190358 327922
rect 193458 370350 194078 387922
rect 196476 402058 196532 402068
rect 196476 382004 196532 402002
rect 198156 401878 198212 401888
rect 198044 393238 198100 393248
rect 197484 391798 197540 391808
rect 196476 381938 196532 381948
rect 197372 383796 197428 383806
rect 196364 379652 196420 379662
rect 196140 379428 196196 379438
rect 196140 372988 196196 379372
rect 196364 379428 196420 379596
rect 196364 379362 196420 379372
rect 196140 372932 196532 372988
rect 193458 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 194078 370350
rect 193458 370226 194078 370294
rect 193458 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 194078 370226
rect 193458 370102 194078 370170
rect 193458 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 194078 370102
rect 193458 369978 194078 370046
rect 193458 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 194078 369978
rect 193458 352350 194078 369922
rect 194448 364350 194768 364384
rect 194448 364294 194518 364350
rect 194574 364294 194642 364350
rect 194698 364294 194768 364350
rect 194448 364226 194768 364294
rect 194448 364170 194518 364226
rect 194574 364170 194642 364226
rect 194698 364170 194768 364226
rect 194448 364102 194768 364170
rect 194448 364046 194518 364102
rect 194574 364046 194642 364102
rect 194698 364046 194768 364102
rect 194448 363978 194768 364046
rect 194448 363922 194518 363978
rect 194574 363922 194642 363978
rect 194698 363922 194768 363978
rect 194448 363888 194768 363922
rect 193458 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 194078 352350
rect 193458 352226 194078 352294
rect 193458 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 194078 352226
rect 193458 352102 194078 352170
rect 193458 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 194078 352102
rect 193458 351978 194078 352046
rect 193458 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 194078 351978
rect 193458 334350 194078 351922
rect 194448 346350 194768 346384
rect 194448 346294 194518 346350
rect 194574 346294 194642 346350
rect 194698 346294 194768 346350
rect 194448 346226 194768 346294
rect 194448 346170 194518 346226
rect 194574 346170 194642 346226
rect 194698 346170 194768 346226
rect 194448 346102 194768 346170
rect 194448 346046 194518 346102
rect 194574 346046 194642 346102
rect 194698 346046 194768 346102
rect 194448 345978 194768 346046
rect 194448 345922 194518 345978
rect 194574 345922 194642 345978
rect 194698 345922 194768 345978
rect 194448 345888 194768 345922
rect 193458 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 194078 334350
rect 193458 334226 194078 334294
rect 193458 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 194078 334226
rect 193458 334102 194078 334170
rect 193458 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 194078 334102
rect 193458 333978 194078 334046
rect 193458 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 194078 333978
rect 190652 323428 190708 323438
rect 190652 323332 190708 323342
rect 192332 323398 192388 323408
rect 189738 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 190358 310350
rect 189738 310226 190358 310294
rect 189738 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 190358 310226
rect 189738 310102 190358 310170
rect 189738 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 190358 310102
rect 189738 309978 190358 310046
rect 189738 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 190358 309978
rect 189738 292350 190358 309922
rect 189738 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 190358 292350
rect 189738 292226 190358 292294
rect 189738 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 190358 292226
rect 189738 292102 190358 292170
rect 189738 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 190358 292102
rect 189738 291978 190358 292046
rect 189738 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 190358 291978
rect 188076 286692 188132 286702
rect 188076 285778 188132 286636
rect 188076 285712 188132 285722
rect 187852 281392 187908 281402
rect 189738 274350 190358 291922
rect 189738 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 190358 274350
rect 189738 274226 190358 274294
rect 189738 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 190358 274226
rect 189738 274102 190358 274170
rect 189738 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 190358 274102
rect 189738 273978 190358 274046
rect 189738 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 190358 273978
rect 189738 256350 190358 273922
rect 189738 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 190358 256350
rect 189738 256226 190358 256294
rect 189738 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 190358 256226
rect 189738 256102 190358 256170
rect 189738 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 190358 256102
rect 189738 255978 190358 256046
rect 189738 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 190358 255978
rect 187740 221106 187796 221116
rect 187852 251524 187908 251534
rect 187628 216514 187684 216524
rect 187516 216402 187572 216412
rect 187852 214138 187908 251468
rect 187852 214072 187908 214082
rect 189738 238350 190358 255922
rect 189738 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 190358 238350
rect 189738 238226 190358 238294
rect 189738 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 190358 238226
rect 189738 238102 190358 238170
rect 189738 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 190358 238102
rect 189738 237978 190358 238046
rect 189738 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 190358 237978
rect 189738 220350 190358 237922
rect 189738 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 190358 220350
rect 189738 220226 190358 220294
rect 189738 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 190358 220226
rect 189738 220102 190358 220170
rect 189738 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 190358 220102
rect 189738 219978 190358 220046
rect 189738 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 190358 219978
rect 189738 210462 190358 219922
rect 190428 309316 190484 309326
rect 190428 209860 190484 309260
rect 190652 288484 190708 288494
rect 190540 285796 190596 285806
rect 190540 275940 190596 285740
rect 190540 250348 190596 275884
rect 190652 280420 190708 288428
rect 190652 255388 190708 280364
rect 190652 255332 191044 255388
rect 190540 250292 190932 250348
rect 190652 249844 190708 249854
rect 190652 249778 190708 249788
rect 190652 249712 190708 249722
rect 190652 248836 190708 248846
rect 190652 248698 190708 248780
rect 190652 248632 190708 248642
rect 190652 247268 190708 247296
rect 190652 247192 190708 247202
rect 190540 244804 190596 244814
rect 190540 231868 190596 244748
rect 190876 243118 190932 250292
rect 190876 243052 190932 243062
rect 190652 242676 190708 242686
rect 190652 242038 190708 242620
rect 190652 241972 190708 241982
rect 190988 238588 191044 255332
rect 190764 238532 191044 238588
rect 190652 235018 190708 235028
rect 190764 235018 190820 238532
rect 190708 234962 190820 235018
rect 190652 234952 190708 234962
rect 190540 231812 190932 231868
rect 190876 216132 190932 231812
rect 190876 216066 190932 216076
rect 192332 214498 192388 323342
rect 192332 214432 192388 214442
rect 193458 316350 194078 333922
rect 194448 328350 194768 328384
rect 194448 328294 194518 328350
rect 194574 328294 194642 328350
rect 194698 328294 194768 328350
rect 194448 328226 194768 328294
rect 194448 328170 194518 328226
rect 194574 328170 194642 328226
rect 194698 328170 194768 328226
rect 194448 328102 194768 328170
rect 194448 328046 194518 328102
rect 194574 328046 194642 328102
rect 194698 328046 194768 328102
rect 194448 327978 194768 328046
rect 194448 327922 194518 327978
rect 194574 327922 194642 327978
rect 194698 327922 194768 327978
rect 194448 327888 194768 327922
rect 193458 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 194078 316350
rect 193458 316226 194078 316294
rect 193458 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 194078 316226
rect 193458 316102 194078 316170
rect 193458 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 194078 316102
rect 193458 315978 194078 316046
rect 193458 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 194078 315978
rect 193458 298350 194078 315922
rect 194448 310350 194768 310384
rect 194448 310294 194518 310350
rect 194574 310294 194642 310350
rect 194698 310294 194768 310350
rect 194448 310226 194768 310294
rect 194448 310170 194518 310226
rect 194574 310170 194642 310226
rect 194698 310170 194768 310226
rect 194448 310102 194768 310170
rect 194448 310046 194518 310102
rect 194574 310046 194642 310102
rect 194698 310046 194768 310102
rect 194448 309978 194768 310046
rect 194448 309922 194518 309978
rect 194574 309922 194642 309978
rect 194698 309922 194768 309978
rect 194448 309888 194768 309922
rect 193458 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 194078 298350
rect 193458 298226 194078 298294
rect 193458 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 194078 298226
rect 193458 298102 194078 298170
rect 193458 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 194078 298102
rect 193458 297978 194078 298046
rect 193458 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 194078 297978
rect 193458 280350 194078 297922
rect 194448 292350 194768 292384
rect 194448 292294 194518 292350
rect 194574 292294 194642 292350
rect 194698 292294 194768 292350
rect 194448 292226 194768 292294
rect 194448 292170 194518 292226
rect 194574 292170 194642 292226
rect 194698 292170 194768 292226
rect 194448 292102 194768 292170
rect 194448 292046 194518 292102
rect 194574 292046 194642 292102
rect 194698 292046 194768 292102
rect 194448 291978 194768 292046
rect 194448 291922 194518 291978
rect 194574 291922 194642 291978
rect 194698 291922 194768 291978
rect 194448 291888 194768 291922
rect 193458 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 194078 280350
rect 193458 280226 194078 280294
rect 193458 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 194078 280226
rect 193458 280102 194078 280170
rect 193458 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 194078 280102
rect 193458 279978 194078 280046
rect 193458 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 194078 279978
rect 193458 262350 194078 279922
rect 194448 274350 194768 274384
rect 194448 274294 194518 274350
rect 194574 274294 194642 274350
rect 194698 274294 194768 274350
rect 194448 274226 194768 274294
rect 194448 274170 194518 274226
rect 194574 274170 194642 274226
rect 194698 274170 194768 274226
rect 194448 274102 194768 274170
rect 194448 274046 194518 274102
rect 194574 274046 194642 274102
rect 194698 274046 194768 274102
rect 194448 273978 194768 274046
rect 194448 273922 194518 273978
rect 194574 273922 194642 273978
rect 194698 273922 194768 273978
rect 194448 273888 194768 273922
rect 193458 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 194078 262350
rect 193458 262226 194078 262294
rect 193458 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 194078 262226
rect 193458 262102 194078 262170
rect 193458 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 194078 262102
rect 193458 261978 194078 262046
rect 193458 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 194078 261978
rect 193458 244350 194078 261922
rect 194448 256350 194768 256384
rect 194448 256294 194518 256350
rect 194574 256294 194642 256350
rect 194698 256294 194768 256350
rect 194448 256226 194768 256294
rect 194448 256170 194518 256226
rect 194574 256170 194642 256226
rect 194698 256170 194768 256226
rect 194448 256102 194768 256170
rect 194448 256046 194518 256102
rect 194574 256046 194642 256102
rect 194698 256046 194768 256102
rect 194448 255978 194768 256046
rect 194448 255922 194518 255978
rect 194574 255922 194642 255978
rect 194698 255922 194768 255978
rect 194448 255888 194768 255922
rect 193458 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 194078 244350
rect 193458 244226 194078 244294
rect 193458 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 194078 244226
rect 193458 244102 194078 244170
rect 193458 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 194078 244102
rect 193458 243978 194078 244046
rect 193458 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 194078 243978
rect 193458 226350 194078 243922
rect 193458 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 194078 226350
rect 193458 226226 194078 226294
rect 193458 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 194078 226226
rect 193458 226102 194078 226170
rect 193458 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 194078 226102
rect 193458 225978 194078 226046
rect 193458 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 194078 225978
rect 193458 210462 194078 225922
rect 194236 248698 194292 248708
rect 194236 214564 194292 248642
rect 194236 214498 194292 214508
rect 196476 211438 196532 372932
rect 197372 240212 197428 383740
rect 197484 287218 197540 391742
rect 198044 382004 198100 393182
rect 198156 382228 198212 401822
rect 199836 401698 199892 401708
rect 199724 393598 199780 393608
rect 198156 382162 198212 382172
rect 199500 383684 199556 383694
rect 198044 381938 198100 381948
rect 197596 378868 197652 378878
rect 197596 340138 197652 378812
rect 199388 373798 199444 373808
rect 197596 340072 197652 340082
rect 199276 368758 199332 368768
rect 197484 287152 197540 287162
rect 197596 289018 197652 289028
rect 197484 281458 197540 281468
rect 197484 240436 197540 281402
rect 197484 240370 197540 240380
rect 197372 240146 197428 240156
rect 197596 235956 197652 288962
rect 197708 285778 197764 285788
rect 197708 240324 197764 285722
rect 198044 268858 198100 268868
rect 197708 240258 197764 240268
rect 197820 249778 197876 249788
rect 197596 235890 197652 235900
rect 196476 211372 196532 211382
rect 197820 210898 197876 249722
rect 197932 247258 197988 247268
rect 197932 214318 197988 247202
rect 198044 241668 198100 268802
rect 198044 241602 198100 241612
rect 197932 214252 197988 214262
rect 199276 211258 199332 368702
rect 199388 214676 199444 373742
rect 199500 219604 199556 383628
rect 199724 382004 199780 393542
rect 199836 382228 199892 401642
rect 201516 393418 201572 393428
rect 199836 382162 199892 382172
rect 201404 391978 201460 391988
rect 199724 381938 199780 381948
rect 201404 382004 201460 391922
rect 201516 382228 201572 393362
rect 201516 382162 201572 382172
rect 204876 392158 204932 392168
rect 201404 381938 201460 381948
rect 204876 382004 204932 392102
rect 204876 381938 204932 381948
rect 206556 382004 206612 404162
rect 208236 382228 208292 404342
rect 208236 382162 208292 382172
rect 209916 382228 209972 404522
rect 220458 400350 221078 410034
rect 220458 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 221078 400350
rect 220458 400226 221078 400294
rect 220458 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 221078 400226
rect 220458 400102 221078 400170
rect 220458 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 221078 400102
rect 220458 399978 221078 400046
rect 220458 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 221078 399978
rect 215068 391438 215124 391448
rect 215068 390964 215124 391382
rect 216636 391438 216692 391448
rect 216636 391344 216692 391356
rect 215068 390898 215124 390908
rect 209916 382162 209972 382172
rect 220458 382350 221078 399922
rect 220458 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 221078 382350
rect 220458 382226 221078 382294
rect 220458 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 221078 382226
rect 220458 382102 221078 382170
rect 220458 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 221078 382102
rect 206556 381938 206612 381948
rect 206780 382004 206836 382014
rect 199836 381892 199892 381902
rect 199500 219538 199556 219548
rect 199612 381444 199668 381454
rect 199612 216356 199668 381388
rect 199836 372988 199892 381836
rect 206780 381444 206836 381948
rect 206780 381378 206836 381388
rect 220458 381978 221078 382046
rect 220458 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 221078 381978
rect 210364 379764 210420 379774
rect 202412 379652 202468 379662
rect 202412 379204 202468 379596
rect 202412 379138 202468 379148
rect 210364 378868 210420 379708
rect 210364 378802 210420 378812
rect 199612 216290 199668 216300
rect 199724 372932 199892 372988
rect 199724 216244 199780 372932
rect 209808 370350 210128 370384
rect 209808 370294 209878 370350
rect 209934 370294 210002 370350
rect 210058 370294 210128 370350
rect 209808 370226 210128 370294
rect 209808 370170 209878 370226
rect 209934 370170 210002 370226
rect 210058 370170 210128 370226
rect 209808 370102 210128 370170
rect 209808 370046 209878 370102
rect 209934 370046 210002 370102
rect 210058 370046 210128 370102
rect 209808 369978 210128 370046
rect 209808 369922 209878 369978
rect 209934 369922 210002 369978
rect 210058 369922 210128 369978
rect 209808 369888 210128 369922
rect 220458 367758 221078 381922
rect 224178 406350 224798 410034
rect 243516 407988 243572 407998
rect 243516 407638 243572 407932
rect 243516 407572 243572 407582
rect 248892 407540 248948 407550
rect 248892 406918 248948 407484
rect 248892 406852 248948 406862
rect 224178 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 224798 406350
rect 224178 406226 224798 406294
rect 224178 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 224798 406226
rect 224178 406102 224798 406170
rect 224178 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 224798 406102
rect 224178 405978 224798 406046
rect 224178 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 224798 405978
rect 224178 388350 224798 405922
rect 227612 406738 227668 406748
rect 227612 406644 227668 406682
rect 227612 395780 227668 406588
rect 227612 395714 227668 395724
rect 251178 400350 251798 410034
rect 251178 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 251798 400350
rect 251178 400226 251798 400294
rect 251178 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 251798 400226
rect 251178 400102 251798 400170
rect 251178 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 251798 400102
rect 251178 399978 251798 400046
rect 251178 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 251798 399978
rect 231644 395218 231700 395228
rect 224178 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 224798 388350
rect 224178 388226 224798 388294
rect 224178 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 224798 388226
rect 224178 388102 224798 388170
rect 224178 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 224798 388102
rect 224178 387978 224798 388046
rect 224178 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 224798 387978
rect 221564 379502 221956 379558
rect 221564 379428 221620 379502
rect 221564 379362 221620 379372
rect 221788 379428 221844 379438
rect 221788 378868 221844 379372
rect 221900 379204 221956 379502
rect 221900 379138 221956 379148
rect 222684 379428 222740 379438
rect 222684 378980 222740 379372
rect 222684 378914 222740 378924
rect 221788 378802 221844 378812
rect 224178 370350 224798 387922
rect 230076 393778 230132 393788
rect 230076 382228 230132 393722
rect 231644 382340 231700 395162
rect 231644 382274 231700 382284
rect 231756 395038 231812 395048
rect 230076 382162 230132 382172
rect 231756 382228 231812 394982
rect 231756 382162 231812 382172
rect 251178 382350 251798 399922
rect 251178 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 251798 382350
rect 251178 382226 251798 382294
rect 251178 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 251798 382226
rect 251178 382102 251798 382170
rect 251178 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 251798 382102
rect 251178 381978 251798 382046
rect 251178 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 251798 381978
rect 236124 379764 236180 379774
rect 236124 379670 236180 379682
rect 224178 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 224798 370350
rect 224178 370226 224798 370294
rect 224178 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 224798 370226
rect 224178 370102 224798 370170
rect 224178 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 224798 370102
rect 224178 369978 224798 370046
rect 224178 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 224798 369978
rect 224178 367758 224798 369922
rect 235228 379428 235284 379438
rect 235228 368758 235284 379372
rect 237020 379428 237076 379438
rect 237020 373798 237076 379372
rect 237020 373732 237076 373742
rect 238476 379428 238532 379438
rect 250124 379428 250180 379438
rect 235228 368692 235284 368702
rect 238476 368758 238532 379372
rect 249116 379372 250124 379378
rect 249116 379322 250180 379372
rect 249116 379316 249172 379322
rect 249116 379250 249172 379260
rect 249340 379204 249396 379214
rect 250012 379204 250068 379214
rect 249396 379148 250012 379198
rect 249340 379142 250068 379148
rect 249340 379138 249396 379142
rect 250012 379138 250068 379142
rect 240528 370350 240848 370384
rect 240528 370294 240598 370350
rect 240654 370294 240722 370350
rect 240778 370294 240848 370350
rect 240528 370226 240848 370294
rect 240528 370170 240598 370226
rect 240654 370170 240722 370226
rect 240778 370170 240848 370226
rect 240528 370102 240848 370170
rect 240528 370046 240598 370102
rect 240654 370046 240722 370102
rect 240778 370046 240848 370102
rect 240528 369978 240848 370046
rect 240528 369922 240598 369978
rect 240654 369922 240722 369978
rect 240778 369922 240848 369978
rect 240528 369888 240848 369922
rect 238476 368692 238532 368702
rect 251178 367758 251798 381922
rect 254898 406350 255518 410034
rect 277116 407458 277172 407468
rect 254898 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 255518 406350
rect 254898 406226 255518 406294
rect 254898 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 255518 406226
rect 254898 406102 255518 406170
rect 254898 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 255518 406102
rect 254898 405978 255518 406046
rect 254898 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 255518 405978
rect 254898 388350 255518 405922
rect 254898 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 255518 388350
rect 254898 388226 255518 388294
rect 254898 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 255518 388226
rect 254898 388102 255518 388170
rect 254898 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 255518 388102
rect 254898 387978 255518 388046
rect 254898 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 255518 387978
rect 253372 379540 253428 379550
rect 253372 378980 253428 379484
rect 253372 378914 253428 378924
rect 254898 370350 255518 387922
rect 266252 406644 266308 406654
rect 264460 379428 264516 379438
rect 264460 379092 264516 379372
rect 264460 379026 264516 379036
rect 254898 370294 254994 370350
rect 255050 370294 255118 370350
rect 255174 370294 255242 370350
rect 255298 370294 255366 370350
rect 255422 370294 255518 370350
rect 254898 370226 255518 370294
rect 254898 370170 254994 370226
rect 255050 370170 255118 370226
rect 255174 370170 255242 370226
rect 255298 370170 255366 370226
rect 255422 370170 255518 370226
rect 254898 370102 255518 370170
rect 254898 370046 254994 370102
rect 255050 370046 255118 370102
rect 255174 370046 255242 370102
rect 255298 370046 255366 370102
rect 255422 370046 255518 370102
rect 254898 369978 255518 370046
rect 254898 369922 254994 369978
rect 255050 369922 255118 369978
rect 255174 369922 255242 369978
rect 255298 369922 255366 369978
rect 255422 369922 255518 369978
rect 254898 367758 255518 369922
rect 266252 368938 266308 406588
rect 266252 368872 266308 368882
rect 270396 406644 270452 406654
rect 270396 367858 270452 406588
rect 276332 406644 276388 406654
rect 276332 373078 276388 406588
rect 277116 382116 277172 407402
rect 277116 382050 277172 382060
rect 281372 406644 281428 406654
rect 281372 373798 281428 406588
rect 281372 373732 281428 373742
rect 281898 400350 282518 410034
rect 281898 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 282518 400350
rect 281898 400226 282518 400294
rect 281898 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 282518 400226
rect 281898 400102 282518 400170
rect 281898 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 282518 400102
rect 281898 399978 282518 400046
rect 281898 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 282518 399978
rect 281898 382350 282518 399922
rect 281898 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 282518 382350
rect 281898 382226 282518 382294
rect 281898 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 282518 382226
rect 281898 382102 282518 382170
rect 281898 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 282518 382102
rect 281898 381978 282518 382046
rect 281898 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 282518 381978
rect 271248 370350 271568 370384
rect 271248 370294 271318 370350
rect 271374 370294 271442 370350
rect 271498 370294 271568 370350
rect 271248 370226 271568 370294
rect 271248 370170 271318 370226
rect 271374 370170 271442 370226
rect 271498 370170 271568 370226
rect 271248 370102 271568 370170
rect 271248 370046 271318 370102
rect 271374 370046 271442 370102
rect 271498 370046 271568 370102
rect 271248 369978 271568 370046
rect 271248 369922 271318 369978
rect 271374 369922 271442 369978
rect 271498 369922 271568 369978
rect 271248 369888 271568 369922
rect 270396 367802 270564 367858
rect 270508 365878 270564 367802
rect 276332 367138 276388 373022
rect 281898 367758 282518 381922
rect 285618 406350 286238 410034
rect 285618 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 286238 406350
rect 285618 406226 286238 406294
rect 285618 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 286238 406226
rect 285618 406102 286238 406170
rect 285618 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 286238 406102
rect 285618 405978 286238 406046
rect 285618 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 286238 405978
rect 285618 388350 286238 405922
rect 285618 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 286238 388350
rect 285618 388226 286238 388294
rect 285618 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 286238 388226
rect 285618 388102 286238 388170
rect 285618 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 286238 388102
rect 285618 387978 286238 388046
rect 285618 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 286238 387978
rect 285618 370350 286238 387922
rect 286412 406644 286468 406654
rect 286412 372178 286468 406588
rect 312618 400350 313238 410034
rect 312618 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 313238 400350
rect 312618 400226 313238 400294
rect 312618 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 313238 400226
rect 312618 400102 313238 400170
rect 312618 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 313238 400102
rect 312618 399978 313238 400046
rect 312618 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 313238 399978
rect 307356 399178 307412 399188
rect 305676 398998 305732 399008
rect 305676 382116 305732 398942
rect 305676 382050 305732 382060
rect 307356 382116 307412 399122
rect 307356 382050 307412 382060
rect 312618 382350 313238 399922
rect 312618 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 313238 382350
rect 312618 382226 313238 382294
rect 312618 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 313238 382226
rect 312618 382102 313238 382170
rect 286412 372112 286468 372122
rect 312618 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 313238 382102
rect 312618 381978 313238 382046
rect 312618 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 313238 381978
rect 285618 370294 285714 370350
rect 285770 370294 285838 370350
rect 285894 370294 285962 370350
rect 286018 370294 286086 370350
rect 286142 370294 286238 370350
rect 285618 370226 286238 370294
rect 285618 370170 285714 370226
rect 285770 370170 285838 370226
rect 285894 370170 285962 370226
rect 286018 370170 286086 370226
rect 286142 370170 286238 370226
rect 285618 370102 286238 370170
rect 285618 370046 285714 370102
rect 285770 370046 285838 370102
rect 285894 370046 285962 370102
rect 286018 370046 286086 370102
rect 286142 370046 286238 370102
rect 285618 369978 286238 370046
rect 285618 369922 285714 369978
rect 285770 369922 285838 369978
rect 285894 369922 285962 369978
rect 286018 369922 286086 369978
rect 286142 369922 286238 369978
rect 285618 367758 286238 369922
rect 301968 370350 302288 370384
rect 301968 370294 302038 370350
rect 302094 370294 302162 370350
rect 302218 370294 302288 370350
rect 301968 370226 302288 370294
rect 301968 370170 302038 370226
rect 302094 370170 302162 370226
rect 302218 370170 302288 370226
rect 301968 370102 302288 370170
rect 301968 370046 302038 370102
rect 302094 370046 302162 370102
rect 302218 370046 302288 370102
rect 301968 369978 302288 370046
rect 301968 369922 302038 369978
rect 302094 369922 302162 369978
rect 302218 369922 302288 369978
rect 301968 369888 302288 369922
rect 312618 367758 313238 381922
rect 316338 406350 316958 410034
rect 316338 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 316958 406350
rect 316338 406226 316958 406294
rect 316338 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 316958 406226
rect 316338 406102 316958 406170
rect 316338 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 316958 406102
rect 316338 405978 316958 406046
rect 316338 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 316958 405978
rect 316338 388350 316958 405922
rect 323372 406644 323428 406654
rect 316338 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 316958 388350
rect 316338 388226 316958 388294
rect 316338 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 316958 388226
rect 316338 388102 316958 388170
rect 316338 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 316958 388102
rect 316338 387978 316958 388046
rect 316338 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 316958 387978
rect 316338 370350 316958 387922
rect 319116 400618 319172 400628
rect 319116 382116 319172 400562
rect 319116 382050 319172 382060
rect 320796 399358 320852 399368
rect 320796 382116 320852 399302
rect 320796 382050 320852 382060
rect 323372 376318 323428 406588
rect 324156 382116 324212 410642
rect 329196 409258 329252 409268
rect 324156 382050 324212 382060
rect 329084 388164 329140 388174
rect 323372 376252 323428 376262
rect 316338 370294 316434 370350
rect 316490 370294 316558 370350
rect 316614 370294 316682 370350
rect 316738 370294 316806 370350
rect 316862 370294 316958 370350
rect 316338 370226 316958 370294
rect 316338 370170 316434 370226
rect 316490 370170 316558 370226
rect 316614 370170 316682 370226
rect 316738 370170 316806 370226
rect 316862 370170 316958 370226
rect 316338 370102 316958 370170
rect 316338 370046 316434 370102
rect 316490 370046 316558 370102
rect 316614 370046 316682 370102
rect 316738 370046 316806 370102
rect 316862 370046 316958 370102
rect 316338 369978 316958 370046
rect 316338 369922 316434 369978
rect 316490 369922 316558 369978
rect 316614 369922 316682 369978
rect 316738 369922 316806 369978
rect 316862 369922 316958 369978
rect 316338 367758 316958 369922
rect 329084 369118 329140 388108
rect 329196 382116 329252 409202
rect 329196 382050 329252 382060
rect 330876 405658 330932 405668
rect 330876 382116 330932 405602
rect 330876 382050 330932 382060
rect 334236 382116 334292 410822
rect 339276 408996 339332 409006
rect 334236 382050 334292 382060
rect 335916 406644 335972 406654
rect 332688 370350 333008 370384
rect 332688 370294 332758 370350
rect 332814 370294 332882 370350
rect 332938 370294 333008 370350
rect 332688 370226 333008 370294
rect 332688 370170 332758 370226
rect 332814 370170 332882 370226
rect 332938 370170 333008 370226
rect 332688 370102 333008 370170
rect 332688 370046 332758 370102
rect 332814 370046 332882 370102
rect 332938 370046 333008 370102
rect 332688 369978 333008 370046
rect 332688 369922 332758 369978
rect 332814 369922 332882 369978
rect 332938 369922 333008 369978
rect 332688 369888 333008 369922
rect 329084 369052 329140 369062
rect 276332 367072 276388 367082
rect 270508 365812 270564 365822
rect 272076 366598 272132 366608
rect 272076 365878 272132 366542
rect 272076 365812 272132 365822
rect 225168 364350 225488 364384
rect 225168 364294 225238 364350
rect 225294 364294 225362 364350
rect 225418 364294 225488 364350
rect 225168 364226 225488 364294
rect 225168 364170 225238 364226
rect 225294 364170 225362 364226
rect 225418 364170 225488 364226
rect 225168 364102 225488 364170
rect 225168 364046 225238 364102
rect 225294 364046 225362 364102
rect 225418 364046 225488 364102
rect 225168 363978 225488 364046
rect 225168 363922 225238 363978
rect 225294 363922 225362 363978
rect 225418 363922 225488 363978
rect 225168 363888 225488 363922
rect 255888 364350 256208 364384
rect 255888 364294 255958 364350
rect 256014 364294 256082 364350
rect 256138 364294 256208 364350
rect 255888 364226 256208 364294
rect 255888 364170 255958 364226
rect 256014 364170 256082 364226
rect 256138 364170 256208 364226
rect 255888 364102 256208 364170
rect 255888 364046 255958 364102
rect 256014 364046 256082 364102
rect 256138 364046 256208 364102
rect 255888 363978 256208 364046
rect 255888 363922 255958 363978
rect 256014 363922 256082 363978
rect 256138 363922 256208 363978
rect 255888 363888 256208 363922
rect 286608 364350 286928 364384
rect 286608 364294 286678 364350
rect 286734 364294 286802 364350
rect 286858 364294 286928 364350
rect 286608 364226 286928 364294
rect 286608 364170 286678 364226
rect 286734 364170 286802 364226
rect 286858 364170 286928 364226
rect 286608 364102 286928 364170
rect 286608 364046 286678 364102
rect 286734 364046 286802 364102
rect 286858 364046 286928 364102
rect 286608 363978 286928 364046
rect 286608 363922 286678 363978
rect 286734 363922 286802 363978
rect 286858 363922 286928 363978
rect 286608 363888 286928 363922
rect 317328 364350 317648 364384
rect 317328 364294 317398 364350
rect 317454 364294 317522 364350
rect 317578 364294 317648 364350
rect 317328 364226 317648 364294
rect 317328 364170 317398 364226
rect 317454 364170 317522 364226
rect 317578 364170 317648 364226
rect 317328 364102 317648 364170
rect 317328 364046 317398 364102
rect 317454 364046 317522 364102
rect 317578 364046 317648 364102
rect 317328 363978 317648 364046
rect 317328 363922 317398 363978
rect 317454 363922 317522 363978
rect 317578 363922 317648 363978
rect 317328 363888 317648 363922
rect 335916 356158 335972 406588
rect 338492 385812 338548 385822
rect 336924 380548 336980 380558
rect 336812 379540 336868 379550
rect 335916 356092 335972 356102
rect 336028 368758 336084 368768
rect 209808 352350 210128 352384
rect 209808 352294 209878 352350
rect 209934 352294 210002 352350
rect 210058 352294 210128 352350
rect 209808 352226 210128 352294
rect 209808 352170 209878 352226
rect 209934 352170 210002 352226
rect 210058 352170 210128 352226
rect 209808 352102 210128 352170
rect 209808 352046 209878 352102
rect 209934 352046 210002 352102
rect 210058 352046 210128 352102
rect 209808 351978 210128 352046
rect 209808 351922 209878 351978
rect 209934 351922 210002 351978
rect 210058 351922 210128 351978
rect 209808 351888 210128 351922
rect 240528 352350 240848 352384
rect 240528 352294 240598 352350
rect 240654 352294 240722 352350
rect 240778 352294 240848 352350
rect 240528 352226 240848 352294
rect 240528 352170 240598 352226
rect 240654 352170 240722 352226
rect 240778 352170 240848 352226
rect 240528 352102 240848 352170
rect 240528 352046 240598 352102
rect 240654 352046 240722 352102
rect 240778 352046 240848 352102
rect 240528 351978 240848 352046
rect 240528 351922 240598 351978
rect 240654 351922 240722 351978
rect 240778 351922 240848 351978
rect 240528 351888 240848 351922
rect 271248 352350 271568 352384
rect 271248 352294 271318 352350
rect 271374 352294 271442 352350
rect 271498 352294 271568 352350
rect 271248 352226 271568 352294
rect 271248 352170 271318 352226
rect 271374 352170 271442 352226
rect 271498 352170 271568 352226
rect 271248 352102 271568 352170
rect 271248 352046 271318 352102
rect 271374 352046 271442 352102
rect 271498 352046 271568 352102
rect 271248 351978 271568 352046
rect 271248 351922 271318 351978
rect 271374 351922 271442 351978
rect 271498 351922 271568 351978
rect 271248 351888 271568 351922
rect 301968 352350 302288 352384
rect 301968 352294 302038 352350
rect 302094 352294 302162 352350
rect 302218 352294 302288 352350
rect 301968 352226 302288 352294
rect 301968 352170 302038 352226
rect 302094 352170 302162 352226
rect 302218 352170 302288 352226
rect 301968 352102 302288 352170
rect 301968 352046 302038 352102
rect 302094 352046 302162 352102
rect 302218 352046 302288 352102
rect 301968 351978 302288 352046
rect 301968 351922 302038 351978
rect 302094 351922 302162 351978
rect 302218 351922 302288 351978
rect 301968 351888 302288 351922
rect 332688 352350 333008 352384
rect 332688 352294 332758 352350
rect 332814 352294 332882 352350
rect 332938 352294 333008 352350
rect 332688 352226 333008 352294
rect 332688 352170 332758 352226
rect 332814 352170 332882 352226
rect 332938 352170 333008 352226
rect 332688 352102 333008 352170
rect 332688 352046 332758 352102
rect 332814 352046 332882 352102
rect 332938 352046 333008 352102
rect 332688 351978 333008 352046
rect 332688 351922 332758 351978
rect 332814 351922 332882 351978
rect 332938 351922 333008 351978
rect 332688 351888 333008 351922
rect 225168 346350 225488 346384
rect 225168 346294 225238 346350
rect 225294 346294 225362 346350
rect 225418 346294 225488 346350
rect 225168 346226 225488 346294
rect 225168 346170 225238 346226
rect 225294 346170 225362 346226
rect 225418 346170 225488 346226
rect 225168 346102 225488 346170
rect 225168 346046 225238 346102
rect 225294 346046 225362 346102
rect 225418 346046 225488 346102
rect 225168 345978 225488 346046
rect 225168 345922 225238 345978
rect 225294 345922 225362 345978
rect 225418 345922 225488 345978
rect 225168 345888 225488 345922
rect 255888 346350 256208 346384
rect 255888 346294 255958 346350
rect 256014 346294 256082 346350
rect 256138 346294 256208 346350
rect 255888 346226 256208 346294
rect 255888 346170 255958 346226
rect 256014 346170 256082 346226
rect 256138 346170 256208 346226
rect 255888 346102 256208 346170
rect 255888 346046 255958 346102
rect 256014 346046 256082 346102
rect 256138 346046 256208 346102
rect 255888 345978 256208 346046
rect 255888 345922 255958 345978
rect 256014 345922 256082 345978
rect 256138 345922 256208 345978
rect 255888 345888 256208 345922
rect 286608 346350 286928 346384
rect 286608 346294 286678 346350
rect 286734 346294 286802 346350
rect 286858 346294 286928 346350
rect 286608 346226 286928 346294
rect 286608 346170 286678 346226
rect 286734 346170 286802 346226
rect 286858 346170 286928 346226
rect 286608 346102 286928 346170
rect 286608 346046 286678 346102
rect 286734 346046 286802 346102
rect 286858 346046 286928 346102
rect 286608 345978 286928 346046
rect 286608 345922 286678 345978
rect 286734 345922 286802 345978
rect 286858 345922 286928 345978
rect 286608 345888 286928 345922
rect 317328 346350 317648 346384
rect 317328 346294 317398 346350
rect 317454 346294 317522 346350
rect 317578 346294 317648 346350
rect 317328 346226 317648 346294
rect 317328 346170 317398 346226
rect 317454 346170 317522 346226
rect 317578 346170 317648 346226
rect 317328 346102 317648 346170
rect 317328 346046 317398 346102
rect 317454 346046 317522 346102
rect 317578 346046 317648 346102
rect 317328 345978 317648 346046
rect 317328 345922 317398 345978
rect 317454 345922 317522 345978
rect 317578 345922 317648 345978
rect 317328 345888 317648 345922
rect 209808 334350 210128 334384
rect 209808 334294 209878 334350
rect 209934 334294 210002 334350
rect 210058 334294 210128 334350
rect 209808 334226 210128 334294
rect 209808 334170 209878 334226
rect 209934 334170 210002 334226
rect 210058 334170 210128 334226
rect 209808 334102 210128 334170
rect 209808 334046 209878 334102
rect 209934 334046 210002 334102
rect 210058 334046 210128 334102
rect 209808 333978 210128 334046
rect 209808 333922 209878 333978
rect 209934 333922 210002 333978
rect 210058 333922 210128 333978
rect 209808 333888 210128 333922
rect 240528 334350 240848 334384
rect 240528 334294 240598 334350
rect 240654 334294 240722 334350
rect 240778 334294 240848 334350
rect 240528 334226 240848 334294
rect 240528 334170 240598 334226
rect 240654 334170 240722 334226
rect 240778 334170 240848 334226
rect 240528 334102 240848 334170
rect 240528 334046 240598 334102
rect 240654 334046 240722 334102
rect 240778 334046 240848 334102
rect 240528 333978 240848 334046
rect 240528 333922 240598 333978
rect 240654 333922 240722 333978
rect 240778 333922 240848 333978
rect 240528 333888 240848 333922
rect 271248 334350 271568 334384
rect 271248 334294 271318 334350
rect 271374 334294 271442 334350
rect 271498 334294 271568 334350
rect 271248 334226 271568 334294
rect 271248 334170 271318 334226
rect 271374 334170 271442 334226
rect 271498 334170 271568 334226
rect 271248 334102 271568 334170
rect 271248 334046 271318 334102
rect 271374 334046 271442 334102
rect 271498 334046 271568 334102
rect 271248 333978 271568 334046
rect 271248 333922 271318 333978
rect 271374 333922 271442 333978
rect 271498 333922 271568 333978
rect 271248 333888 271568 333922
rect 301968 334350 302288 334384
rect 301968 334294 302038 334350
rect 302094 334294 302162 334350
rect 302218 334294 302288 334350
rect 301968 334226 302288 334294
rect 301968 334170 302038 334226
rect 302094 334170 302162 334226
rect 302218 334170 302288 334226
rect 301968 334102 302288 334170
rect 301968 334046 302038 334102
rect 302094 334046 302162 334102
rect 302218 334046 302288 334102
rect 301968 333978 302288 334046
rect 301968 333922 302038 333978
rect 302094 333922 302162 333978
rect 302218 333922 302288 333978
rect 301968 333888 302288 333922
rect 332688 334350 333008 334384
rect 332688 334294 332758 334350
rect 332814 334294 332882 334350
rect 332938 334294 333008 334350
rect 332688 334226 333008 334294
rect 332688 334170 332758 334226
rect 332814 334170 332882 334226
rect 332938 334170 333008 334226
rect 332688 334102 333008 334170
rect 332688 334046 332758 334102
rect 332814 334046 332882 334102
rect 332938 334046 333008 334102
rect 332688 333978 333008 334046
rect 332688 333922 332758 333978
rect 332814 333922 332882 333978
rect 332938 333922 333008 333978
rect 332688 333888 333008 333922
rect 225168 328350 225488 328384
rect 225168 328294 225238 328350
rect 225294 328294 225362 328350
rect 225418 328294 225488 328350
rect 225168 328226 225488 328294
rect 225168 328170 225238 328226
rect 225294 328170 225362 328226
rect 225418 328170 225488 328226
rect 225168 328102 225488 328170
rect 225168 328046 225238 328102
rect 225294 328046 225362 328102
rect 225418 328046 225488 328102
rect 225168 327978 225488 328046
rect 225168 327922 225238 327978
rect 225294 327922 225362 327978
rect 225418 327922 225488 327978
rect 225168 327888 225488 327922
rect 255888 328350 256208 328384
rect 255888 328294 255958 328350
rect 256014 328294 256082 328350
rect 256138 328294 256208 328350
rect 255888 328226 256208 328294
rect 255888 328170 255958 328226
rect 256014 328170 256082 328226
rect 256138 328170 256208 328226
rect 255888 328102 256208 328170
rect 255888 328046 255958 328102
rect 256014 328046 256082 328102
rect 256138 328046 256208 328102
rect 255888 327978 256208 328046
rect 255888 327922 255958 327978
rect 256014 327922 256082 327978
rect 256138 327922 256208 327978
rect 255888 327888 256208 327922
rect 286608 328350 286928 328384
rect 286608 328294 286678 328350
rect 286734 328294 286802 328350
rect 286858 328294 286928 328350
rect 286608 328226 286928 328294
rect 286608 328170 286678 328226
rect 286734 328170 286802 328226
rect 286858 328170 286928 328226
rect 286608 328102 286928 328170
rect 286608 328046 286678 328102
rect 286734 328046 286802 328102
rect 286858 328046 286928 328102
rect 286608 327978 286928 328046
rect 286608 327922 286678 327978
rect 286734 327922 286802 327978
rect 286858 327922 286928 327978
rect 286608 327888 286928 327922
rect 317328 328350 317648 328384
rect 317328 328294 317398 328350
rect 317454 328294 317522 328350
rect 317578 328294 317648 328350
rect 317328 328226 317648 328294
rect 317328 328170 317398 328226
rect 317454 328170 317522 328226
rect 317578 328170 317648 328226
rect 317328 328102 317648 328170
rect 317328 328046 317398 328102
rect 317454 328046 317522 328102
rect 317578 328046 317648 328102
rect 317328 327978 317648 328046
rect 317328 327922 317398 327978
rect 317454 327922 317522 327978
rect 317578 327922 317648 327978
rect 317328 327888 317648 327922
rect 209808 316350 210128 316384
rect 209808 316294 209878 316350
rect 209934 316294 210002 316350
rect 210058 316294 210128 316350
rect 209808 316226 210128 316294
rect 209808 316170 209878 316226
rect 209934 316170 210002 316226
rect 210058 316170 210128 316226
rect 209808 316102 210128 316170
rect 209808 316046 209878 316102
rect 209934 316046 210002 316102
rect 210058 316046 210128 316102
rect 209808 315978 210128 316046
rect 209808 315922 209878 315978
rect 209934 315922 210002 315978
rect 210058 315922 210128 315978
rect 209808 315888 210128 315922
rect 240528 316350 240848 316384
rect 240528 316294 240598 316350
rect 240654 316294 240722 316350
rect 240778 316294 240848 316350
rect 240528 316226 240848 316294
rect 240528 316170 240598 316226
rect 240654 316170 240722 316226
rect 240778 316170 240848 316226
rect 240528 316102 240848 316170
rect 240528 316046 240598 316102
rect 240654 316046 240722 316102
rect 240778 316046 240848 316102
rect 240528 315978 240848 316046
rect 240528 315922 240598 315978
rect 240654 315922 240722 315978
rect 240778 315922 240848 315978
rect 240528 315888 240848 315922
rect 271248 316350 271568 316384
rect 271248 316294 271318 316350
rect 271374 316294 271442 316350
rect 271498 316294 271568 316350
rect 271248 316226 271568 316294
rect 271248 316170 271318 316226
rect 271374 316170 271442 316226
rect 271498 316170 271568 316226
rect 271248 316102 271568 316170
rect 271248 316046 271318 316102
rect 271374 316046 271442 316102
rect 271498 316046 271568 316102
rect 271248 315978 271568 316046
rect 271248 315922 271318 315978
rect 271374 315922 271442 315978
rect 271498 315922 271568 315978
rect 271248 315888 271568 315922
rect 301968 316350 302288 316384
rect 301968 316294 302038 316350
rect 302094 316294 302162 316350
rect 302218 316294 302288 316350
rect 301968 316226 302288 316294
rect 301968 316170 302038 316226
rect 302094 316170 302162 316226
rect 302218 316170 302288 316226
rect 301968 316102 302288 316170
rect 301968 316046 302038 316102
rect 302094 316046 302162 316102
rect 302218 316046 302288 316102
rect 301968 315978 302288 316046
rect 301968 315922 302038 315978
rect 302094 315922 302162 315978
rect 302218 315922 302288 315978
rect 301968 315888 302288 315922
rect 332688 316350 333008 316384
rect 332688 316294 332758 316350
rect 332814 316294 332882 316350
rect 332938 316294 333008 316350
rect 332688 316226 333008 316294
rect 332688 316170 332758 316226
rect 332814 316170 332882 316226
rect 332938 316170 333008 316226
rect 332688 316102 333008 316170
rect 332688 316046 332758 316102
rect 332814 316046 332882 316102
rect 332938 316046 333008 316102
rect 332688 315978 333008 316046
rect 332688 315922 332758 315978
rect 332814 315922 332882 315978
rect 332938 315922 333008 315978
rect 332688 315888 333008 315922
rect 225168 310350 225488 310384
rect 225168 310294 225238 310350
rect 225294 310294 225362 310350
rect 225418 310294 225488 310350
rect 225168 310226 225488 310294
rect 225168 310170 225238 310226
rect 225294 310170 225362 310226
rect 225418 310170 225488 310226
rect 225168 310102 225488 310170
rect 225168 310046 225238 310102
rect 225294 310046 225362 310102
rect 225418 310046 225488 310102
rect 225168 309978 225488 310046
rect 225168 309922 225238 309978
rect 225294 309922 225362 309978
rect 225418 309922 225488 309978
rect 225168 309888 225488 309922
rect 255888 310350 256208 310384
rect 255888 310294 255958 310350
rect 256014 310294 256082 310350
rect 256138 310294 256208 310350
rect 255888 310226 256208 310294
rect 255888 310170 255958 310226
rect 256014 310170 256082 310226
rect 256138 310170 256208 310226
rect 255888 310102 256208 310170
rect 255888 310046 255958 310102
rect 256014 310046 256082 310102
rect 256138 310046 256208 310102
rect 255888 309978 256208 310046
rect 255888 309922 255958 309978
rect 256014 309922 256082 309978
rect 256138 309922 256208 309978
rect 255888 309888 256208 309922
rect 286608 310350 286928 310384
rect 286608 310294 286678 310350
rect 286734 310294 286802 310350
rect 286858 310294 286928 310350
rect 286608 310226 286928 310294
rect 286608 310170 286678 310226
rect 286734 310170 286802 310226
rect 286858 310170 286928 310226
rect 286608 310102 286928 310170
rect 286608 310046 286678 310102
rect 286734 310046 286802 310102
rect 286858 310046 286928 310102
rect 286608 309978 286928 310046
rect 286608 309922 286678 309978
rect 286734 309922 286802 309978
rect 286858 309922 286928 309978
rect 286608 309888 286928 309922
rect 317328 310350 317648 310384
rect 317328 310294 317398 310350
rect 317454 310294 317522 310350
rect 317578 310294 317648 310350
rect 317328 310226 317648 310294
rect 317328 310170 317398 310226
rect 317454 310170 317522 310226
rect 317578 310170 317648 310226
rect 317328 310102 317648 310170
rect 317328 310046 317398 310102
rect 317454 310046 317522 310102
rect 317578 310046 317648 310102
rect 317328 309978 317648 310046
rect 317328 309922 317398 309978
rect 317454 309922 317522 309978
rect 317578 309922 317648 309978
rect 317328 309888 317648 309922
rect 209808 298350 210128 298384
rect 209808 298294 209878 298350
rect 209934 298294 210002 298350
rect 210058 298294 210128 298350
rect 209808 298226 210128 298294
rect 209808 298170 209878 298226
rect 209934 298170 210002 298226
rect 210058 298170 210128 298226
rect 209808 298102 210128 298170
rect 209808 298046 209878 298102
rect 209934 298046 210002 298102
rect 210058 298046 210128 298102
rect 209808 297978 210128 298046
rect 209808 297922 209878 297978
rect 209934 297922 210002 297978
rect 210058 297922 210128 297978
rect 209808 297888 210128 297922
rect 240528 298350 240848 298384
rect 240528 298294 240598 298350
rect 240654 298294 240722 298350
rect 240778 298294 240848 298350
rect 240528 298226 240848 298294
rect 240528 298170 240598 298226
rect 240654 298170 240722 298226
rect 240778 298170 240848 298226
rect 240528 298102 240848 298170
rect 240528 298046 240598 298102
rect 240654 298046 240722 298102
rect 240778 298046 240848 298102
rect 240528 297978 240848 298046
rect 240528 297922 240598 297978
rect 240654 297922 240722 297978
rect 240778 297922 240848 297978
rect 240528 297888 240848 297922
rect 271248 298350 271568 298384
rect 271248 298294 271318 298350
rect 271374 298294 271442 298350
rect 271498 298294 271568 298350
rect 271248 298226 271568 298294
rect 271248 298170 271318 298226
rect 271374 298170 271442 298226
rect 271498 298170 271568 298226
rect 271248 298102 271568 298170
rect 271248 298046 271318 298102
rect 271374 298046 271442 298102
rect 271498 298046 271568 298102
rect 271248 297978 271568 298046
rect 271248 297922 271318 297978
rect 271374 297922 271442 297978
rect 271498 297922 271568 297978
rect 271248 297888 271568 297922
rect 301968 298350 302288 298384
rect 301968 298294 302038 298350
rect 302094 298294 302162 298350
rect 302218 298294 302288 298350
rect 301968 298226 302288 298294
rect 301968 298170 302038 298226
rect 302094 298170 302162 298226
rect 302218 298170 302288 298226
rect 301968 298102 302288 298170
rect 301968 298046 302038 298102
rect 302094 298046 302162 298102
rect 302218 298046 302288 298102
rect 301968 297978 302288 298046
rect 301968 297922 302038 297978
rect 302094 297922 302162 297978
rect 302218 297922 302288 297978
rect 301968 297888 302288 297922
rect 332688 298350 333008 298384
rect 332688 298294 332758 298350
rect 332814 298294 332882 298350
rect 332938 298294 333008 298350
rect 332688 298226 333008 298294
rect 332688 298170 332758 298226
rect 332814 298170 332882 298226
rect 332938 298170 333008 298226
rect 332688 298102 333008 298170
rect 332688 298046 332758 298102
rect 332814 298046 332882 298102
rect 332938 298046 333008 298102
rect 332688 297978 333008 298046
rect 332688 297922 332758 297978
rect 332814 297922 332882 297978
rect 332938 297922 333008 297978
rect 332688 297888 333008 297922
rect 225168 292350 225488 292384
rect 225168 292294 225238 292350
rect 225294 292294 225362 292350
rect 225418 292294 225488 292350
rect 225168 292226 225488 292294
rect 225168 292170 225238 292226
rect 225294 292170 225362 292226
rect 225418 292170 225488 292226
rect 225168 292102 225488 292170
rect 225168 292046 225238 292102
rect 225294 292046 225362 292102
rect 225418 292046 225488 292102
rect 225168 291978 225488 292046
rect 225168 291922 225238 291978
rect 225294 291922 225362 291978
rect 225418 291922 225488 291978
rect 225168 291888 225488 291922
rect 255888 292350 256208 292384
rect 255888 292294 255958 292350
rect 256014 292294 256082 292350
rect 256138 292294 256208 292350
rect 255888 292226 256208 292294
rect 255888 292170 255958 292226
rect 256014 292170 256082 292226
rect 256138 292170 256208 292226
rect 255888 292102 256208 292170
rect 255888 292046 255958 292102
rect 256014 292046 256082 292102
rect 256138 292046 256208 292102
rect 255888 291978 256208 292046
rect 255888 291922 255958 291978
rect 256014 291922 256082 291978
rect 256138 291922 256208 291978
rect 255888 291888 256208 291922
rect 286608 292350 286928 292384
rect 286608 292294 286678 292350
rect 286734 292294 286802 292350
rect 286858 292294 286928 292350
rect 286608 292226 286928 292294
rect 286608 292170 286678 292226
rect 286734 292170 286802 292226
rect 286858 292170 286928 292226
rect 286608 292102 286928 292170
rect 286608 292046 286678 292102
rect 286734 292046 286802 292102
rect 286858 292046 286928 292102
rect 286608 291978 286928 292046
rect 286608 291922 286678 291978
rect 286734 291922 286802 291978
rect 286858 291922 286928 291978
rect 286608 291888 286928 291922
rect 317328 292350 317648 292384
rect 317328 292294 317398 292350
rect 317454 292294 317522 292350
rect 317578 292294 317648 292350
rect 317328 292226 317648 292294
rect 317328 292170 317398 292226
rect 317454 292170 317522 292226
rect 317578 292170 317648 292226
rect 317328 292102 317648 292170
rect 317328 292046 317398 292102
rect 317454 292046 317522 292102
rect 317578 292046 317648 292102
rect 317328 291978 317648 292046
rect 317328 291922 317398 291978
rect 317454 291922 317522 291978
rect 317578 291922 317648 291978
rect 317328 291888 317648 291922
rect 209808 280350 210128 280384
rect 209808 280294 209878 280350
rect 209934 280294 210002 280350
rect 210058 280294 210128 280350
rect 209808 280226 210128 280294
rect 209808 280170 209878 280226
rect 209934 280170 210002 280226
rect 210058 280170 210128 280226
rect 209808 280102 210128 280170
rect 209808 280046 209878 280102
rect 209934 280046 210002 280102
rect 210058 280046 210128 280102
rect 209808 279978 210128 280046
rect 209808 279922 209878 279978
rect 209934 279922 210002 279978
rect 210058 279922 210128 279978
rect 209808 279888 210128 279922
rect 240528 280350 240848 280384
rect 240528 280294 240598 280350
rect 240654 280294 240722 280350
rect 240778 280294 240848 280350
rect 240528 280226 240848 280294
rect 240528 280170 240598 280226
rect 240654 280170 240722 280226
rect 240778 280170 240848 280226
rect 240528 280102 240848 280170
rect 240528 280046 240598 280102
rect 240654 280046 240722 280102
rect 240778 280046 240848 280102
rect 240528 279978 240848 280046
rect 240528 279922 240598 279978
rect 240654 279922 240722 279978
rect 240778 279922 240848 279978
rect 240528 279888 240848 279922
rect 271248 280350 271568 280384
rect 271248 280294 271318 280350
rect 271374 280294 271442 280350
rect 271498 280294 271568 280350
rect 271248 280226 271568 280294
rect 271248 280170 271318 280226
rect 271374 280170 271442 280226
rect 271498 280170 271568 280226
rect 271248 280102 271568 280170
rect 271248 280046 271318 280102
rect 271374 280046 271442 280102
rect 271498 280046 271568 280102
rect 271248 279978 271568 280046
rect 271248 279922 271318 279978
rect 271374 279922 271442 279978
rect 271498 279922 271568 279978
rect 271248 279888 271568 279922
rect 301968 280350 302288 280384
rect 301968 280294 302038 280350
rect 302094 280294 302162 280350
rect 302218 280294 302288 280350
rect 301968 280226 302288 280294
rect 301968 280170 302038 280226
rect 302094 280170 302162 280226
rect 302218 280170 302288 280226
rect 301968 280102 302288 280170
rect 301968 280046 302038 280102
rect 302094 280046 302162 280102
rect 302218 280046 302288 280102
rect 301968 279978 302288 280046
rect 301968 279922 302038 279978
rect 302094 279922 302162 279978
rect 302218 279922 302288 279978
rect 301968 279888 302288 279922
rect 332688 280350 333008 280384
rect 332688 280294 332758 280350
rect 332814 280294 332882 280350
rect 332938 280294 333008 280350
rect 332688 280226 333008 280294
rect 332688 280170 332758 280226
rect 332814 280170 332882 280226
rect 332938 280170 333008 280226
rect 332688 280102 333008 280170
rect 332688 280046 332758 280102
rect 332814 280046 332882 280102
rect 332938 280046 333008 280102
rect 332688 279978 333008 280046
rect 332688 279922 332758 279978
rect 332814 279922 332882 279978
rect 332938 279922 333008 279978
rect 332688 279888 333008 279922
rect 225168 274350 225488 274384
rect 225168 274294 225238 274350
rect 225294 274294 225362 274350
rect 225418 274294 225488 274350
rect 225168 274226 225488 274294
rect 225168 274170 225238 274226
rect 225294 274170 225362 274226
rect 225418 274170 225488 274226
rect 225168 274102 225488 274170
rect 225168 274046 225238 274102
rect 225294 274046 225362 274102
rect 225418 274046 225488 274102
rect 225168 273978 225488 274046
rect 225168 273922 225238 273978
rect 225294 273922 225362 273978
rect 225418 273922 225488 273978
rect 225168 273888 225488 273922
rect 255888 274350 256208 274384
rect 255888 274294 255958 274350
rect 256014 274294 256082 274350
rect 256138 274294 256208 274350
rect 255888 274226 256208 274294
rect 255888 274170 255958 274226
rect 256014 274170 256082 274226
rect 256138 274170 256208 274226
rect 255888 274102 256208 274170
rect 255888 274046 255958 274102
rect 256014 274046 256082 274102
rect 256138 274046 256208 274102
rect 255888 273978 256208 274046
rect 255888 273922 255958 273978
rect 256014 273922 256082 273978
rect 256138 273922 256208 273978
rect 255888 273888 256208 273922
rect 286608 274350 286928 274384
rect 286608 274294 286678 274350
rect 286734 274294 286802 274350
rect 286858 274294 286928 274350
rect 286608 274226 286928 274294
rect 286608 274170 286678 274226
rect 286734 274170 286802 274226
rect 286858 274170 286928 274226
rect 286608 274102 286928 274170
rect 286608 274046 286678 274102
rect 286734 274046 286802 274102
rect 286858 274046 286928 274102
rect 286608 273978 286928 274046
rect 286608 273922 286678 273978
rect 286734 273922 286802 273978
rect 286858 273922 286928 273978
rect 286608 273888 286928 273922
rect 317328 274350 317648 274384
rect 317328 274294 317398 274350
rect 317454 274294 317522 274350
rect 317578 274294 317648 274350
rect 317328 274226 317648 274294
rect 317328 274170 317398 274226
rect 317454 274170 317522 274226
rect 317578 274170 317648 274226
rect 317328 274102 317648 274170
rect 317328 274046 317398 274102
rect 317454 274046 317522 274102
rect 317578 274046 317648 274102
rect 317328 273978 317648 274046
rect 317328 273922 317398 273978
rect 317454 273922 317522 273978
rect 317578 273922 317648 273978
rect 317328 273888 317648 273922
rect 209808 262350 210128 262384
rect 209808 262294 209878 262350
rect 209934 262294 210002 262350
rect 210058 262294 210128 262350
rect 209808 262226 210128 262294
rect 209808 262170 209878 262226
rect 209934 262170 210002 262226
rect 210058 262170 210128 262226
rect 209808 262102 210128 262170
rect 209808 262046 209878 262102
rect 209934 262046 210002 262102
rect 210058 262046 210128 262102
rect 209808 261978 210128 262046
rect 209808 261922 209878 261978
rect 209934 261922 210002 261978
rect 210058 261922 210128 261978
rect 209808 261888 210128 261922
rect 240528 262350 240848 262384
rect 240528 262294 240598 262350
rect 240654 262294 240722 262350
rect 240778 262294 240848 262350
rect 240528 262226 240848 262294
rect 240528 262170 240598 262226
rect 240654 262170 240722 262226
rect 240778 262170 240848 262226
rect 240528 262102 240848 262170
rect 240528 262046 240598 262102
rect 240654 262046 240722 262102
rect 240778 262046 240848 262102
rect 240528 261978 240848 262046
rect 240528 261922 240598 261978
rect 240654 261922 240722 261978
rect 240778 261922 240848 261978
rect 240528 261888 240848 261922
rect 271248 262350 271568 262384
rect 271248 262294 271318 262350
rect 271374 262294 271442 262350
rect 271498 262294 271568 262350
rect 271248 262226 271568 262294
rect 271248 262170 271318 262226
rect 271374 262170 271442 262226
rect 271498 262170 271568 262226
rect 271248 262102 271568 262170
rect 271248 262046 271318 262102
rect 271374 262046 271442 262102
rect 271498 262046 271568 262102
rect 271248 261978 271568 262046
rect 271248 261922 271318 261978
rect 271374 261922 271442 261978
rect 271498 261922 271568 261978
rect 271248 261888 271568 261922
rect 301968 262350 302288 262384
rect 301968 262294 302038 262350
rect 302094 262294 302162 262350
rect 302218 262294 302288 262350
rect 301968 262226 302288 262294
rect 301968 262170 302038 262226
rect 302094 262170 302162 262226
rect 302218 262170 302288 262226
rect 301968 262102 302288 262170
rect 301968 262046 302038 262102
rect 302094 262046 302162 262102
rect 302218 262046 302288 262102
rect 301968 261978 302288 262046
rect 301968 261922 302038 261978
rect 302094 261922 302162 261978
rect 302218 261922 302288 261978
rect 301968 261888 302288 261922
rect 332688 262350 333008 262384
rect 332688 262294 332758 262350
rect 332814 262294 332882 262350
rect 332938 262294 333008 262350
rect 332688 262226 333008 262294
rect 332688 262170 332758 262226
rect 332814 262170 332882 262226
rect 332938 262170 333008 262226
rect 332688 262102 333008 262170
rect 332688 262046 332758 262102
rect 332814 262046 332882 262102
rect 332938 262046 333008 262102
rect 332688 261978 333008 262046
rect 332688 261922 332758 261978
rect 332814 261922 332882 261978
rect 332938 261922 333008 261978
rect 332688 261888 333008 261922
rect 225168 256350 225488 256384
rect 225168 256294 225238 256350
rect 225294 256294 225362 256350
rect 225418 256294 225488 256350
rect 225168 256226 225488 256294
rect 225168 256170 225238 256226
rect 225294 256170 225362 256226
rect 225418 256170 225488 256226
rect 225168 256102 225488 256170
rect 225168 256046 225238 256102
rect 225294 256046 225362 256102
rect 225418 256046 225488 256102
rect 225168 255978 225488 256046
rect 225168 255922 225238 255978
rect 225294 255922 225362 255978
rect 225418 255922 225488 255978
rect 225168 255888 225488 255922
rect 255888 256350 256208 256384
rect 255888 256294 255958 256350
rect 256014 256294 256082 256350
rect 256138 256294 256208 256350
rect 255888 256226 256208 256294
rect 255888 256170 255958 256226
rect 256014 256170 256082 256226
rect 256138 256170 256208 256226
rect 255888 256102 256208 256170
rect 255888 256046 255958 256102
rect 256014 256046 256082 256102
rect 256138 256046 256208 256102
rect 255888 255978 256208 256046
rect 255888 255922 255958 255978
rect 256014 255922 256082 255978
rect 256138 255922 256208 255978
rect 255888 255888 256208 255922
rect 286608 256350 286928 256384
rect 286608 256294 286678 256350
rect 286734 256294 286802 256350
rect 286858 256294 286928 256350
rect 286608 256226 286928 256294
rect 286608 256170 286678 256226
rect 286734 256170 286802 256226
rect 286858 256170 286928 256226
rect 286608 256102 286928 256170
rect 286608 256046 286678 256102
rect 286734 256046 286802 256102
rect 286858 256046 286928 256102
rect 286608 255978 286928 256046
rect 286608 255922 286678 255978
rect 286734 255922 286802 255978
rect 286858 255922 286928 255978
rect 286608 255888 286928 255922
rect 317328 256350 317648 256384
rect 317328 256294 317398 256350
rect 317454 256294 317522 256350
rect 317578 256294 317648 256350
rect 317328 256226 317648 256294
rect 317328 256170 317398 256226
rect 317454 256170 317522 256226
rect 317578 256170 317648 256226
rect 317328 256102 317648 256170
rect 317328 256046 317398 256102
rect 317454 256046 317522 256102
rect 317578 256046 317648 256102
rect 317328 255978 317648 256046
rect 317328 255922 317398 255978
rect 317454 255922 317522 255978
rect 317578 255922 317648 255978
rect 317328 255888 317648 255922
rect 335804 253558 335860 253568
rect 209808 244350 210128 244384
rect 209808 244294 209878 244350
rect 209934 244294 210002 244350
rect 210058 244294 210128 244350
rect 209808 244226 210128 244294
rect 209808 244170 209878 244226
rect 209934 244170 210002 244226
rect 210058 244170 210128 244226
rect 209808 244102 210128 244170
rect 209808 244046 209878 244102
rect 209934 244046 210002 244102
rect 210058 244046 210128 244102
rect 209808 243978 210128 244046
rect 209808 243922 209878 243978
rect 209934 243922 210002 243978
rect 210058 243922 210128 243978
rect 209808 243888 210128 243922
rect 240528 244350 240848 244384
rect 240528 244294 240598 244350
rect 240654 244294 240722 244350
rect 240778 244294 240848 244350
rect 240528 244226 240848 244294
rect 240528 244170 240598 244226
rect 240654 244170 240722 244226
rect 240778 244170 240848 244226
rect 240528 244102 240848 244170
rect 240528 244046 240598 244102
rect 240654 244046 240722 244102
rect 240778 244046 240848 244102
rect 240528 243978 240848 244046
rect 240528 243922 240598 243978
rect 240654 243922 240722 243978
rect 240778 243922 240848 243978
rect 240528 243888 240848 243922
rect 271248 244350 271568 244384
rect 271248 244294 271318 244350
rect 271374 244294 271442 244350
rect 271498 244294 271568 244350
rect 271248 244226 271568 244294
rect 271248 244170 271318 244226
rect 271374 244170 271442 244226
rect 271498 244170 271568 244226
rect 271248 244102 271568 244170
rect 271248 244046 271318 244102
rect 271374 244046 271442 244102
rect 271498 244046 271568 244102
rect 271248 243978 271568 244046
rect 271248 243922 271318 243978
rect 271374 243922 271442 243978
rect 271498 243922 271568 243978
rect 271248 243888 271568 243922
rect 301968 244350 302288 244384
rect 301968 244294 302038 244350
rect 302094 244294 302162 244350
rect 302218 244294 302288 244350
rect 301968 244226 302288 244294
rect 301968 244170 302038 244226
rect 302094 244170 302162 244226
rect 302218 244170 302288 244226
rect 301968 244102 302288 244170
rect 301968 244046 302038 244102
rect 302094 244046 302162 244102
rect 302218 244046 302288 244102
rect 301968 243978 302288 244046
rect 301968 243922 302038 243978
rect 302094 243922 302162 243978
rect 302218 243922 302288 243978
rect 301968 243888 302288 243922
rect 332688 244350 333008 244384
rect 332688 244294 332758 244350
rect 332814 244294 332882 244350
rect 332938 244294 333008 244350
rect 332688 244226 333008 244294
rect 332688 244170 332758 244226
rect 332814 244170 332882 244226
rect 332938 244170 333008 244226
rect 332688 244102 333008 244170
rect 332688 244046 332758 244102
rect 332814 244046 332882 244102
rect 332938 244046 333008 244102
rect 332688 243978 333008 244046
rect 332688 243922 332758 243978
rect 332814 243922 332882 243978
rect 332938 243922 333008 243978
rect 332688 243888 333008 243922
rect 323260 242758 323316 242768
rect 278012 242038 278068 242048
rect 273868 241332 273924 241342
rect 220458 238350 221078 241154
rect 220458 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 221078 238350
rect 220458 238226 221078 238294
rect 220458 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 221078 238226
rect 220458 238102 221078 238170
rect 220458 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 221078 238102
rect 220458 237978 221078 238046
rect 220458 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 221078 237978
rect 219996 237076 220052 237086
rect 218316 236964 218372 236974
rect 218316 231238 218372 236908
rect 219996 231418 220052 237020
rect 219996 231352 220052 231362
rect 218316 231172 218372 231182
rect 199724 216178 199780 216188
rect 220458 220350 221078 237922
rect 241948 238532 242004 238542
rect 233212 237300 233268 237310
rect 228508 236964 228564 236974
rect 228508 231058 228564 236908
rect 233212 234478 233268 237244
rect 233212 234412 233268 234422
rect 235900 237300 235956 237310
rect 235900 234478 235956 237244
rect 241948 236998 242004 238476
rect 242620 238532 242676 238542
rect 242620 237178 242676 238476
rect 242620 237112 242676 237122
rect 251178 238350 251798 241154
rect 272748 239316 272804 239326
rect 251178 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 251798 238350
rect 251178 238226 251798 238294
rect 251178 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 251798 238226
rect 251178 238102 251798 238170
rect 251178 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 251798 238102
rect 251178 237978 251798 238046
rect 251178 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 251798 237978
rect 235900 234412 235956 234422
rect 236796 236964 236852 236974
rect 241948 236932 242004 236942
rect 228508 230992 228564 231002
rect 236796 227818 236852 236908
rect 236796 227752 236852 227762
rect 220458 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 221078 220350
rect 220458 220226 221078 220294
rect 220458 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 221078 220226
rect 220458 220102 221078 220170
rect 220458 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 221078 220102
rect 220458 219978 221078 220046
rect 220458 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 221078 219978
rect 199388 214610 199444 214620
rect 199276 211192 199332 211202
rect 197820 210832 197876 210842
rect 220458 210462 221078 219922
rect 251178 220350 251798 237922
rect 267260 238420 267316 238430
rect 251178 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 251798 220350
rect 251178 220226 251798 220294
rect 251178 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 251798 220226
rect 251178 220102 251798 220170
rect 251178 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 251798 220102
rect 251178 219978 251798 220046
rect 251178 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 251798 219978
rect 251178 210462 251798 219922
rect 266812 235060 266868 235070
rect 190428 209794 190484 209804
rect 185836 209682 185892 209692
rect 181356 209346 181412 209356
rect 75168 202350 75488 202384
rect 75168 202294 75238 202350
rect 75294 202294 75362 202350
rect 75418 202294 75488 202350
rect 75168 202226 75488 202294
rect 75168 202170 75238 202226
rect 75294 202170 75362 202226
rect 75418 202170 75488 202226
rect 75168 202102 75488 202170
rect 75168 202046 75238 202102
rect 75294 202046 75362 202102
rect 75418 202046 75488 202102
rect 75168 201978 75488 202046
rect 75168 201922 75238 201978
rect 75294 201922 75362 201978
rect 75418 201922 75488 201978
rect 75168 201888 75488 201922
rect 105888 202350 106208 202384
rect 105888 202294 105958 202350
rect 106014 202294 106082 202350
rect 106138 202294 106208 202350
rect 105888 202226 106208 202294
rect 105888 202170 105958 202226
rect 106014 202170 106082 202226
rect 106138 202170 106208 202226
rect 105888 202102 106208 202170
rect 105888 202046 105958 202102
rect 106014 202046 106082 202102
rect 106138 202046 106208 202102
rect 105888 201978 106208 202046
rect 105888 201922 105958 201978
rect 106014 201922 106082 201978
rect 106138 201922 106208 201978
rect 105888 201888 106208 201922
rect 136608 202350 136928 202384
rect 136608 202294 136678 202350
rect 136734 202294 136802 202350
rect 136858 202294 136928 202350
rect 136608 202226 136928 202294
rect 136608 202170 136678 202226
rect 136734 202170 136802 202226
rect 136858 202170 136928 202226
rect 136608 202102 136928 202170
rect 136608 202046 136678 202102
rect 136734 202046 136802 202102
rect 136858 202046 136928 202102
rect 136608 201978 136928 202046
rect 136608 201922 136678 201978
rect 136734 201922 136802 201978
rect 136858 201922 136928 201978
rect 136608 201888 136928 201922
rect 167328 202350 167648 202384
rect 167328 202294 167398 202350
rect 167454 202294 167522 202350
rect 167578 202294 167648 202350
rect 167328 202226 167648 202294
rect 167328 202170 167398 202226
rect 167454 202170 167522 202226
rect 167578 202170 167648 202226
rect 167328 202102 167648 202170
rect 167328 202046 167398 202102
rect 167454 202046 167522 202102
rect 167578 202046 167648 202102
rect 167328 201978 167648 202046
rect 167328 201922 167398 201978
rect 167454 201922 167522 201978
rect 167578 201922 167648 201978
rect 167328 201888 167648 201922
rect 198048 202350 198368 202384
rect 198048 202294 198118 202350
rect 198174 202294 198242 202350
rect 198298 202294 198368 202350
rect 198048 202226 198368 202294
rect 198048 202170 198118 202226
rect 198174 202170 198242 202226
rect 198298 202170 198368 202226
rect 198048 202102 198368 202170
rect 198048 202046 198118 202102
rect 198174 202046 198242 202102
rect 198298 202046 198368 202102
rect 198048 201978 198368 202046
rect 198048 201922 198118 201978
rect 198174 201922 198242 201978
rect 198298 201922 198368 201978
rect 198048 201888 198368 201922
rect 228768 202350 229088 202384
rect 228768 202294 228838 202350
rect 228894 202294 228962 202350
rect 229018 202294 229088 202350
rect 228768 202226 229088 202294
rect 228768 202170 228838 202226
rect 228894 202170 228962 202226
rect 229018 202170 229088 202226
rect 228768 202102 229088 202170
rect 228768 202046 228838 202102
rect 228894 202046 228962 202102
rect 229018 202046 229088 202102
rect 228768 201978 229088 202046
rect 228768 201922 228838 201978
rect 228894 201922 228962 201978
rect 229018 201922 229088 201978
rect 228768 201888 229088 201922
rect 259488 202350 259808 202384
rect 259488 202294 259558 202350
rect 259614 202294 259682 202350
rect 259738 202294 259808 202350
rect 259488 202226 259808 202294
rect 259488 202170 259558 202226
rect 259614 202170 259682 202226
rect 259738 202170 259808 202226
rect 259488 202102 259808 202170
rect 259488 202046 259558 202102
rect 259614 202046 259682 202102
rect 259738 202046 259808 202102
rect 259488 201978 259808 202046
rect 259488 201922 259558 201978
rect 259614 201922 259682 201978
rect 259738 201922 259808 201978
rect 259488 201888 259808 201922
rect 59808 190350 60128 190384
rect 59808 190294 59878 190350
rect 59934 190294 60002 190350
rect 60058 190294 60128 190350
rect 59808 190226 60128 190294
rect 59808 190170 59878 190226
rect 59934 190170 60002 190226
rect 60058 190170 60128 190226
rect 59808 190102 60128 190170
rect 59808 190046 59878 190102
rect 59934 190046 60002 190102
rect 60058 190046 60128 190102
rect 59808 189978 60128 190046
rect 59808 189922 59878 189978
rect 59934 189922 60002 189978
rect 60058 189922 60128 189978
rect 59808 189888 60128 189922
rect 90528 190350 90848 190384
rect 90528 190294 90598 190350
rect 90654 190294 90722 190350
rect 90778 190294 90848 190350
rect 90528 190226 90848 190294
rect 90528 190170 90598 190226
rect 90654 190170 90722 190226
rect 90778 190170 90848 190226
rect 90528 190102 90848 190170
rect 90528 190046 90598 190102
rect 90654 190046 90722 190102
rect 90778 190046 90848 190102
rect 90528 189978 90848 190046
rect 90528 189922 90598 189978
rect 90654 189922 90722 189978
rect 90778 189922 90848 189978
rect 90528 189888 90848 189922
rect 121248 190350 121568 190384
rect 121248 190294 121318 190350
rect 121374 190294 121442 190350
rect 121498 190294 121568 190350
rect 121248 190226 121568 190294
rect 121248 190170 121318 190226
rect 121374 190170 121442 190226
rect 121498 190170 121568 190226
rect 121248 190102 121568 190170
rect 121248 190046 121318 190102
rect 121374 190046 121442 190102
rect 121498 190046 121568 190102
rect 121248 189978 121568 190046
rect 121248 189922 121318 189978
rect 121374 189922 121442 189978
rect 121498 189922 121568 189978
rect 121248 189888 121568 189922
rect 151968 190350 152288 190384
rect 151968 190294 152038 190350
rect 152094 190294 152162 190350
rect 152218 190294 152288 190350
rect 151968 190226 152288 190294
rect 151968 190170 152038 190226
rect 152094 190170 152162 190226
rect 152218 190170 152288 190226
rect 151968 190102 152288 190170
rect 151968 190046 152038 190102
rect 152094 190046 152162 190102
rect 152218 190046 152288 190102
rect 151968 189978 152288 190046
rect 151968 189922 152038 189978
rect 152094 189922 152162 189978
rect 152218 189922 152288 189978
rect 151968 189888 152288 189922
rect 182688 190350 183008 190384
rect 182688 190294 182758 190350
rect 182814 190294 182882 190350
rect 182938 190294 183008 190350
rect 182688 190226 183008 190294
rect 182688 190170 182758 190226
rect 182814 190170 182882 190226
rect 182938 190170 183008 190226
rect 182688 190102 183008 190170
rect 182688 190046 182758 190102
rect 182814 190046 182882 190102
rect 182938 190046 183008 190102
rect 182688 189978 183008 190046
rect 182688 189922 182758 189978
rect 182814 189922 182882 189978
rect 182938 189922 183008 189978
rect 182688 189888 183008 189922
rect 213408 190350 213728 190384
rect 213408 190294 213478 190350
rect 213534 190294 213602 190350
rect 213658 190294 213728 190350
rect 213408 190226 213728 190294
rect 213408 190170 213478 190226
rect 213534 190170 213602 190226
rect 213658 190170 213728 190226
rect 213408 190102 213728 190170
rect 213408 190046 213478 190102
rect 213534 190046 213602 190102
rect 213658 190046 213728 190102
rect 213408 189978 213728 190046
rect 213408 189922 213478 189978
rect 213534 189922 213602 189978
rect 213658 189922 213728 189978
rect 213408 189888 213728 189922
rect 244128 190350 244448 190384
rect 244128 190294 244198 190350
rect 244254 190294 244322 190350
rect 244378 190294 244448 190350
rect 244128 190226 244448 190294
rect 244128 190170 244198 190226
rect 244254 190170 244322 190226
rect 244378 190170 244448 190226
rect 244128 190102 244448 190170
rect 244128 190046 244198 190102
rect 244254 190046 244322 190102
rect 244378 190046 244448 190102
rect 244128 189978 244448 190046
rect 244128 189922 244198 189978
rect 244254 189922 244322 189978
rect 244378 189922 244448 189978
rect 244128 189888 244448 189922
rect 75168 184350 75488 184384
rect 75168 184294 75238 184350
rect 75294 184294 75362 184350
rect 75418 184294 75488 184350
rect 75168 184226 75488 184294
rect 75168 184170 75238 184226
rect 75294 184170 75362 184226
rect 75418 184170 75488 184226
rect 75168 184102 75488 184170
rect 75168 184046 75238 184102
rect 75294 184046 75362 184102
rect 75418 184046 75488 184102
rect 75168 183978 75488 184046
rect 75168 183922 75238 183978
rect 75294 183922 75362 183978
rect 75418 183922 75488 183978
rect 75168 183888 75488 183922
rect 105888 184350 106208 184384
rect 105888 184294 105958 184350
rect 106014 184294 106082 184350
rect 106138 184294 106208 184350
rect 105888 184226 106208 184294
rect 105888 184170 105958 184226
rect 106014 184170 106082 184226
rect 106138 184170 106208 184226
rect 105888 184102 106208 184170
rect 105888 184046 105958 184102
rect 106014 184046 106082 184102
rect 106138 184046 106208 184102
rect 105888 183978 106208 184046
rect 105888 183922 105958 183978
rect 106014 183922 106082 183978
rect 106138 183922 106208 183978
rect 105888 183888 106208 183922
rect 136608 184350 136928 184384
rect 136608 184294 136678 184350
rect 136734 184294 136802 184350
rect 136858 184294 136928 184350
rect 136608 184226 136928 184294
rect 136608 184170 136678 184226
rect 136734 184170 136802 184226
rect 136858 184170 136928 184226
rect 136608 184102 136928 184170
rect 136608 184046 136678 184102
rect 136734 184046 136802 184102
rect 136858 184046 136928 184102
rect 136608 183978 136928 184046
rect 136608 183922 136678 183978
rect 136734 183922 136802 183978
rect 136858 183922 136928 183978
rect 136608 183888 136928 183922
rect 167328 184350 167648 184384
rect 167328 184294 167398 184350
rect 167454 184294 167522 184350
rect 167578 184294 167648 184350
rect 167328 184226 167648 184294
rect 167328 184170 167398 184226
rect 167454 184170 167522 184226
rect 167578 184170 167648 184226
rect 167328 184102 167648 184170
rect 167328 184046 167398 184102
rect 167454 184046 167522 184102
rect 167578 184046 167648 184102
rect 167328 183978 167648 184046
rect 167328 183922 167398 183978
rect 167454 183922 167522 183978
rect 167578 183922 167648 183978
rect 167328 183888 167648 183922
rect 198048 184350 198368 184384
rect 198048 184294 198118 184350
rect 198174 184294 198242 184350
rect 198298 184294 198368 184350
rect 198048 184226 198368 184294
rect 198048 184170 198118 184226
rect 198174 184170 198242 184226
rect 198298 184170 198368 184226
rect 198048 184102 198368 184170
rect 198048 184046 198118 184102
rect 198174 184046 198242 184102
rect 198298 184046 198368 184102
rect 198048 183978 198368 184046
rect 198048 183922 198118 183978
rect 198174 183922 198242 183978
rect 198298 183922 198368 183978
rect 198048 183888 198368 183922
rect 228768 184350 229088 184384
rect 228768 184294 228838 184350
rect 228894 184294 228962 184350
rect 229018 184294 229088 184350
rect 228768 184226 229088 184294
rect 228768 184170 228838 184226
rect 228894 184170 228962 184226
rect 229018 184170 229088 184226
rect 228768 184102 229088 184170
rect 228768 184046 228838 184102
rect 228894 184046 228962 184102
rect 229018 184046 229088 184102
rect 228768 183978 229088 184046
rect 228768 183922 228838 183978
rect 228894 183922 228962 183978
rect 229018 183922 229088 183978
rect 228768 183888 229088 183922
rect 259488 184350 259808 184384
rect 259488 184294 259558 184350
rect 259614 184294 259682 184350
rect 259738 184294 259808 184350
rect 259488 184226 259808 184294
rect 259488 184170 259558 184226
rect 259614 184170 259682 184226
rect 259738 184170 259808 184226
rect 259488 184102 259808 184170
rect 259488 184046 259558 184102
rect 259614 184046 259682 184102
rect 259738 184046 259808 184102
rect 259488 183978 259808 184046
rect 259488 183922 259558 183978
rect 259614 183922 259682 183978
rect 259738 183922 259808 183978
rect 259488 183888 259808 183922
rect 59808 172350 60128 172384
rect 59808 172294 59878 172350
rect 59934 172294 60002 172350
rect 60058 172294 60128 172350
rect 59808 172226 60128 172294
rect 59808 172170 59878 172226
rect 59934 172170 60002 172226
rect 60058 172170 60128 172226
rect 59808 172102 60128 172170
rect 59808 172046 59878 172102
rect 59934 172046 60002 172102
rect 60058 172046 60128 172102
rect 59808 171978 60128 172046
rect 59808 171922 59878 171978
rect 59934 171922 60002 171978
rect 60058 171922 60128 171978
rect 59808 171888 60128 171922
rect 90528 172350 90848 172384
rect 90528 172294 90598 172350
rect 90654 172294 90722 172350
rect 90778 172294 90848 172350
rect 90528 172226 90848 172294
rect 90528 172170 90598 172226
rect 90654 172170 90722 172226
rect 90778 172170 90848 172226
rect 90528 172102 90848 172170
rect 90528 172046 90598 172102
rect 90654 172046 90722 172102
rect 90778 172046 90848 172102
rect 90528 171978 90848 172046
rect 90528 171922 90598 171978
rect 90654 171922 90722 171978
rect 90778 171922 90848 171978
rect 90528 171888 90848 171922
rect 121248 172350 121568 172384
rect 121248 172294 121318 172350
rect 121374 172294 121442 172350
rect 121498 172294 121568 172350
rect 121248 172226 121568 172294
rect 121248 172170 121318 172226
rect 121374 172170 121442 172226
rect 121498 172170 121568 172226
rect 121248 172102 121568 172170
rect 121248 172046 121318 172102
rect 121374 172046 121442 172102
rect 121498 172046 121568 172102
rect 121248 171978 121568 172046
rect 121248 171922 121318 171978
rect 121374 171922 121442 171978
rect 121498 171922 121568 171978
rect 121248 171888 121568 171922
rect 151968 172350 152288 172384
rect 151968 172294 152038 172350
rect 152094 172294 152162 172350
rect 152218 172294 152288 172350
rect 151968 172226 152288 172294
rect 151968 172170 152038 172226
rect 152094 172170 152162 172226
rect 152218 172170 152288 172226
rect 151968 172102 152288 172170
rect 151968 172046 152038 172102
rect 152094 172046 152162 172102
rect 152218 172046 152288 172102
rect 151968 171978 152288 172046
rect 151968 171922 152038 171978
rect 152094 171922 152162 171978
rect 152218 171922 152288 171978
rect 151968 171888 152288 171922
rect 182688 172350 183008 172384
rect 182688 172294 182758 172350
rect 182814 172294 182882 172350
rect 182938 172294 183008 172350
rect 182688 172226 183008 172294
rect 182688 172170 182758 172226
rect 182814 172170 182882 172226
rect 182938 172170 183008 172226
rect 182688 172102 183008 172170
rect 182688 172046 182758 172102
rect 182814 172046 182882 172102
rect 182938 172046 183008 172102
rect 182688 171978 183008 172046
rect 182688 171922 182758 171978
rect 182814 171922 182882 171978
rect 182938 171922 183008 171978
rect 182688 171888 183008 171922
rect 213408 172350 213728 172384
rect 213408 172294 213478 172350
rect 213534 172294 213602 172350
rect 213658 172294 213728 172350
rect 213408 172226 213728 172294
rect 213408 172170 213478 172226
rect 213534 172170 213602 172226
rect 213658 172170 213728 172226
rect 213408 172102 213728 172170
rect 213408 172046 213478 172102
rect 213534 172046 213602 172102
rect 213658 172046 213728 172102
rect 213408 171978 213728 172046
rect 213408 171922 213478 171978
rect 213534 171922 213602 171978
rect 213658 171922 213728 171978
rect 213408 171888 213728 171922
rect 244128 172350 244448 172384
rect 244128 172294 244198 172350
rect 244254 172294 244322 172350
rect 244378 172294 244448 172350
rect 244128 172226 244448 172294
rect 244128 172170 244198 172226
rect 244254 172170 244322 172226
rect 244378 172170 244448 172226
rect 244128 172102 244448 172170
rect 244128 172046 244198 172102
rect 244254 172046 244322 172102
rect 244378 172046 244448 172102
rect 244128 171978 244448 172046
rect 244128 171922 244198 171978
rect 244254 171922 244322 171978
rect 244378 171922 244448 171978
rect 244128 171888 244448 171922
rect 75168 166350 75488 166384
rect 75168 166294 75238 166350
rect 75294 166294 75362 166350
rect 75418 166294 75488 166350
rect 75168 166226 75488 166294
rect 75168 166170 75238 166226
rect 75294 166170 75362 166226
rect 75418 166170 75488 166226
rect 75168 166102 75488 166170
rect 75168 166046 75238 166102
rect 75294 166046 75362 166102
rect 75418 166046 75488 166102
rect 75168 165978 75488 166046
rect 75168 165922 75238 165978
rect 75294 165922 75362 165978
rect 75418 165922 75488 165978
rect 75168 165888 75488 165922
rect 105888 166350 106208 166384
rect 105888 166294 105958 166350
rect 106014 166294 106082 166350
rect 106138 166294 106208 166350
rect 105888 166226 106208 166294
rect 105888 166170 105958 166226
rect 106014 166170 106082 166226
rect 106138 166170 106208 166226
rect 105888 166102 106208 166170
rect 105888 166046 105958 166102
rect 106014 166046 106082 166102
rect 106138 166046 106208 166102
rect 105888 165978 106208 166046
rect 105888 165922 105958 165978
rect 106014 165922 106082 165978
rect 106138 165922 106208 165978
rect 105888 165888 106208 165922
rect 136608 166350 136928 166384
rect 136608 166294 136678 166350
rect 136734 166294 136802 166350
rect 136858 166294 136928 166350
rect 136608 166226 136928 166294
rect 136608 166170 136678 166226
rect 136734 166170 136802 166226
rect 136858 166170 136928 166226
rect 136608 166102 136928 166170
rect 136608 166046 136678 166102
rect 136734 166046 136802 166102
rect 136858 166046 136928 166102
rect 136608 165978 136928 166046
rect 136608 165922 136678 165978
rect 136734 165922 136802 165978
rect 136858 165922 136928 165978
rect 136608 165888 136928 165922
rect 167328 166350 167648 166384
rect 167328 166294 167398 166350
rect 167454 166294 167522 166350
rect 167578 166294 167648 166350
rect 167328 166226 167648 166294
rect 167328 166170 167398 166226
rect 167454 166170 167522 166226
rect 167578 166170 167648 166226
rect 167328 166102 167648 166170
rect 167328 166046 167398 166102
rect 167454 166046 167522 166102
rect 167578 166046 167648 166102
rect 167328 165978 167648 166046
rect 167328 165922 167398 165978
rect 167454 165922 167522 165978
rect 167578 165922 167648 165978
rect 167328 165888 167648 165922
rect 198048 166350 198368 166384
rect 198048 166294 198118 166350
rect 198174 166294 198242 166350
rect 198298 166294 198368 166350
rect 198048 166226 198368 166294
rect 198048 166170 198118 166226
rect 198174 166170 198242 166226
rect 198298 166170 198368 166226
rect 198048 166102 198368 166170
rect 198048 166046 198118 166102
rect 198174 166046 198242 166102
rect 198298 166046 198368 166102
rect 198048 165978 198368 166046
rect 198048 165922 198118 165978
rect 198174 165922 198242 165978
rect 198298 165922 198368 165978
rect 198048 165888 198368 165922
rect 228768 166350 229088 166384
rect 228768 166294 228838 166350
rect 228894 166294 228962 166350
rect 229018 166294 229088 166350
rect 228768 166226 229088 166294
rect 228768 166170 228838 166226
rect 228894 166170 228962 166226
rect 229018 166170 229088 166226
rect 228768 166102 229088 166170
rect 228768 166046 228838 166102
rect 228894 166046 228962 166102
rect 229018 166046 229088 166102
rect 228768 165978 229088 166046
rect 228768 165922 228838 165978
rect 228894 165922 228962 165978
rect 229018 165922 229088 165978
rect 228768 165888 229088 165922
rect 259488 166350 259808 166384
rect 259488 166294 259558 166350
rect 259614 166294 259682 166350
rect 259738 166294 259808 166350
rect 259488 166226 259808 166294
rect 259488 166170 259558 166226
rect 259614 166170 259682 166226
rect 259738 166170 259808 166226
rect 259488 166102 259808 166170
rect 259488 166046 259558 166102
rect 259614 166046 259682 166102
rect 259738 166046 259808 166102
rect 259488 165978 259808 166046
rect 259488 165922 259558 165978
rect 259614 165922 259682 165978
rect 259738 165922 259808 165978
rect 259488 165888 259808 165922
rect 59808 154350 60128 154384
rect 59808 154294 59878 154350
rect 59934 154294 60002 154350
rect 60058 154294 60128 154350
rect 59808 154226 60128 154294
rect 59808 154170 59878 154226
rect 59934 154170 60002 154226
rect 60058 154170 60128 154226
rect 59808 154102 60128 154170
rect 59808 154046 59878 154102
rect 59934 154046 60002 154102
rect 60058 154046 60128 154102
rect 59808 153978 60128 154046
rect 59808 153922 59878 153978
rect 59934 153922 60002 153978
rect 60058 153922 60128 153978
rect 59808 153888 60128 153922
rect 90528 154350 90848 154384
rect 90528 154294 90598 154350
rect 90654 154294 90722 154350
rect 90778 154294 90848 154350
rect 90528 154226 90848 154294
rect 90528 154170 90598 154226
rect 90654 154170 90722 154226
rect 90778 154170 90848 154226
rect 90528 154102 90848 154170
rect 90528 154046 90598 154102
rect 90654 154046 90722 154102
rect 90778 154046 90848 154102
rect 90528 153978 90848 154046
rect 90528 153922 90598 153978
rect 90654 153922 90722 153978
rect 90778 153922 90848 153978
rect 90528 153888 90848 153922
rect 121248 154350 121568 154384
rect 121248 154294 121318 154350
rect 121374 154294 121442 154350
rect 121498 154294 121568 154350
rect 121248 154226 121568 154294
rect 121248 154170 121318 154226
rect 121374 154170 121442 154226
rect 121498 154170 121568 154226
rect 121248 154102 121568 154170
rect 121248 154046 121318 154102
rect 121374 154046 121442 154102
rect 121498 154046 121568 154102
rect 121248 153978 121568 154046
rect 121248 153922 121318 153978
rect 121374 153922 121442 153978
rect 121498 153922 121568 153978
rect 121248 153888 121568 153922
rect 151968 154350 152288 154384
rect 151968 154294 152038 154350
rect 152094 154294 152162 154350
rect 152218 154294 152288 154350
rect 151968 154226 152288 154294
rect 151968 154170 152038 154226
rect 152094 154170 152162 154226
rect 152218 154170 152288 154226
rect 151968 154102 152288 154170
rect 151968 154046 152038 154102
rect 152094 154046 152162 154102
rect 152218 154046 152288 154102
rect 151968 153978 152288 154046
rect 151968 153922 152038 153978
rect 152094 153922 152162 153978
rect 152218 153922 152288 153978
rect 151968 153888 152288 153922
rect 182688 154350 183008 154384
rect 182688 154294 182758 154350
rect 182814 154294 182882 154350
rect 182938 154294 183008 154350
rect 182688 154226 183008 154294
rect 182688 154170 182758 154226
rect 182814 154170 182882 154226
rect 182938 154170 183008 154226
rect 182688 154102 183008 154170
rect 182688 154046 182758 154102
rect 182814 154046 182882 154102
rect 182938 154046 183008 154102
rect 182688 153978 183008 154046
rect 182688 153922 182758 153978
rect 182814 153922 182882 153978
rect 182938 153922 183008 153978
rect 182688 153888 183008 153922
rect 213408 154350 213728 154384
rect 213408 154294 213478 154350
rect 213534 154294 213602 154350
rect 213658 154294 213728 154350
rect 213408 154226 213728 154294
rect 213408 154170 213478 154226
rect 213534 154170 213602 154226
rect 213658 154170 213728 154226
rect 213408 154102 213728 154170
rect 213408 154046 213478 154102
rect 213534 154046 213602 154102
rect 213658 154046 213728 154102
rect 213408 153978 213728 154046
rect 213408 153922 213478 153978
rect 213534 153922 213602 153978
rect 213658 153922 213728 153978
rect 213408 153888 213728 153922
rect 244128 154350 244448 154384
rect 244128 154294 244198 154350
rect 244254 154294 244322 154350
rect 244378 154294 244448 154350
rect 244128 154226 244448 154294
rect 244128 154170 244198 154226
rect 244254 154170 244322 154226
rect 244378 154170 244448 154226
rect 244128 154102 244448 154170
rect 244128 154046 244198 154102
rect 244254 154046 244322 154102
rect 244378 154046 244448 154102
rect 244128 153978 244448 154046
rect 244128 153922 244198 153978
rect 244254 153922 244322 153978
rect 244378 153922 244448 153978
rect 244128 153888 244448 153922
rect 75168 148350 75488 148384
rect 75168 148294 75238 148350
rect 75294 148294 75362 148350
rect 75418 148294 75488 148350
rect 75168 148226 75488 148294
rect 75168 148170 75238 148226
rect 75294 148170 75362 148226
rect 75418 148170 75488 148226
rect 75168 148102 75488 148170
rect 75168 148046 75238 148102
rect 75294 148046 75362 148102
rect 75418 148046 75488 148102
rect 75168 147978 75488 148046
rect 75168 147922 75238 147978
rect 75294 147922 75362 147978
rect 75418 147922 75488 147978
rect 75168 147888 75488 147922
rect 105888 148350 106208 148384
rect 105888 148294 105958 148350
rect 106014 148294 106082 148350
rect 106138 148294 106208 148350
rect 105888 148226 106208 148294
rect 105888 148170 105958 148226
rect 106014 148170 106082 148226
rect 106138 148170 106208 148226
rect 105888 148102 106208 148170
rect 105888 148046 105958 148102
rect 106014 148046 106082 148102
rect 106138 148046 106208 148102
rect 105888 147978 106208 148046
rect 105888 147922 105958 147978
rect 106014 147922 106082 147978
rect 106138 147922 106208 147978
rect 105888 147888 106208 147922
rect 136608 148350 136928 148384
rect 136608 148294 136678 148350
rect 136734 148294 136802 148350
rect 136858 148294 136928 148350
rect 136608 148226 136928 148294
rect 136608 148170 136678 148226
rect 136734 148170 136802 148226
rect 136858 148170 136928 148226
rect 136608 148102 136928 148170
rect 136608 148046 136678 148102
rect 136734 148046 136802 148102
rect 136858 148046 136928 148102
rect 136608 147978 136928 148046
rect 136608 147922 136678 147978
rect 136734 147922 136802 147978
rect 136858 147922 136928 147978
rect 136608 147888 136928 147922
rect 167328 148350 167648 148384
rect 167328 148294 167398 148350
rect 167454 148294 167522 148350
rect 167578 148294 167648 148350
rect 167328 148226 167648 148294
rect 167328 148170 167398 148226
rect 167454 148170 167522 148226
rect 167578 148170 167648 148226
rect 167328 148102 167648 148170
rect 167328 148046 167398 148102
rect 167454 148046 167522 148102
rect 167578 148046 167648 148102
rect 167328 147978 167648 148046
rect 167328 147922 167398 147978
rect 167454 147922 167522 147978
rect 167578 147922 167648 147978
rect 167328 147888 167648 147922
rect 198048 148350 198368 148384
rect 198048 148294 198118 148350
rect 198174 148294 198242 148350
rect 198298 148294 198368 148350
rect 198048 148226 198368 148294
rect 198048 148170 198118 148226
rect 198174 148170 198242 148226
rect 198298 148170 198368 148226
rect 198048 148102 198368 148170
rect 198048 148046 198118 148102
rect 198174 148046 198242 148102
rect 198298 148046 198368 148102
rect 198048 147978 198368 148046
rect 198048 147922 198118 147978
rect 198174 147922 198242 147978
rect 198298 147922 198368 147978
rect 198048 147888 198368 147922
rect 228768 148350 229088 148384
rect 228768 148294 228838 148350
rect 228894 148294 228962 148350
rect 229018 148294 229088 148350
rect 228768 148226 229088 148294
rect 228768 148170 228838 148226
rect 228894 148170 228962 148226
rect 229018 148170 229088 148226
rect 228768 148102 229088 148170
rect 228768 148046 228838 148102
rect 228894 148046 228962 148102
rect 229018 148046 229088 148102
rect 228768 147978 229088 148046
rect 228768 147922 228838 147978
rect 228894 147922 228962 147978
rect 229018 147922 229088 147978
rect 228768 147888 229088 147922
rect 259488 148350 259808 148384
rect 259488 148294 259558 148350
rect 259614 148294 259682 148350
rect 259738 148294 259808 148350
rect 259488 148226 259808 148294
rect 259488 148170 259558 148226
rect 259614 148170 259682 148226
rect 259738 148170 259808 148226
rect 259488 148102 259808 148170
rect 259488 148046 259558 148102
rect 259614 148046 259682 148102
rect 259738 148046 259808 148102
rect 259488 147978 259808 148046
rect 259488 147922 259558 147978
rect 259614 147922 259682 147978
rect 259738 147922 259808 147978
rect 259488 147888 259808 147922
rect 59808 136350 60128 136384
rect 59808 136294 59878 136350
rect 59934 136294 60002 136350
rect 60058 136294 60128 136350
rect 59808 136226 60128 136294
rect 59808 136170 59878 136226
rect 59934 136170 60002 136226
rect 60058 136170 60128 136226
rect 59808 136102 60128 136170
rect 59808 136046 59878 136102
rect 59934 136046 60002 136102
rect 60058 136046 60128 136102
rect 59808 135978 60128 136046
rect 59808 135922 59878 135978
rect 59934 135922 60002 135978
rect 60058 135922 60128 135978
rect 59808 135888 60128 135922
rect 90528 136350 90848 136384
rect 90528 136294 90598 136350
rect 90654 136294 90722 136350
rect 90778 136294 90848 136350
rect 90528 136226 90848 136294
rect 90528 136170 90598 136226
rect 90654 136170 90722 136226
rect 90778 136170 90848 136226
rect 90528 136102 90848 136170
rect 90528 136046 90598 136102
rect 90654 136046 90722 136102
rect 90778 136046 90848 136102
rect 90528 135978 90848 136046
rect 90528 135922 90598 135978
rect 90654 135922 90722 135978
rect 90778 135922 90848 135978
rect 90528 135888 90848 135922
rect 121248 136350 121568 136384
rect 121248 136294 121318 136350
rect 121374 136294 121442 136350
rect 121498 136294 121568 136350
rect 121248 136226 121568 136294
rect 121248 136170 121318 136226
rect 121374 136170 121442 136226
rect 121498 136170 121568 136226
rect 121248 136102 121568 136170
rect 121248 136046 121318 136102
rect 121374 136046 121442 136102
rect 121498 136046 121568 136102
rect 121248 135978 121568 136046
rect 121248 135922 121318 135978
rect 121374 135922 121442 135978
rect 121498 135922 121568 135978
rect 121248 135888 121568 135922
rect 151968 136350 152288 136384
rect 151968 136294 152038 136350
rect 152094 136294 152162 136350
rect 152218 136294 152288 136350
rect 151968 136226 152288 136294
rect 151968 136170 152038 136226
rect 152094 136170 152162 136226
rect 152218 136170 152288 136226
rect 151968 136102 152288 136170
rect 151968 136046 152038 136102
rect 152094 136046 152162 136102
rect 152218 136046 152288 136102
rect 151968 135978 152288 136046
rect 151968 135922 152038 135978
rect 152094 135922 152162 135978
rect 152218 135922 152288 135978
rect 151968 135888 152288 135922
rect 182688 136350 183008 136384
rect 182688 136294 182758 136350
rect 182814 136294 182882 136350
rect 182938 136294 183008 136350
rect 182688 136226 183008 136294
rect 182688 136170 182758 136226
rect 182814 136170 182882 136226
rect 182938 136170 183008 136226
rect 182688 136102 183008 136170
rect 182688 136046 182758 136102
rect 182814 136046 182882 136102
rect 182938 136046 183008 136102
rect 182688 135978 183008 136046
rect 182688 135922 182758 135978
rect 182814 135922 182882 135978
rect 182938 135922 183008 135978
rect 182688 135888 183008 135922
rect 213408 136350 213728 136384
rect 213408 136294 213478 136350
rect 213534 136294 213602 136350
rect 213658 136294 213728 136350
rect 213408 136226 213728 136294
rect 213408 136170 213478 136226
rect 213534 136170 213602 136226
rect 213658 136170 213728 136226
rect 213408 136102 213728 136170
rect 213408 136046 213478 136102
rect 213534 136046 213602 136102
rect 213658 136046 213728 136102
rect 213408 135978 213728 136046
rect 213408 135922 213478 135978
rect 213534 135922 213602 135978
rect 213658 135922 213728 135978
rect 213408 135888 213728 135922
rect 244128 136350 244448 136384
rect 244128 136294 244198 136350
rect 244254 136294 244322 136350
rect 244378 136294 244448 136350
rect 244128 136226 244448 136294
rect 244128 136170 244198 136226
rect 244254 136170 244322 136226
rect 244378 136170 244448 136226
rect 244128 136102 244448 136170
rect 244128 136046 244198 136102
rect 244254 136046 244322 136102
rect 244378 136046 244448 136102
rect 244128 135978 244448 136046
rect 244128 135922 244198 135978
rect 244254 135922 244322 135978
rect 244378 135922 244448 135978
rect 244128 135888 244448 135922
rect 75168 130350 75488 130384
rect 75168 130294 75238 130350
rect 75294 130294 75362 130350
rect 75418 130294 75488 130350
rect 75168 130226 75488 130294
rect 75168 130170 75238 130226
rect 75294 130170 75362 130226
rect 75418 130170 75488 130226
rect 75168 130102 75488 130170
rect 75168 130046 75238 130102
rect 75294 130046 75362 130102
rect 75418 130046 75488 130102
rect 75168 129978 75488 130046
rect 75168 129922 75238 129978
rect 75294 129922 75362 129978
rect 75418 129922 75488 129978
rect 75168 129888 75488 129922
rect 105888 130350 106208 130384
rect 105888 130294 105958 130350
rect 106014 130294 106082 130350
rect 106138 130294 106208 130350
rect 105888 130226 106208 130294
rect 105888 130170 105958 130226
rect 106014 130170 106082 130226
rect 106138 130170 106208 130226
rect 105888 130102 106208 130170
rect 105888 130046 105958 130102
rect 106014 130046 106082 130102
rect 106138 130046 106208 130102
rect 105888 129978 106208 130046
rect 105888 129922 105958 129978
rect 106014 129922 106082 129978
rect 106138 129922 106208 129978
rect 105888 129888 106208 129922
rect 136608 130350 136928 130384
rect 136608 130294 136678 130350
rect 136734 130294 136802 130350
rect 136858 130294 136928 130350
rect 136608 130226 136928 130294
rect 136608 130170 136678 130226
rect 136734 130170 136802 130226
rect 136858 130170 136928 130226
rect 136608 130102 136928 130170
rect 136608 130046 136678 130102
rect 136734 130046 136802 130102
rect 136858 130046 136928 130102
rect 136608 129978 136928 130046
rect 136608 129922 136678 129978
rect 136734 129922 136802 129978
rect 136858 129922 136928 129978
rect 136608 129888 136928 129922
rect 167328 130350 167648 130384
rect 167328 130294 167398 130350
rect 167454 130294 167522 130350
rect 167578 130294 167648 130350
rect 167328 130226 167648 130294
rect 167328 130170 167398 130226
rect 167454 130170 167522 130226
rect 167578 130170 167648 130226
rect 167328 130102 167648 130170
rect 167328 130046 167398 130102
rect 167454 130046 167522 130102
rect 167578 130046 167648 130102
rect 167328 129978 167648 130046
rect 167328 129922 167398 129978
rect 167454 129922 167522 129978
rect 167578 129922 167648 129978
rect 167328 129888 167648 129922
rect 198048 130350 198368 130384
rect 198048 130294 198118 130350
rect 198174 130294 198242 130350
rect 198298 130294 198368 130350
rect 198048 130226 198368 130294
rect 198048 130170 198118 130226
rect 198174 130170 198242 130226
rect 198298 130170 198368 130226
rect 198048 130102 198368 130170
rect 198048 130046 198118 130102
rect 198174 130046 198242 130102
rect 198298 130046 198368 130102
rect 198048 129978 198368 130046
rect 198048 129922 198118 129978
rect 198174 129922 198242 129978
rect 198298 129922 198368 129978
rect 198048 129888 198368 129922
rect 228768 130350 229088 130384
rect 228768 130294 228838 130350
rect 228894 130294 228962 130350
rect 229018 130294 229088 130350
rect 228768 130226 229088 130294
rect 228768 130170 228838 130226
rect 228894 130170 228962 130226
rect 229018 130170 229088 130226
rect 228768 130102 229088 130170
rect 228768 130046 228838 130102
rect 228894 130046 228962 130102
rect 229018 130046 229088 130102
rect 228768 129978 229088 130046
rect 228768 129922 228838 129978
rect 228894 129922 228962 129978
rect 229018 129922 229088 129978
rect 228768 129888 229088 129922
rect 259488 130350 259808 130384
rect 259488 130294 259558 130350
rect 259614 130294 259682 130350
rect 259738 130294 259808 130350
rect 259488 130226 259808 130294
rect 259488 130170 259558 130226
rect 259614 130170 259682 130226
rect 259738 130170 259808 130226
rect 259488 130102 259808 130170
rect 259488 130046 259558 130102
rect 259614 130046 259682 130102
rect 259738 130046 259808 130102
rect 259488 129978 259808 130046
rect 259488 129922 259558 129978
rect 259614 129922 259682 129978
rect 259738 129922 259808 129978
rect 259488 129888 259808 129922
rect 59808 118350 60128 118384
rect 59808 118294 59878 118350
rect 59934 118294 60002 118350
rect 60058 118294 60128 118350
rect 59808 118226 60128 118294
rect 59808 118170 59878 118226
rect 59934 118170 60002 118226
rect 60058 118170 60128 118226
rect 59808 118102 60128 118170
rect 59808 118046 59878 118102
rect 59934 118046 60002 118102
rect 60058 118046 60128 118102
rect 59808 117978 60128 118046
rect 59808 117922 59878 117978
rect 59934 117922 60002 117978
rect 60058 117922 60128 117978
rect 59808 117888 60128 117922
rect 90528 118350 90848 118384
rect 90528 118294 90598 118350
rect 90654 118294 90722 118350
rect 90778 118294 90848 118350
rect 90528 118226 90848 118294
rect 90528 118170 90598 118226
rect 90654 118170 90722 118226
rect 90778 118170 90848 118226
rect 90528 118102 90848 118170
rect 90528 118046 90598 118102
rect 90654 118046 90722 118102
rect 90778 118046 90848 118102
rect 90528 117978 90848 118046
rect 90528 117922 90598 117978
rect 90654 117922 90722 117978
rect 90778 117922 90848 117978
rect 90528 117888 90848 117922
rect 121248 118350 121568 118384
rect 121248 118294 121318 118350
rect 121374 118294 121442 118350
rect 121498 118294 121568 118350
rect 121248 118226 121568 118294
rect 121248 118170 121318 118226
rect 121374 118170 121442 118226
rect 121498 118170 121568 118226
rect 121248 118102 121568 118170
rect 121248 118046 121318 118102
rect 121374 118046 121442 118102
rect 121498 118046 121568 118102
rect 121248 117978 121568 118046
rect 121248 117922 121318 117978
rect 121374 117922 121442 117978
rect 121498 117922 121568 117978
rect 121248 117888 121568 117922
rect 151968 118350 152288 118384
rect 151968 118294 152038 118350
rect 152094 118294 152162 118350
rect 152218 118294 152288 118350
rect 151968 118226 152288 118294
rect 151968 118170 152038 118226
rect 152094 118170 152162 118226
rect 152218 118170 152288 118226
rect 151968 118102 152288 118170
rect 151968 118046 152038 118102
rect 152094 118046 152162 118102
rect 152218 118046 152288 118102
rect 151968 117978 152288 118046
rect 151968 117922 152038 117978
rect 152094 117922 152162 117978
rect 152218 117922 152288 117978
rect 151968 117888 152288 117922
rect 182688 118350 183008 118384
rect 182688 118294 182758 118350
rect 182814 118294 182882 118350
rect 182938 118294 183008 118350
rect 182688 118226 183008 118294
rect 182688 118170 182758 118226
rect 182814 118170 182882 118226
rect 182938 118170 183008 118226
rect 182688 118102 183008 118170
rect 182688 118046 182758 118102
rect 182814 118046 182882 118102
rect 182938 118046 183008 118102
rect 182688 117978 183008 118046
rect 182688 117922 182758 117978
rect 182814 117922 182882 117978
rect 182938 117922 183008 117978
rect 182688 117888 183008 117922
rect 213408 118350 213728 118384
rect 213408 118294 213478 118350
rect 213534 118294 213602 118350
rect 213658 118294 213728 118350
rect 213408 118226 213728 118294
rect 213408 118170 213478 118226
rect 213534 118170 213602 118226
rect 213658 118170 213728 118226
rect 213408 118102 213728 118170
rect 213408 118046 213478 118102
rect 213534 118046 213602 118102
rect 213658 118046 213728 118102
rect 213408 117978 213728 118046
rect 213408 117922 213478 117978
rect 213534 117922 213602 117978
rect 213658 117922 213728 117978
rect 213408 117888 213728 117922
rect 244128 118350 244448 118384
rect 244128 118294 244198 118350
rect 244254 118294 244322 118350
rect 244378 118294 244448 118350
rect 244128 118226 244448 118294
rect 244128 118170 244198 118226
rect 244254 118170 244322 118226
rect 244378 118170 244448 118226
rect 244128 118102 244448 118170
rect 244128 118046 244198 118102
rect 244254 118046 244322 118102
rect 244378 118046 244448 118102
rect 244128 117978 244448 118046
rect 244128 117922 244198 117978
rect 244254 117922 244322 117978
rect 244378 117922 244448 117978
rect 244128 117888 244448 117922
rect 75168 112350 75488 112384
rect 75168 112294 75238 112350
rect 75294 112294 75362 112350
rect 75418 112294 75488 112350
rect 75168 112226 75488 112294
rect 75168 112170 75238 112226
rect 75294 112170 75362 112226
rect 75418 112170 75488 112226
rect 75168 112102 75488 112170
rect 75168 112046 75238 112102
rect 75294 112046 75362 112102
rect 75418 112046 75488 112102
rect 75168 111978 75488 112046
rect 75168 111922 75238 111978
rect 75294 111922 75362 111978
rect 75418 111922 75488 111978
rect 75168 111888 75488 111922
rect 105888 112350 106208 112384
rect 105888 112294 105958 112350
rect 106014 112294 106082 112350
rect 106138 112294 106208 112350
rect 105888 112226 106208 112294
rect 105888 112170 105958 112226
rect 106014 112170 106082 112226
rect 106138 112170 106208 112226
rect 105888 112102 106208 112170
rect 105888 112046 105958 112102
rect 106014 112046 106082 112102
rect 106138 112046 106208 112102
rect 105888 111978 106208 112046
rect 105888 111922 105958 111978
rect 106014 111922 106082 111978
rect 106138 111922 106208 111978
rect 105888 111888 106208 111922
rect 136608 112350 136928 112384
rect 136608 112294 136678 112350
rect 136734 112294 136802 112350
rect 136858 112294 136928 112350
rect 136608 112226 136928 112294
rect 136608 112170 136678 112226
rect 136734 112170 136802 112226
rect 136858 112170 136928 112226
rect 136608 112102 136928 112170
rect 136608 112046 136678 112102
rect 136734 112046 136802 112102
rect 136858 112046 136928 112102
rect 136608 111978 136928 112046
rect 136608 111922 136678 111978
rect 136734 111922 136802 111978
rect 136858 111922 136928 111978
rect 136608 111888 136928 111922
rect 167328 112350 167648 112384
rect 167328 112294 167398 112350
rect 167454 112294 167522 112350
rect 167578 112294 167648 112350
rect 167328 112226 167648 112294
rect 167328 112170 167398 112226
rect 167454 112170 167522 112226
rect 167578 112170 167648 112226
rect 167328 112102 167648 112170
rect 167328 112046 167398 112102
rect 167454 112046 167522 112102
rect 167578 112046 167648 112102
rect 167328 111978 167648 112046
rect 167328 111922 167398 111978
rect 167454 111922 167522 111978
rect 167578 111922 167648 111978
rect 167328 111888 167648 111922
rect 198048 112350 198368 112384
rect 198048 112294 198118 112350
rect 198174 112294 198242 112350
rect 198298 112294 198368 112350
rect 198048 112226 198368 112294
rect 198048 112170 198118 112226
rect 198174 112170 198242 112226
rect 198298 112170 198368 112226
rect 198048 112102 198368 112170
rect 198048 112046 198118 112102
rect 198174 112046 198242 112102
rect 198298 112046 198368 112102
rect 198048 111978 198368 112046
rect 198048 111922 198118 111978
rect 198174 111922 198242 111978
rect 198298 111922 198368 111978
rect 198048 111888 198368 111922
rect 228768 112350 229088 112384
rect 228768 112294 228838 112350
rect 228894 112294 228962 112350
rect 229018 112294 229088 112350
rect 228768 112226 229088 112294
rect 228768 112170 228838 112226
rect 228894 112170 228962 112226
rect 229018 112170 229088 112226
rect 228768 112102 229088 112170
rect 228768 112046 228838 112102
rect 228894 112046 228962 112102
rect 229018 112046 229088 112102
rect 228768 111978 229088 112046
rect 228768 111922 228838 111978
rect 228894 111922 228962 111978
rect 229018 111922 229088 111978
rect 228768 111888 229088 111922
rect 259488 112350 259808 112384
rect 259488 112294 259558 112350
rect 259614 112294 259682 112350
rect 259738 112294 259808 112350
rect 259488 112226 259808 112294
rect 259488 112170 259558 112226
rect 259614 112170 259682 112226
rect 259738 112170 259808 112226
rect 259488 112102 259808 112170
rect 259488 112046 259558 112102
rect 259614 112046 259682 112102
rect 259738 112046 259808 112102
rect 259488 111978 259808 112046
rect 259488 111922 259558 111978
rect 259614 111922 259682 111978
rect 259738 111922 259808 111978
rect 259488 111888 259808 111922
rect 59808 100350 60128 100384
rect 59808 100294 59878 100350
rect 59934 100294 60002 100350
rect 60058 100294 60128 100350
rect 59808 100226 60128 100294
rect 59808 100170 59878 100226
rect 59934 100170 60002 100226
rect 60058 100170 60128 100226
rect 59808 100102 60128 100170
rect 59808 100046 59878 100102
rect 59934 100046 60002 100102
rect 60058 100046 60128 100102
rect 59808 99978 60128 100046
rect 59808 99922 59878 99978
rect 59934 99922 60002 99978
rect 60058 99922 60128 99978
rect 59808 99888 60128 99922
rect 90528 100350 90848 100384
rect 90528 100294 90598 100350
rect 90654 100294 90722 100350
rect 90778 100294 90848 100350
rect 90528 100226 90848 100294
rect 90528 100170 90598 100226
rect 90654 100170 90722 100226
rect 90778 100170 90848 100226
rect 90528 100102 90848 100170
rect 90528 100046 90598 100102
rect 90654 100046 90722 100102
rect 90778 100046 90848 100102
rect 90528 99978 90848 100046
rect 90528 99922 90598 99978
rect 90654 99922 90722 99978
rect 90778 99922 90848 99978
rect 90528 99888 90848 99922
rect 121248 100350 121568 100384
rect 121248 100294 121318 100350
rect 121374 100294 121442 100350
rect 121498 100294 121568 100350
rect 121248 100226 121568 100294
rect 121248 100170 121318 100226
rect 121374 100170 121442 100226
rect 121498 100170 121568 100226
rect 121248 100102 121568 100170
rect 121248 100046 121318 100102
rect 121374 100046 121442 100102
rect 121498 100046 121568 100102
rect 121248 99978 121568 100046
rect 121248 99922 121318 99978
rect 121374 99922 121442 99978
rect 121498 99922 121568 99978
rect 121248 99888 121568 99922
rect 151968 100350 152288 100384
rect 151968 100294 152038 100350
rect 152094 100294 152162 100350
rect 152218 100294 152288 100350
rect 151968 100226 152288 100294
rect 151968 100170 152038 100226
rect 152094 100170 152162 100226
rect 152218 100170 152288 100226
rect 151968 100102 152288 100170
rect 151968 100046 152038 100102
rect 152094 100046 152162 100102
rect 152218 100046 152288 100102
rect 151968 99978 152288 100046
rect 151968 99922 152038 99978
rect 152094 99922 152162 99978
rect 152218 99922 152288 99978
rect 151968 99888 152288 99922
rect 182688 100350 183008 100384
rect 182688 100294 182758 100350
rect 182814 100294 182882 100350
rect 182938 100294 183008 100350
rect 182688 100226 183008 100294
rect 182688 100170 182758 100226
rect 182814 100170 182882 100226
rect 182938 100170 183008 100226
rect 182688 100102 183008 100170
rect 182688 100046 182758 100102
rect 182814 100046 182882 100102
rect 182938 100046 183008 100102
rect 182688 99978 183008 100046
rect 182688 99922 182758 99978
rect 182814 99922 182882 99978
rect 182938 99922 183008 99978
rect 182688 99888 183008 99922
rect 213408 100350 213728 100384
rect 213408 100294 213478 100350
rect 213534 100294 213602 100350
rect 213658 100294 213728 100350
rect 213408 100226 213728 100294
rect 213408 100170 213478 100226
rect 213534 100170 213602 100226
rect 213658 100170 213728 100226
rect 213408 100102 213728 100170
rect 213408 100046 213478 100102
rect 213534 100046 213602 100102
rect 213658 100046 213728 100102
rect 213408 99978 213728 100046
rect 213408 99922 213478 99978
rect 213534 99922 213602 99978
rect 213658 99922 213728 99978
rect 213408 99888 213728 99922
rect 244128 100350 244448 100384
rect 244128 100294 244198 100350
rect 244254 100294 244322 100350
rect 244378 100294 244448 100350
rect 244128 100226 244448 100294
rect 244128 100170 244198 100226
rect 244254 100170 244322 100226
rect 244378 100170 244448 100226
rect 244128 100102 244448 100170
rect 244128 100046 244198 100102
rect 244254 100046 244322 100102
rect 244378 100046 244448 100102
rect 244128 99978 244448 100046
rect 244128 99922 244198 99978
rect 244254 99922 244322 99978
rect 244378 99922 244448 99978
rect 244128 99888 244448 99922
rect 75168 94350 75488 94384
rect 75168 94294 75238 94350
rect 75294 94294 75362 94350
rect 75418 94294 75488 94350
rect 75168 94226 75488 94294
rect 75168 94170 75238 94226
rect 75294 94170 75362 94226
rect 75418 94170 75488 94226
rect 75168 94102 75488 94170
rect 75168 94046 75238 94102
rect 75294 94046 75362 94102
rect 75418 94046 75488 94102
rect 75168 93978 75488 94046
rect 75168 93922 75238 93978
rect 75294 93922 75362 93978
rect 75418 93922 75488 93978
rect 75168 93888 75488 93922
rect 105888 94350 106208 94384
rect 105888 94294 105958 94350
rect 106014 94294 106082 94350
rect 106138 94294 106208 94350
rect 105888 94226 106208 94294
rect 105888 94170 105958 94226
rect 106014 94170 106082 94226
rect 106138 94170 106208 94226
rect 105888 94102 106208 94170
rect 105888 94046 105958 94102
rect 106014 94046 106082 94102
rect 106138 94046 106208 94102
rect 105888 93978 106208 94046
rect 105888 93922 105958 93978
rect 106014 93922 106082 93978
rect 106138 93922 106208 93978
rect 105888 93888 106208 93922
rect 136608 94350 136928 94384
rect 136608 94294 136678 94350
rect 136734 94294 136802 94350
rect 136858 94294 136928 94350
rect 136608 94226 136928 94294
rect 136608 94170 136678 94226
rect 136734 94170 136802 94226
rect 136858 94170 136928 94226
rect 136608 94102 136928 94170
rect 136608 94046 136678 94102
rect 136734 94046 136802 94102
rect 136858 94046 136928 94102
rect 136608 93978 136928 94046
rect 136608 93922 136678 93978
rect 136734 93922 136802 93978
rect 136858 93922 136928 93978
rect 136608 93888 136928 93922
rect 167328 94350 167648 94384
rect 167328 94294 167398 94350
rect 167454 94294 167522 94350
rect 167578 94294 167648 94350
rect 167328 94226 167648 94294
rect 167328 94170 167398 94226
rect 167454 94170 167522 94226
rect 167578 94170 167648 94226
rect 167328 94102 167648 94170
rect 167328 94046 167398 94102
rect 167454 94046 167522 94102
rect 167578 94046 167648 94102
rect 167328 93978 167648 94046
rect 167328 93922 167398 93978
rect 167454 93922 167522 93978
rect 167578 93922 167648 93978
rect 167328 93888 167648 93922
rect 198048 94350 198368 94384
rect 198048 94294 198118 94350
rect 198174 94294 198242 94350
rect 198298 94294 198368 94350
rect 198048 94226 198368 94294
rect 198048 94170 198118 94226
rect 198174 94170 198242 94226
rect 198298 94170 198368 94226
rect 198048 94102 198368 94170
rect 198048 94046 198118 94102
rect 198174 94046 198242 94102
rect 198298 94046 198368 94102
rect 198048 93978 198368 94046
rect 198048 93922 198118 93978
rect 198174 93922 198242 93978
rect 198298 93922 198368 93978
rect 198048 93888 198368 93922
rect 228768 94350 229088 94384
rect 228768 94294 228838 94350
rect 228894 94294 228962 94350
rect 229018 94294 229088 94350
rect 228768 94226 229088 94294
rect 228768 94170 228838 94226
rect 228894 94170 228962 94226
rect 229018 94170 229088 94226
rect 228768 94102 229088 94170
rect 228768 94046 228838 94102
rect 228894 94046 228962 94102
rect 229018 94046 229088 94102
rect 228768 93978 229088 94046
rect 228768 93922 228838 93978
rect 228894 93922 228962 93978
rect 229018 93922 229088 93978
rect 228768 93888 229088 93922
rect 259488 94350 259808 94384
rect 259488 94294 259558 94350
rect 259614 94294 259682 94350
rect 259738 94294 259808 94350
rect 259488 94226 259808 94294
rect 259488 94170 259558 94226
rect 259614 94170 259682 94226
rect 259738 94170 259808 94226
rect 259488 94102 259808 94170
rect 259488 94046 259558 94102
rect 259614 94046 259682 94102
rect 259738 94046 259808 94102
rect 259488 93978 259808 94046
rect 259488 93922 259558 93978
rect 259614 93922 259682 93978
rect 259738 93922 259808 93978
rect 259488 93888 259808 93922
rect 59808 82350 60128 82384
rect 59808 82294 59878 82350
rect 59934 82294 60002 82350
rect 60058 82294 60128 82350
rect 59808 82226 60128 82294
rect 59808 82170 59878 82226
rect 59934 82170 60002 82226
rect 60058 82170 60128 82226
rect 59808 82102 60128 82170
rect 59808 82046 59878 82102
rect 59934 82046 60002 82102
rect 60058 82046 60128 82102
rect 59808 81978 60128 82046
rect 59808 81922 59878 81978
rect 59934 81922 60002 81978
rect 60058 81922 60128 81978
rect 59808 81888 60128 81922
rect 90528 82350 90848 82384
rect 90528 82294 90598 82350
rect 90654 82294 90722 82350
rect 90778 82294 90848 82350
rect 90528 82226 90848 82294
rect 90528 82170 90598 82226
rect 90654 82170 90722 82226
rect 90778 82170 90848 82226
rect 90528 82102 90848 82170
rect 90528 82046 90598 82102
rect 90654 82046 90722 82102
rect 90778 82046 90848 82102
rect 90528 81978 90848 82046
rect 90528 81922 90598 81978
rect 90654 81922 90722 81978
rect 90778 81922 90848 81978
rect 90528 81888 90848 81922
rect 121248 82350 121568 82384
rect 121248 82294 121318 82350
rect 121374 82294 121442 82350
rect 121498 82294 121568 82350
rect 121248 82226 121568 82294
rect 121248 82170 121318 82226
rect 121374 82170 121442 82226
rect 121498 82170 121568 82226
rect 121248 82102 121568 82170
rect 121248 82046 121318 82102
rect 121374 82046 121442 82102
rect 121498 82046 121568 82102
rect 121248 81978 121568 82046
rect 121248 81922 121318 81978
rect 121374 81922 121442 81978
rect 121498 81922 121568 81978
rect 121248 81888 121568 81922
rect 151968 82350 152288 82384
rect 151968 82294 152038 82350
rect 152094 82294 152162 82350
rect 152218 82294 152288 82350
rect 151968 82226 152288 82294
rect 151968 82170 152038 82226
rect 152094 82170 152162 82226
rect 152218 82170 152288 82226
rect 151968 82102 152288 82170
rect 151968 82046 152038 82102
rect 152094 82046 152162 82102
rect 152218 82046 152288 82102
rect 151968 81978 152288 82046
rect 151968 81922 152038 81978
rect 152094 81922 152162 81978
rect 152218 81922 152288 81978
rect 151968 81888 152288 81922
rect 182688 82350 183008 82384
rect 182688 82294 182758 82350
rect 182814 82294 182882 82350
rect 182938 82294 183008 82350
rect 182688 82226 183008 82294
rect 182688 82170 182758 82226
rect 182814 82170 182882 82226
rect 182938 82170 183008 82226
rect 182688 82102 183008 82170
rect 182688 82046 182758 82102
rect 182814 82046 182882 82102
rect 182938 82046 183008 82102
rect 182688 81978 183008 82046
rect 182688 81922 182758 81978
rect 182814 81922 182882 81978
rect 182938 81922 183008 81978
rect 182688 81888 183008 81922
rect 213408 82350 213728 82384
rect 213408 82294 213478 82350
rect 213534 82294 213602 82350
rect 213658 82294 213728 82350
rect 213408 82226 213728 82294
rect 213408 82170 213478 82226
rect 213534 82170 213602 82226
rect 213658 82170 213728 82226
rect 213408 82102 213728 82170
rect 213408 82046 213478 82102
rect 213534 82046 213602 82102
rect 213658 82046 213728 82102
rect 213408 81978 213728 82046
rect 213408 81922 213478 81978
rect 213534 81922 213602 81978
rect 213658 81922 213728 81978
rect 213408 81888 213728 81922
rect 244128 82350 244448 82384
rect 244128 82294 244198 82350
rect 244254 82294 244322 82350
rect 244378 82294 244448 82350
rect 244128 82226 244448 82294
rect 244128 82170 244198 82226
rect 244254 82170 244322 82226
rect 244378 82170 244448 82226
rect 244128 82102 244448 82170
rect 244128 82046 244198 82102
rect 244254 82046 244322 82102
rect 244378 82046 244448 82102
rect 244128 81978 244448 82046
rect 244128 81922 244198 81978
rect 244254 81922 244322 81978
rect 244378 81922 244448 81978
rect 244128 81888 244448 81922
rect 75168 76350 75488 76384
rect 75168 76294 75238 76350
rect 75294 76294 75362 76350
rect 75418 76294 75488 76350
rect 75168 76226 75488 76294
rect 75168 76170 75238 76226
rect 75294 76170 75362 76226
rect 75418 76170 75488 76226
rect 75168 76102 75488 76170
rect 75168 76046 75238 76102
rect 75294 76046 75362 76102
rect 75418 76046 75488 76102
rect 75168 75978 75488 76046
rect 75168 75922 75238 75978
rect 75294 75922 75362 75978
rect 75418 75922 75488 75978
rect 75168 75888 75488 75922
rect 105888 76350 106208 76384
rect 105888 76294 105958 76350
rect 106014 76294 106082 76350
rect 106138 76294 106208 76350
rect 105888 76226 106208 76294
rect 105888 76170 105958 76226
rect 106014 76170 106082 76226
rect 106138 76170 106208 76226
rect 105888 76102 106208 76170
rect 105888 76046 105958 76102
rect 106014 76046 106082 76102
rect 106138 76046 106208 76102
rect 105888 75978 106208 76046
rect 105888 75922 105958 75978
rect 106014 75922 106082 75978
rect 106138 75922 106208 75978
rect 105888 75888 106208 75922
rect 136608 76350 136928 76384
rect 136608 76294 136678 76350
rect 136734 76294 136802 76350
rect 136858 76294 136928 76350
rect 136608 76226 136928 76294
rect 136608 76170 136678 76226
rect 136734 76170 136802 76226
rect 136858 76170 136928 76226
rect 136608 76102 136928 76170
rect 136608 76046 136678 76102
rect 136734 76046 136802 76102
rect 136858 76046 136928 76102
rect 136608 75978 136928 76046
rect 136608 75922 136678 75978
rect 136734 75922 136802 75978
rect 136858 75922 136928 75978
rect 136608 75888 136928 75922
rect 167328 76350 167648 76384
rect 167328 76294 167398 76350
rect 167454 76294 167522 76350
rect 167578 76294 167648 76350
rect 167328 76226 167648 76294
rect 167328 76170 167398 76226
rect 167454 76170 167522 76226
rect 167578 76170 167648 76226
rect 167328 76102 167648 76170
rect 167328 76046 167398 76102
rect 167454 76046 167522 76102
rect 167578 76046 167648 76102
rect 167328 75978 167648 76046
rect 167328 75922 167398 75978
rect 167454 75922 167522 75978
rect 167578 75922 167648 75978
rect 167328 75888 167648 75922
rect 198048 76350 198368 76384
rect 198048 76294 198118 76350
rect 198174 76294 198242 76350
rect 198298 76294 198368 76350
rect 198048 76226 198368 76294
rect 198048 76170 198118 76226
rect 198174 76170 198242 76226
rect 198298 76170 198368 76226
rect 198048 76102 198368 76170
rect 198048 76046 198118 76102
rect 198174 76046 198242 76102
rect 198298 76046 198368 76102
rect 198048 75978 198368 76046
rect 198048 75922 198118 75978
rect 198174 75922 198242 75978
rect 198298 75922 198368 75978
rect 198048 75888 198368 75922
rect 228768 76350 229088 76384
rect 228768 76294 228838 76350
rect 228894 76294 228962 76350
rect 229018 76294 229088 76350
rect 228768 76226 229088 76294
rect 228768 76170 228838 76226
rect 228894 76170 228962 76226
rect 229018 76170 229088 76226
rect 228768 76102 229088 76170
rect 228768 76046 228838 76102
rect 228894 76046 228962 76102
rect 229018 76046 229088 76102
rect 228768 75978 229088 76046
rect 228768 75922 228838 75978
rect 228894 75922 228962 75978
rect 229018 75922 229088 75978
rect 228768 75888 229088 75922
rect 259488 76350 259808 76384
rect 259488 76294 259558 76350
rect 259614 76294 259682 76350
rect 259738 76294 259808 76350
rect 259488 76226 259808 76294
rect 259488 76170 259558 76226
rect 259614 76170 259682 76226
rect 259738 76170 259808 76226
rect 259488 76102 259808 76170
rect 259488 76046 259558 76102
rect 259614 76046 259682 76102
rect 259738 76046 259808 76102
rect 259488 75978 259808 76046
rect 259488 75922 259558 75978
rect 259614 75922 259682 75978
rect 259738 75922 259808 75978
rect 259488 75888 259808 75922
rect 59808 64350 60128 64384
rect 59808 64294 59878 64350
rect 59934 64294 60002 64350
rect 60058 64294 60128 64350
rect 59808 64226 60128 64294
rect 59808 64170 59878 64226
rect 59934 64170 60002 64226
rect 60058 64170 60128 64226
rect 59808 64102 60128 64170
rect 59808 64046 59878 64102
rect 59934 64046 60002 64102
rect 60058 64046 60128 64102
rect 59808 63978 60128 64046
rect 59808 63922 59878 63978
rect 59934 63922 60002 63978
rect 60058 63922 60128 63978
rect 59808 63888 60128 63922
rect 90528 64350 90848 64384
rect 90528 64294 90598 64350
rect 90654 64294 90722 64350
rect 90778 64294 90848 64350
rect 90528 64226 90848 64294
rect 90528 64170 90598 64226
rect 90654 64170 90722 64226
rect 90778 64170 90848 64226
rect 90528 64102 90848 64170
rect 90528 64046 90598 64102
rect 90654 64046 90722 64102
rect 90778 64046 90848 64102
rect 90528 63978 90848 64046
rect 90528 63922 90598 63978
rect 90654 63922 90722 63978
rect 90778 63922 90848 63978
rect 90528 63888 90848 63922
rect 121248 64350 121568 64384
rect 121248 64294 121318 64350
rect 121374 64294 121442 64350
rect 121498 64294 121568 64350
rect 121248 64226 121568 64294
rect 121248 64170 121318 64226
rect 121374 64170 121442 64226
rect 121498 64170 121568 64226
rect 121248 64102 121568 64170
rect 121248 64046 121318 64102
rect 121374 64046 121442 64102
rect 121498 64046 121568 64102
rect 121248 63978 121568 64046
rect 121248 63922 121318 63978
rect 121374 63922 121442 63978
rect 121498 63922 121568 63978
rect 121248 63888 121568 63922
rect 151968 64350 152288 64384
rect 151968 64294 152038 64350
rect 152094 64294 152162 64350
rect 152218 64294 152288 64350
rect 151968 64226 152288 64294
rect 151968 64170 152038 64226
rect 152094 64170 152162 64226
rect 152218 64170 152288 64226
rect 151968 64102 152288 64170
rect 151968 64046 152038 64102
rect 152094 64046 152162 64102
rect 152218 64046 152288 64102
rect 151968 63978 152288 64046
rect 151968 63922 152038 63978
rect 152094 63922 152162 63978
rect 152218 63922 152288 63978
rect 151968 63888 152288 63922
rect 182688 64350 183008 64384
rect 182688 64294 182758 64350
rect 182814 64294 182882 64350
rect 182938 64294 183008 64350
rect 182688 64226 183008 64294
rect 182688 64170 182758 64226
rect 182814 64170 182882 64226
rect 182938 64170 183008 64226
rect 182688 64102 183008 64170
rect 182688 64046 182758 64102
rect 182814 64046 182882 64102
rect 182938 64046 183008 64102
rect 182688 63978 183008 64046
rect 182688 63922 182758 63978
rect 182814 63922 182882 63978
rect 182938 63922 183008 63978
rect 182688 63888 183008 63922
rect 213408 64350 213728 64384
rect 213408 64294 213478 64350
rect 213534 64294 213602 64350
rect 213658 64294 213728 64350
rect 213408 64226 213728 64294
rect 213408 64170 213478 64226
rect 213534 64170 213602 64226
rect 213658 64170 213728 64226
rect 213408 64102 213728 64170
rect 213408 64046 213478 64102
rect 213534 64046 213602 64102
rect 213658 64046 213728 64102
rect 213408 63978 213728 64046
rect 213408 63922 213478 63978
rect 213534 63922 213602 63978
rect 213658 63922 213728 63978
rect 213408 63888 213728 63922
rect 244128 64350 244448 64384
rect 244128 64294 244198 64350
rect 244254 64294 244322 64350
rect 244378 64294 244448 64350
rect 244128 64226 244448 64294
rect 244128 64170 244198 64226
rect 244254 64170 244322 64226
rect 244378 64170 244448 64226
rect 244128 64102 244448 64170
rect 244128 64046 244198 64102
rect 244254 64046 244322 64102
rect 244378 64046 244448 64102
rect 244128 63978 244448 64046
rect 244128 63922 244198 63978
rect 244254 63922 244322 63978
rect 244378 63922 244448 63978
rect 244128 63888 244448 63922
rect 75168 58350 75488 58384
rect 75168 58294 75238 58350
rect 75294 58294 75362 58350
rect 75418 58294 75488 58350
rect 75168 58226 75488 58294
rect 75168 58170 75238 58226
rect 75294 58170 75362 58226
rect 75418 58170 75488 58226
rect 75168 58102 75488 58170
rect 75168 58046 75238 58102
rect 75294 58046 75362 58102
rect 75418 58046 75488 58102
rect 75168 57978 75488 58046
rect 75168 57922 75238 57978
rect 75294 57922 75362 57978
rect 75418 57922 75488 57978
rect 75168 57888 75488 57922
rect 105888 58350 106208 58384
rect 105888 58294 105958 58350
rect 106014 58294 106082 58350
rect 106138 58294 106208 58350
rect 105888 58226 106208 58294
rect 105888 58170 105958 58226
rect 106014 58170 106082 58226
rect 106138 58170 106208 58226
rect 105888 58102 106208 58170
rect 105888 58046 105958 58102
rect 106014 58046 106082 58102
rect 106138 58046 106208 58102
rect 105888 57978 106208 58046
rect 105888 57922 105958 57978
rect 106014 57922 106082 57978
rect 106138 57922 106208 57978
rect 105888 57888 106208 57922
rect 136608 58350 136928 58384
rect 136608 58294 136678 58350
rect 136734 58294 136802 58350
rect 136858 58294 136928 58350
rect 136608 58226 136928 58294
rect 136608 58170 136678 58226
rect 136734 58170 136802 58226
rect 136858 58170 136928 58226
rect 136608 58102 136928 58170
rect 136608 58046 136678 58102
rect 136734 58046 136802 58102
rect 136858 58046 136928 58102
rect 136608 57978 136928 58046
rect 136608 57922 136678 57978
rect 136734 57922 136802 57978
rect 136858 57922 136928 57978
rect 136608 57888 136928 57922
rect 167328 58350 167648 58384
rect 167328 58294 167398 58350
rect 167454 58294 167522 58350
rect 167578 58294 167648 58350
rect 167328 58226 167648 58294
rect 167328 58170 167398 58226
rect 167454 58170 167522 58226
rect 167578 58170 167648 58226
rect 167328 58102 167648 58170
rect 167328 58046 167398 58102
rect 167454 58046 167522 58102
rect 167578 58046 167648 58102
rect 167328 57978 167648 58046
rect 167328 57922 167398 57978
rect 167454 57922 167522 57978
rect 167578 57922 167648 57978
rect 167328 57888 167648 57922
rect 198048 58350 198368 58384
rect 198048 58294 198118 58350
rect 198174 58294 198242 58350
rect 198298 58294 198368 58350
rect 198048 58226 198368 58294
rect 198048 58170 198118 58226
rect 198174 58170 198242 58226
rect 198298 58170 198368 58226
rect 198048 58102 198368 58170
rect 198048 58046 198118 58102
rect 198174 58046 198242 58102
rect 198298 58046 198368 58102
rect 198048 57978 198368 58046
rect 198048 57922 198118 57978
rect 198174 57922 198242 57978
rect 198298 57922 198368 57978
rect 198048 57888 198368 57922
rect 228768 58350 229088 58384
rect 228768 58294 228838 58350
rect 228894 58294 228962 58350
rect 229018 58294 229088 58350
rect 228768 58226 229088 58294
rect 228768 58170 228838 58226
rect 228894 58170 228962 58226
rect 229018 58170 229088 58226
rect 228768 58102 229088 58170
rect 228768 58046 228838 58102
rect 228894 58046 228962 58102
rect 229018 58046 229088 58102
rect 228768 57978 229088 58046
rect 228768 57922 228838 57978
rect 228894 57922 228962 57978
rect 229018 57922 229088 57978
rect 228768 57888 229088 57922
rect 259488 58350 259808 58384
rect 259488 58294 259558 58350
rect 259614 58294 259682 58350
rect 259738 58294 259808 58350
rect 259488 58226 259808 58294
rect 259488 58170 259558 58226
rect 259614 58170 259682 58226
rect 259738 58170 259808 58226
rect 259488 58102 259808 58170
rect 259488 58046 259558 58102
rect 259614 58046 259682 58102
rect 259738 58046 259808 58102
rect 259488 57978 259808 58046
rect 259488 57922 259558 57978
rect 259614 57922 259682 57978
rect 259738 57922 259808 57978
rect 259488 57888 259808 57922
rect 66858 40350 67478 48802
rect 66858 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 67478 40350
rect 66858 40226 67478 40294
rect 66858 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 67478 40226
rect 66858 40102 67478 40170
rect 66858 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 67478 40102
rect 66858 39978 67478 40046
rect 66858 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 67478 39978
rect 66858 22350 67478 39922
rect 66858 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 67478 22350
rect 66858 22226 67478 22294
rect 66858 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 67478 22226
rect 66858 22102 67478 22170
rect 66858 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 67478 22102
rect 66858 21978 67478 22046
rect 66858 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 67478 21978
rect 60844 4978 60900 4988
rect 51996 4274 52052 4284
rect 55132 4798 55188 4808
rect 48636 4162 48692 4172
rect 55132 3444 55188 4742
rect 55132 3378 55188 3388
rect 60844 3444 60900 4922
rect 60844 3378 60900 3388
rect 66858 4350 67478 21922
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 39858 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 40478 -1120
rect 39858 -1244 40478 -1176
rect 39858 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 40478 -1244
rect 39858 -1368 40478 -1300
rect 39858 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 40478 -1368
rect 39858 -1492 40478 -1424
rect 39858 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 40478 -1492
rect 39858 -1644 40478 -1548
rect 66858 -160 67478 3922
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 70578 46350 71198 48802
rect 70578 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 71198 46350
rect 70578 46226 71198 46294
rect 70578 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 71198 46226
rect 70578 46102 71198 46170
rect 70578 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 71198 46102
rect 70578 45978 71198 46046
rect 70578 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 71198 45978
rect 70578 28350 71198 45922
rect 70578 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 71198 28350
rect 70578 28226 71198 28294
rect 70578 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 71198 28226
rect 70578 28102 71198 28170
rect 70578 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 71198 28102
rect 70578 27978 71198 28046
rect 70578 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 71198 27978
rect 70578 10350 71198 27922
rect 70578 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 71198 10350
rect 70578 10226 71198 10294
rect 70578 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 71198 10226
rect 70578 10102 71198 10170
rect 70578 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 71198 10102
rect 70578 9978 71198 10046
rect 70578 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 71198 9978
rect 70578 -1120 71198 9922
rect 97578 40350 98198 48802
rect 97578 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 98198 40350
rect 97578 40226 98198 40294
rect 97578 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 98198 40226
rect 97578 40102 98198 40170
rect 97578 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 98198 40102
rect 97578 39978 98198 40046
rect 97578 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 98198 39978
rect 97578 22350 98198 39922
rect 97578 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 98198 22350
rect 97578 22226 98198 22294
rect 97578 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 98198 22226
rect 97578 22102 98198 22170
rect 97578 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 98198 22102
rect 97578 21978 98198 22046
rect 97578 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 98198 21978
rect 91532 4978 91588 4988
rect 91532 3444 91588 4922
rect 91532 3378 91588 3388
rect 97578 4350 98198 21922
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 97578 4102 98198 4170
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 70578 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 71198 -1120
rect 70578 -1244 71198 -1176
rect 70578 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 71198 -1244
rect 70578 -1368 71198 -1300
rect 70578 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 71198 -1368
rect 70578 -1492 71198 -1424
rect 70578 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 71198 -1492
rect 70578 -1644 71198 -1548
rect 97578 -160 98198 3922
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 101298 46350 101918 48802
rect 101298 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 101918 46350
rect 101298 46226 101918 46294
rect 101298 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 101918 46226
rect 101298 46102 101918 46170
rect 101298 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 101918 46102
rect 101298 45978 101918 46046
rect 101298 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 101918 45978
rect 101298 28350 101918 45922
rect 101298 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 101918 28350
rect 101298 28226 101918 28294
rect 101298 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 101918 28226
rect 101298 28102 101918 28170
rect 101298 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 101918 28102
rect 101298 27978 101918 28046
rect 101298 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 101918 27978
rect 101298 10350 101918 27922
rect 101298 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 101918 10350
rect 101298 10226 101918 10294
rect 101298 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 101918 10226
rect 101298 10102 101918 10170
rect 101298 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 101918 10102
rect 101298 9978 101918 10046
rect 101298 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 101918 9978
rect 101298 -1120 101918 9922
rect 101298 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 101918 -1120
rect 101298 -1244 101918 -1176
rect 101298 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 101918 -1244
rect 101298 -1368 101918 -1300
rect 101298 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 101918 -1368
rect 101298 -1492 101918 -1424
rect 101298 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 101918 -1492
rect 101298 -1644 101918 -1548
rect 128298 40350 128918 48802
rect 128298 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 128918 40350
rect 128298 40226 128918 40294
rect 128298 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 128918 40226
rect 128298 40102 128918 40170
rect 128298 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 128918 40102
rect 128298 39978 128918 40046
rect 128298 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 128918 39978
rect 128298 22350 128918 39922
rect 128298 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 128918 22350
rect 128298 22226 128918 22294
rect 128298 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 128918 22226
rect 128298 22102 128918 22170
rect 128298 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 128918 22102
rect 128298 21978 128918 22046
rect 128298 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 128918 21978
rect 128298 4350 128918 21922
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 128298 -160 128918 3922
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 132018 46350 132638 48802
rect 132018 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 132638 46350
rect 132018 46226 132638 46294
rect 132018 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 132638 46226
rect 132018 46102 132638 46170
rect 132018 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 132638 46102
rect 132018 45978 132638 46046
rect 132018 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 132638 45978
rect 132018 28350 132638 45922
rect 132018 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 132638 28350
rect 132018 28226 132638 28294
rect 132018 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 132638 28226
rect 132018 28102 132638 28170
rect 132018 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 132638 28102
rect 132018 27978 132638 28046
rect 132018 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 132638 27978
rect 132018 10350 132638 27922
rect 132018 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 132638 10350
rect 132018 10226 132638 10294
rect 132018 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 132638 10226
rect 132018 10102 132638 10170
rect 132018 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 132638 10102
rect 132018 9978 132638 10046
rect 132018 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 132638 9978
rect 132018 -1120 132638 9922
rect 159018 40350 159638 48802
rect 159018 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 159638 40350
rect 159018 40226 159638 40294
rect 159018 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 159638 40226
rect 159018 40102 159638 40170
rect 159018 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 159638 40102
rect 159018 39978 159638 40046
rect 159018 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 159638 39978
rect 159018 22350 159638 39922
rect 159018 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 159638 22350
rect 159018 22226 159638 22294
rect 159018 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 159638 22226
rect 159018 22102 159638 22170
rect 159018 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 159638 22102
rect 159018 21978 159638 22046
rect 159018 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 159638 21978
rect 142940 4798 142996 4808
rect 142940 3444 142996 4742
rect 142940 3378 142996 3388
rect 159018 4350 159638 21922
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 159018 4102 159638 4170
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 132018 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 132638 -1120
rect 132018 -1244 132638 -1176
rect 132018 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 132638 -1244
rect 132018 -1368 132638 -1300
rect 132018 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 132638 -1368
rect 132018 -1492 132638 -1424
rect 132018 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 132638 -1492
rect 132018 -1644 132638 -1548
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 162738 46350 163358 48802
rect 162738 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163358 46350
rect 162738 46226 163358 46294
rect 162738 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163358 46226
rect 162738 46102 163358 46170
rect 162738 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163358 46102
rect 162738 45978 163358 46046
rect 162738 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163358 45978
rect 162738 28350 163358 45922
rect 162738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 163358 28350
rect 162738 28226 163358 28294
rect 162738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 163358 28226
rect 162738 28102 163358 28170
rect 162738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 163358 28102
rect 162738 27978 163358 28046
rect 162738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 163358 27978
rect 162738 10350 163358 27922
rect 162738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 163358 10350
rect 162738 10226 163358 10294
rect 162738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 163358 10226
rect 162738 10102 163358 10170
rect 162738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 163358 10102
rect 162738 9978 163358 10046
rect 162738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 163358 9978
rect 162738 -1120 163358 9922
rect 172956 47818 173012 47828
rect 172956 4116 173012 47762
rect 172956 4050 173012 4060
rect 189738 40350 190358 48802
rect 189738 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 190358 40350
rect 189738 40226 190358 40294
rect 189738 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 190358 40226
rect 189738 40102 190358 40170
rect 189738 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 190358 40102
rect 189738 39978 190358 40046
rect 189738 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 190358 39978
rect 189738 22350 190358 39922
rect 189738 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 190358 22350
rect 189738 22226 190358 22294
rect 189738 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 190358 22226
rect 189738 22102 190358 22170
rect 189738 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 190358 22102
rect 189738 21978 190358 22046
rect 189738 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 190358 21978
rect 189738 4350 190358 21922
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 189738 4102 190358 4170
rect 162738 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 163358 -1120
rect 162738 -1244 163358 -1176
rect 162738 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 163358 -1244
rect 162738 -1368 163358 -1300
rect 162738 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 163358 -1368
rect 162738 -1492 163358 -1424
rect 162738 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 163358 -1492
rect 162738 -1644 163358 -1548
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 189738 -160 190358 3922
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 193458 46350 194078 48802
rect 193458 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 194078 46350
rect 193458 46226 194078 46294
rect 193458 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 194078 46226
rect 193458 46102 194078 46170
rect 193458 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 194078 46102
rect 193458 45978 194078 46046
rect 193458 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 194078 45978
rect 193458 28350 194078 45922
rect 193458 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 194078 28350
rect 193458 28226 194078 28294
rect 193458 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 194078 28226
rect 193458 28102 194078 28170
rect 193458 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 194078 28102
rect 193458 27978 194078 28046
rect 193458 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 194078 27978
rect 193458 10350 194078 27922
rect 193458 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 194078 10350
rect 193458 10226 194078 10294
rect 193458 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 194078 10226
rect 193458 10102 194078 10170
rect 193458 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 194078 10102
rect 193458 9978 194078 10046
rect 193458 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 194078 9978
rect 193458 -1120 194078 9922
rect 209132 47998 209188 48008
rect 209132 4676 209188 47942
rect 209132 4610 209188 4620
rect 220458 40350 221078 48802
rect 220458 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 221078 40350
rect 220458 40226 221078 40294
rect 220458 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 221078 40226
rect 220458 40102 221078 40170
rect 220458 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 221078 40102
rect 220458 39978 221078 40046
rect 220458 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 221078 39978
rect 220458 22350 221078 39922
rect 220458 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 221078 22350
rect 220458 22226 221078 22294
rect 220458 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 221078 22226
rect 220458 22102 221078 22170
rect 220458 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 221078 22102
rect 220458 21978 221078 22046
rect 220458 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 221078 21978
rect 193458 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 194078 -1120
rect 193458 -1244 194078 -1176
rect 193458 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 194078 -1244
rect 193458 -1368 194078 -1300
rect 193458 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 194078 -1368
rect 193458 -1492 194078 -1424
rect 193458 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 194078 -1492
rect 193458 -1644 194078 -1548
rect 220458 4350 221078 21922
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 220458 4102 221078 4170
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 224178 46350 224798 48802
rect 224178 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 224798 46350
rect 224178 46226 224798 46294
rect 224178 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 224798 46226
rect 224178 46102 224798 46170
rect 224178 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 224798 46102
rect 224178 45978 224798 46046
rect 224178 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 224798 45978
rect 224178 28350 224798 45922
rect 224178 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 224798 28350
rect 224178 28226 224798 28294
rect 224178 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 224798 28226
rect 224178 28102 224798 28170
rect 224178 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 224798 28102
rect 224178 27978 224798 28046
rect 224178 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 224798 27978
rect 224178 10350 224798 27922
rect 224178 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 224798 10350
rect 224178 10226 224798 10294
rect 224178 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 224798 10226
rect 224178 10102 224798 10170
rect 224178 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 224798 10102
rect 224178 9978 224798 10046
rect 224178 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 224798 9978
rect 224178 -1120 224798 9922
rect 224178 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 224798 -1120
rect 224178 -1244 224798 -1176
rect 224178 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 224798 -1244
rect 224178 -1368 224798 -1300
rect 224178 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 224798 -1368
rect 224178 -1492 224798 -1424
rect 224178 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 224798 -1492
rect 224178 -1644 224798 -1548
rect 251178 40350 251798 48802
rect 251178 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 251798 40350
rect 251178 40226 251798 40294
rect 251178 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 251798 40226
rect 251178 40102 251798 40170
rect 251178 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 251798 40102
rect 251178 39978 251798 40046
rect 251178 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 251798 39978
rect 251178 22350 251798 39922
rect 251178 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 251798 22350
rect 251178 22226 251798 22294
rect 251178 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 251798 22226
rect 251178 22102 251798 22170
rect 251178 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 251798 22102
rect 251178 21978 251798 22046
rect 251178 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 251798 21978
rect 251178 4350 251798 21922
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 251178 4102 251798 4170
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 251178 -160 251798 3922
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 254898 46350 255518 48802
rect 254898 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 255518 46350
rect 254898 46226 255518 46294
rect 254898 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 255518 46226
rect 254898 46102 255518 46170
rect 254898 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 255518 46102
rect 254898 45978 255518 46046
rect 254898 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 255518 45978
rect 254898 28350 255518 45922
rect 266812 45108 266868 235004
rect 267148 234388 267204 234398
rect 267148 48804 267204 234332
rect 267148 48738 267204 48748
rect 266812 45042 266868 45052
rect 254898 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 255518 28350
rect 254898 28226 255518 28294
rect 254898 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 255518 28226
rect 254898 28102 255518 28170
rect 254898 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 255518 28102
rect 254898 27978 255518 28046
rect 254898 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 255518 27978
rect 254898 10350 255518 27922
rect 267260 17668 267316 238364
rect 268716 237076 268772 237086
rect 268604 236964 268660 236974
rect 267484 235172 267540 235182
rect 267372 234276 267428 234286
rect 267372 45332 267428 234220
rect 267372 45266 267428 45276
rect 267484 45220 267540 235116
rect 267596 230916 267652 230926
rect 267596 48468 267652 230860
rect 268604 136918 268660 236908
rect 268604 136852 268660 136862
rect 268716 133498 268772 237020
rect 270284 237076 270340 237086
rect 269276 234612 269332 234622
rect 269276 215068 269332 234556
rect 269612 231700 269668 231710
rect 269052 215012 269332 215068
rect 269500 224196 269556 224206
rect 269052 196678 269108 215012
rect 269164 208740 269220 208750
rect 269164 202258 269220 208684
rect 269164 202202 269444 202258
rect 269052 196622 269332 196678
rect 268716 133432 268772 133442
rect 267596 48402 267652 48412
rect 269276 48020 269332 196622
rect 269388 140084 269444 202202
rect 269388 140018 269444 140028
rect 269500 49700 269556 224140
rect 269500 49634 269556 49644
rect 269276 47954 269332 47964
rect 267484 45154 267540 45164
rect 269612 44772 269668 231644
rect 269612 44706 269668 44716
rect 269724 231418 269780 231428
rect 269724 44548 269780 231362
rect 269836 227818 269892 227828
rect 269836 49588 269892 227762
rect 270284 197428 270340 237020
rect 270284 197362 270340 197372
rect 270396 236964 270452 236974
rect 270396 161812 270452 236908
rect 270396 161746 270452 161756
rect 270508 234478 270564 234488
rect 269836 49522 269892 49532
rect 269724 44482 269780 44492
rect 270508 41188 270564 234422
rect 270844 231238 270900 231248
rect 270732 228452 270788 228462
rect 270508 41122 270564 41132
rect 270620 227556 270676 227566
rect 270620 38052 270676 227500
rect 270732 41300 270788 228396
rect 270844 48132 270900 231182
rect 272524 219828 272580 219838
rect 271068 218148 271124 218158
rect 270956 216580 271012 216590
rect 270956 154644 271012 216524
rect 271068 163380 271124 218092
rect 272188 214788 272244 214798
rect 272188 210980 272244 214732
rect 272412 213220 272468 213230
rect 272188 210914 272244 210924
rect 272300 212884 272356 212894
rect 272188 209636 272244 209646
rect 272188 204148 272244 209580
rect 272300 207060 272356 212828
rect 272412 211316 272468 213164
rect 272412 211250 272468 211260
rect 272300 206994 272356 207004
rect 272412 211092 272468 211102
rect 272188 204082 272244 204092
rect 272412 203308 272468 211036
rect 272524 209188 272580 219772
rect 272636 211204 272692 211214
rect 272636 209972 272692 211148
rect 272636 209906 272692 209916
rect 272524 209122 272580 209132
rect 272412 203252 272580 203308
rect 272524 189588 272580 203252
rect 272748 192500 272804 239260
rect 272860 219716 272916 219726
rect 272860 198324 272916 219660
rect 272860 198258 272916 198268
rect 272972 212996 273028 213006
rect 272972 195412 273028 212940
rect 273420 212772 273476 212782
rect 273196 210532 273252 210542
rect 272972 195346 273028 195356
rect 273084 209748 273140 209758
rect 272748 192434 272804 192444
rect 272524 189522 272580 189532
rect 273084 183764 273140 209692
rect 273196 186676 273252 210476
rect 273196 186610 273252 186620
rect 273308 205828 273364 205838
rect 273084 183698 273140 183708
rect 271068 163314 271124 163324
rect 270956 154578 271012 154588
rect 272524 153658 272580 153674
rect 272524 153570 272580 153580
rect 273308 110964 273364 205772
rect 273420 201236 273476 212716
rect 273420 201170 273476 201180
rect 273868 157556 273924 241276
rect 275548 237178 275604 237188
rect 274092 221172 274148 221182
rect 273868 157490 273924 157500
rect 273980 211764 274036 211774
rect 273980 154308 274036 211708
rect 274092 169204 274148 221116
rect 274092 169138 274148 169148
rect 274652 215908 274708 215918
rect 273980 154242 274036 154252
rect 273308 110898 273364 110908
rect 270844 48066 270900 48076
rect 270732 41234 270788 41244
rect 270620 37986 270676 37996
rect 274652 24612 274708 215852
rect 275436 154532 275492 154542
rect 275436 154308 275492 154476
rect 275436 154242 275492 154252
rect 274652 24546 274708 24556
rect 267260 17602 267316 17612
rect 254898 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 255518 10350
rect 254898 10226 255518 10294
rect 254898 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 255518 10226
rect 254898 10102 255518 10170
rect 254898 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 255518 10102
rect 254898 9978 255518 10046
rect 254898 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 255518 9978
rect 254898 -1120 255518 9922
rect 275548 7588 275604 237122
rect 275660 236998 275716 237008
rect 275660 26068 275716 236942
rect 275884 218036 275940 218046
rect 275772 216468 275828 216478
rect 275772 148820 275828 216412
rect 275884 166292 275940 217980
rect 275884 166226 275940 166236
rect 278012 150418 278068 241982
rect 322588 241444 322644 241454
rect 318556 241332 318612 241342
rect 278908 241220 278964 241230
rect 278908 151732 278964 241164
rect 288204 241220 288260 241230
rect 281372 240598 281428 240608
rect 278908 151666 278964 151676
rect 279692 239338 279748 239348
rect 278012 150352 278068 150362
rect 275772 148754 275828 148764
rect 279692 90580 279748 239282
rect 279692 90514 279748 90524
rect 275660 26002 275716 26012
rect 275548 7522 275604 7532
rect 281372 4452 281428 240542
rect 281372 4386 281428 4396
rect 281898 238350 282518 241154
rect 284956 240778 285012 240788
rect 281898 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 282518 238350
rect 281898 238226 282518 238294
rect 281898 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 282518 238226
rect 281898 238102 282518 238170
rect 281898 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 282518 238102
rect 281898 237978 282518 238046
rect 281898 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 282518 237978
rect 281898 220350 282518 237922
rect 284732 240418 284788 240428
rect 281898 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 282518 220350
rect 281898 220226 282518 220294
rect 281898 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 282518 220226
rect 281898 220102 282518 220170
rect 281898 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 282518 220102
rect 281898 219978 282518 220046
rect 281898 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 282518 219978
rect 281898 202350 282518 219922
rect 281898 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 282518 202350
rect 281898 202226 282518 202294
rect 281898 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 282518 202226
rect 281898 202102 282518 202170
rect 281898 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 282518 202102
rect 281898 201978 282518 202046
rect 281898 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 282518 201978
rect 281898 184350 282518 201922
rect 281898 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 282518 184350
rect 281898 184226 282518 184294
rect 281898 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 282518 184226
rect 281898 184102 282518 184170
rect 281898 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 282518 184102
rect 281898 183978 282518 184046
rect 281898 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 282518 183978
rect 281898 166350 282518 183922
rect 281898 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 282518 166350
rect 281898 166226 282518 166294
rect 281898 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 282518 166226
rect 281898 166102 282518 166170
rect 281898 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 282518 166102
rect 281898 165978 282518 166046
rect 281898 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 282518 165978
rect 281898 148350 282518 165922
rect 281898 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 282518 148350
rect 281898 148226 282518 148294
rect 281898 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 282518 148226
rect 281898 148102 282518 148170
rect 281898 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 282518 148102
rect 281898 147978 282518 148046
rect 281898 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 282518 147978
rect 281898 130350 282518 147922
rect 281898 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 282518 130350
rect 281898 130226 282518 130294
rect 281898 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 282518 130226
rect 281898 130102 282518 130170
rect 281898 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 282518 130102
rect 281898 129978 282518 130046
rect 281898 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 282518 129978
rect 281898 112350 282518 129922
rect 281898 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 282518 112350
rect 281898 112226 282518 112294
rect 281898 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 282518 112226
rect 281898 112102 282518 112170
rect 281898 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 282518 112102
rect 281898 111978 282518 112046
rect 281898 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 282518 111978
rect 281898 94350 282518 111922
rect 281898 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 282518 94350
rect 281898 94226 282518 94294
rect 281898 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 282518 94226
rect 281898 94102 282518 94170
rect 281898 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 282518 94102
rect 281898 93978 282518 94046
rect 281898 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 282518 93978
rect 281898 76350 282518 93922
rect 281898 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 282518 76350
rect 281898 76226 282518 76294
rect 281898 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 282518 76226
rect 281898 76102 282518 76170
rect 281898 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 282518 76102
rect 281898 75978 282518 76046
rect 281898 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 282518 75978
rect 281898 58350 282518 75922
rect 281898 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 282518 58350
rect 281898 58226 282518 58294
rect 281898 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 282518 58226
rect 281898 58102 282518 58170
rect 281898 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 282518 58102
rect 281898 57978 282518 58046
rect 281898 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 282518 57978
rect 281898 40350 282518 57922
rect 281898 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 282518 40350
rect 281898 40226 282518 40294
rect 281898 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 282518 40226
rect 281898 40102 282518 40170
rect 281898 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 282518 40102
rect 281898 39978 282518 40046
rect 281898 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 282518 39978
rect 281898 22350 282518 39922
rect 281898 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 282518 22350
rect 281898 22226 282518 22294
rect 281898 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 282518 22226
rect 281898 22102 282518 22170
rect 281898 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 282518 22102
rect 281898 21978 282518 22046
rect 281898 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 282518 21978
rect 254898 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 255518 -1120
rect 254898 -1244 255518 -1176
rect 254898 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 255518 -1244
rect 254898 -1368 255518 -1300
rect 254898 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 255518 -1368
rect 254898 -1492 255518 -1424
rect 254898 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 255518 -1492
rect 254898 -1644 255518 -1548
rect 281898 4350 282518 21922
rect 283052 234478 283108 234488
rect 283052 4564 283108 234422
rect 284732 4798 284788 240362
rect 284732 4732 284788 4742
rect 283052 4498 283108 4508
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 281898 4226 282518 4294
rect 284956 4340 285012 240722
rect 285180 236098 285236 236108
rect 285180 4788 285236 236042
rect 285180 4722 285236 4732
rect 285618 226350 286238 241154
rect 288204 239316 288260 241164
rect 304892 240772 304948 240782
rect 304892 239428 304948 240716
rect 304892 239362 304948 239372
rect 288204 239250 288260 239260
rect 312618 238350 313238 241154
rect 314972 240100 315028 240110
rect 314972 239428 315028 240044
rect 314972 239362 315028 239372
rect 312618 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 313238 238350
rect 312618 238226 313238 238294
rect 312618 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 313238 238226
rect 312618 238102 313238 238170
rect 312618 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 313238 238102
rect 312618 237978 313238 238046
rect 312618 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 313238 237978
rect 293916 237076 293972 237086
rect 285618 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 286238 226350
rect 285618 226226 286238 226294
rect 285618 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 286238 226226
rect 285618 226102 286238 226170
rect 285618 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 286238 226102
rect 285618 225978 286238 226046
rect 285618 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 286238 225978
rect 285618 208350 286238 225922
rect 293804 236964 293860 236974
rect 289772 214498 289828 214508
rect 285618 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 286238 208350
rect 285618 208226 286238 208294
rect 285618 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 286238 208226
rect 285618 208102 286238 208170
rect 285618 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 286238 208102
rect 285618 207978 286238 208046
rect 285618 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 286238 207978
rect 285618 190350 286238 207922
rect 285618 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 286238 190350
rect 285618 190226 286238 190294
rect 285618 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 286238 190226
rect 285618 190102 286238 190170
rect 285618 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 286238 190102
rect 285618 189978 286238 190046
rect 285618 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 286238 189978
rect 285618 172350 286238 189922
rect 285618 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 286238 172350
rect 285618 172226 286238 172294
rect 285618 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 286238 172226
rect 285618 172102 286238 172170
rect 285618 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 286238 172102
rect 285618 171978 286238 172046
rect 285618 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 286238 171978
rect 285618 154350 286238 171922
rect 285618 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 286238 154350
rect 285618 154226 286238 154294
rect 285618 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 286238 154226
rect 285618 154102 286238 154170
rect 285618 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 286238 154102
rect 285618 153978 286238 154046
rect 285618 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 286238 153978
rect 285618 136350 286238 153922
rect 285618 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 286238 136350
rect 285618 136226 286238 136294
rect 285618 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 286238 136226
rect 285618 136102 286238 136170
rect 285618 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 286238 136102
rect 285618 135978 286238 136046
rect 285618 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 286238 135978
rect 285618 118350 286238 135922
rect 285618 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 286238 118350
rect 285618 118226 286238 118294
rect 285618 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 286238 118226
rect 285618 118102 286238 118170
rect 285618 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 286238 118102
rect 285618 117978 286238 118046
rect 285618 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 286238 117978
rect 285618 100350 286238 117922
rect 285618 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 286238 100350
rect 285618 100226 286238 100294
rect 285618 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 286238 100226
rect 285618 100102 286238 100170
rect 285618 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 286238 100102
rect 285618 99978 286238 100046
rect 285618 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 286238 99978
rect 285618 82350 286238 99922
rect 285618 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 286238 82350
rect 285618 82226 286238 82294
rect 285618 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 286238 82226
rect 285618 82102 286238 82170
rect 285618 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 286238 82102
rect 285618 81978 286238 82046
rect 285618 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 286238 81978
rect 285618 64350 286238 81922
rect 285618 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 286238 64350
rect 285618 64226 286238 64294
rect 285618 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 286238 64226
rect 285618 64102 286238 64170
rect 285618 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 286238 64102
rect 285618 63978 286238 64046
rect 285618 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 286238 63978
rect 285618 46350 286238 63922
rect 285618 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 286238 46350
rect 285618 46226 286238 46294
rect 285618 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 286238 46226
rect 285618 46102 286238 46170
rect 285618 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 286238 46102
rect 285618 45978 286238 46046
rect 285618 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 286238 45978
rect 285618 28350 286238 45922
rect 285618 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 286238 28350
rect 285618 28226 286238 28294
rect 285618 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 286238 28226
rect 285618 28102 286238 28170
rect 285618 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 286238 28102
rect 285618 27978 286238 28046
rect 285618 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 286238 27978
rect 285618 10350 286238 27922
rect 285618 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 286238 10350
rect 285618 10226 286238 10294
rect 285618 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 286238 10226
rect 285618 10102 286238 10170
rect 285618 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 286238 10102
rect 285618 9978 286238 10046
rect 285618 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 286238 9978
rect 284956 4274 285012 4284
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 281898 4102 282518 4170
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 281898 -160 282518 3922
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 285618 -1120 286238 9922
rect 288092 211438 288148 211448
rect 288092 7140 288148 211382
rect 289772 52052 289828 214442
rect 293804 160498 293860 236908
rect 293804 160432 293860 160442
rect 293916 158698 293972 237020
rect 293916 158632 293972 158642
rect 295596 236964 295652 236974
rect 295596 155458 295652 236908
rect 298956 236964 299012 236974
rect 295596 155392 295652 155402
rect 298172 214116 298228 214126
rect 298172 124318 298228 214060
rect 298956 160678 299012 236908
rect 298956 160612 299012 160622
rect 300636 236964 300692 236974
rect 300636 158878 300692 236908
rect 306572 236628 306628 236638
rect 300636 158812 300692 158822
rect 304892 226548 304948 226558
rect 298172 124252 298228 124262
rect 304892 124138 304948 226492
rect 304892 124072 304948 124082
rect 306572 123958 306628 236572
rect 307356 236068 307412 236078
rect 306572 123892 306628 123902
rect 306796 229460 306852 229470
rect 306796 123598 306852 229404
rect 307356 146098 307412 236012
rect 312396 231700 312452 231710
rect 311724 231588 311780 231598
rect 311612 231058 311668 231068
rect 309932 229572 309988 229582
rect 307356 145460 307412 146042
rect 307356 145394 307412 145404
rect 307468 216244 307524 216254
rect 306796 123532 306852 123542
rect 299500 82147 299820 82204
rect 299500 82091 299528 82147
rect 299584 82091 299632 82147
rect 299688 82091 299736 82147
rect 299792 82091 299820 82147
rect 299500 82043 299820 82091
rect 299500 81987 299528 82043
rect 299584 81987 299632 82043
rect 299688 81987 299736 82043
rect 299792 81987 299820 82043
rect 299500 81939 299820 81987
rect 299500 81883 299528 81939
rect 299584 81883 299632 81939
rect 299688 81883 299736 81939
rect 299792 81883 299820 81939
rect 299500 81826 299820 81883
rect 295342 76350 295662 76384
rect 295342 76294 295412 76350
rect 295468 76294 295536 76350
rect 295592 76294 295662 76350
rect 295342 76226 295662 76294
rect 295342 76170 295412 76226
rect 295468 76170 295536 76226
rect 295592 76170 295662 76226
rect 295342 76102 295662 76170
rect 295342 76046 295412 76102
rect 295468 76046 295536 76102
rect 295592 76046 295662 76102
rect 295342 75978 295662 76046
rect 295342 75922 295412 75978
rect 295468 75922 295536 75978
rect 295592 75922 295662 75978
rect 295342 75888 295662 75922
rect 303658 76350 303978 76384
rect 303658 76294 303728 76350
rect 303784 76294 303852 76350
rect 303908 76294 303978 76350
rect 303658 76226 303978 76294
rect 303658 76170 303728 76226
rect 303784 76170 303852 76226
rect 303908 76170 303978 76226
rect 303658 76102 303978 76170
rect 303658 76046 303728 76102
rect 303784 76046 303852 76102
rect 303908 76046 303978 76102
rect 303658 75978 303978 76046
rect 303658 75922 303728 75978
rect 303784 75922 303852 75978
rect 303908 75922 303978 75978
rect 303658 75888 303978 75922
rect 299500 64350 299820 64384
rect 299500 64294 299570 64350
rect 299626 64294 299694 64350
rect 299750 64294 299820 64350
rect 299500 64226 299820 64294
rect 299500 64170 299570 64226
rect 299626 64170 299694 64226
rect 299750 64170 299820 64226
rect 299500 64102 299820 64170
rect 299500 64046 299570 64102
rect 299626 64046 299694 64102
rect 299750 64046 299820 64102
rect 299500 63978 299820 64046
rect 299500 63922 299570 63978
rect 299626 63922 299694 63978
rect 299750 63922 299820 63978
rect 299500 63888 299820 63922
rect 295342 58350 295662 58384
rect 295342 58294 295412 58350
rect 295468 58294 295536 58350
rect 295592 58294 295662 58350
rect 295342 58226 295662 58294
rect 295342 58170 295412 58226
rect 295468 58170 295536 58226
rect 295592 58170 295662 58226
rect 295342 58102 295662 58170
rect 295342 58046 295412 58102
rect 295468 58046 295536 58102
rect 295592 58046 295662 58102
rect 295342 57978 295662 58046
rect 295342 57922 295412 57978
rect 295468 57922 295536 57978
rect 295592 57922 295662 57978
rect 295342 57888 295662 57922
rect 303658 58350 303978 58384
rect 303658 58294 303728 58350
rect 303784 58294 303852 58350
rect 303908 58294 303978 58350
rect 303658 58226 303978 58294
rect 303658 58170 303728 58226
rect 303784 58170 303852 58226
rect 303908 58170 303978 58226
rect 303658 58102 303978 58170
rect 303658 58046 303728 58102
rect 303784 58046 303852 58102
rect 303908 58046 303978 58102
rect 303658 57978 303978 58046
rect 303658 57922 303728 57978
rect 303784 57922 303852 57978
rect 303908 57922 303978 57978
rect 303658 57888 303978 57922
rect 289772 51986 289828 51996
rect 307468 50372 307524 216188
rect 308252 211428 308308 211438
rect 308252 123778 308308 211372
rect 308252 123712 308308 123722
rect 307816 82147 308136 82204
rect 307816 82091 307844 82147
rect 307900 82091 307948 82147
rect 308004 82091 308052 82147
rect 308108 82091 308136 82147
rect 307816 82043 308136 82091
rect 307816 81987 307844 82043
rect 307900 81987 307948 82043
rect 308004 81987 308052 82043
rect 308108 81987 308136 82043
rect 307816 81939 308136 81987
rect 307816 81883 307844 81939
rect 307900 81883 307948 81939
rect 308004 81883 308052 81939
rect 308108 81883 308136 81939
rect 307816 81826 308136 81883
rect 307816 64350 308136 64384
rect 307816 64294 307886 64350
rect 307942 64294 308010 64350
rect 308066 64294 308136 64350
rect 307816 64226 308136 64294
rect 307816 64170 307886 64226
rect 307942 64170 308010 64226
rect 308066 64170 308136 64226
rect 307816 64102 308136 64170
rect 307816 64046 307886 64102
rect 307942 64046 308010 64102
rect 308066 64046 308136 64102
rect 307816 63978 308136 64046
rect 307816 63922 307886 63978
rect 307942 63922 308010 63978
rect 308066 63922 308136 63978
rect 307816 63888 308136 63922
rect 307468 50306 307524 50316
rect 309932 27748 309988 229516
rect 311612 37940 311668 231002
rect 311724 47818 311780 231532
rect 311948 231364 312004 231374
rect 311724 47752 311780 47762
rect 311836 230698 311892 230708
rect 311612 37874 311668 37884
rect 311836 37828 311892 230642
rect 311948 108052 312004 231308
rect 312060 230518 312116 230528
rect 312060 113876 312116 230462
rect 312060 113810 312116 113820
rect 311948 107986 312004 107996
rect 311974 76350 312294 76384
rect 311974 76294 312044 76350
rect 312100 76294 312168 76350
rect 312224 76294 312294 76350
rect 311974 76226 312294 76294
rect 311974 76170 312044 76226
rect 312100 76170 312168 76226
rect 312224 76170 312294 76226
rect 311974 76102 312294 76170
rect 311974 76046 312044 76102
rect 312100 76046 312168 76102
rect 312224 76046 312294 76102
rect 311974 75978 312294 76046
rect 311974 75922 312044 75978
rect 312100 75922 312168 75978
rect 312224 75922 312294 75978
rect 311974 75888 312294 75922
rect 311974 58350 312294 58384
rect 311974 58294 312044 58350
rect 312100 58294 312168 58350
rect 312224 58294 312294 58350
rect 311974 58226 312294 58294
rect 311974 58170 312044 58226
rect 312100 58170 312168 58226
rect 312224 58170 312294 58226
rect 311974 58102 312294 58170
rect 311974 58046 312044 58102
rect 312100 58046 312168 58102
rect 312224 58046 312294 58102
rect 311974 57978 312294 58046
rect 311974 57922 312044 57978
rect 312100 57922 312168 57978
rect 312224 57922 312294 57978
rect 311974 57888 312294 57922
rect 312396 47998 312452 231644
rect 312396 47932 312452 47942
rect 312618 220350 313238 237922
rect 312618 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 313238 220350
rect 312618 220226 313238 220294
rect 312618 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 313238 220226
rect 312618 220102 313238 220170
rect 312618 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 313238 220102
rect 312618 219978 313238 220046
rect 312618 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 313238 219978
rect 312618 202350 313238 219922
rect 312618 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 313238 202350
rect 312618 202226 313238 202294
rect 312618 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 313238 202226
rect 312618 202102 313238 202170
rect 312618 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 313238 202102
rect 312618 201978 313238 202046
rect 312618 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 313238 201978
rect 312618 184350 313238 201922
rect 314860 239204 314916 239214
rect 312618 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 313238 184350
rect 312618 184226 313238 184294
rect 312618 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 313238 184226
rect 312618 184102 313238 184170
rect 312618 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 313238 184102
rect 312618 183978 313238 184046
rect 312618 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 313238 183978
rect 312618 166350 313238 183922
rect 312618 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 313238 166350
rect 312618 166226 313238 166294
rect 312618 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 313238 166226
rect 312618 166102 313238 166170
rect 312618 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 313238 166102
rect 312618 165978 313238 166046
rect 312618 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 313238 165978
rect 312618 148350 313238 165922
rect 313404 194740 313460 194750
rect 313404 160692 313460 194684
rect 313404 160626 313460 160636
rect 314860 160132 314916 239148
rect 314860 160066 314916 160076
rect 314972 234658 315028 234668
rect 312618 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 313238 148350
rect 312618 148226 313238 148294
rect 312618 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 313238 148226
rect 312618 148102 313238 148170
rect 312618 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 313238 148102
rect 312618 147978 313238 148046
rect 312618 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 313238 147978
rect 312618 130350 313238 147922
rect 312618 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 313238 130350
rect 312618 130226 313238 130294
rect 312618 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 313238 130226
rect 312618 130102 313238 130170
rect 312618 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 313238 130102
rect 312618 129978 313238 130046
rect 312618 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 313238 129978
rect 312618 112350 313238 129922
rect 312618 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 313238 112350
rect 312618 112226 313238 112294
rect 312618 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 313238 112226
rect 312618 112102 313238 112170
rect 312618 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 313238 112102
rect 312618 111978 313238 112046
rect 312618 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 313238 111978
rect 312618 94350 313238 111922
rect 312618 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 313238 94350
rect 312618 94226 313238 94294
rect 312618 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 313238 94226
rect 312618 94102 313238 94170
rect 312618 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 313238 94102
rect 312618 93978 313238 94046
rect 312618 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 313238 93978
rect 312618 76350 313238 93922
rect 312618 76294 312714 76350
rect 312770 76294 312838 76350
rect 312894 76294 312962 76350
rect 313018 76294 313086 76350
rect 313142 76294 313238 76350
rect 312618 76226 313238 76294
rect 312618 76170 312714 76226
rect 312770 76170 312838 76226
rect 312894 76170 312962 76226
rect 313018 76170 313086 76226
rect 313142 76170 313238 76226
rect 312618 76102 313238 76170
rect 312618 76046 312714 76102
rect 312770 76046 312838 76102
rect 312894 76046 312962 76102
rect 313018 76046 313086 76102
rect 313142 76046 313238 76102
rect 312618 75978 313238 76046
rect 312618 75922 312714 75978
rect 312770 75922 312838 75978
rect 312894 75922 312962 75978
rect 313018 75922 313086 75978
rect 313142 75922 313238 75978
rect 312618 58350 313238 75922
rect 312618 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 313238 58350
rect 312618 58226 313238 58294
rect 312618 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 313238 58226
rect 312618 58102 313238 58170
rect 312618 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 313238 58102
rect 312618 57978 313238 58046
rect 312618 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 313238 57978
rect 311836 37762 311892 37772
rect 312618 40350 313238 57922
rect 312618 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 313238 40350
rect 312618 40226 313238 40294
rect 312618 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 313238 40226
rect 312618 40102 313238 40170
rect 312618 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 313238 40102
rect 312618 39978 313238 40046
rect 312618 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 313238 39978
rect 309932 27682 309988 27692
rect 288092 7074 288148 7084
rect 312618 22350 313238 39922
rect 312618 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 313238 22350
rect 312618 22226 313238 22294
rect 312618 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 313238 22226
rect 312618 22102 313238 22170
rect 312618 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 313238 22102
rect 312618 21978 313238 22046
rect 312618 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 313238 21978
rect 285618 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 286238 -1120
rect 285618 -1244 286238 -1176
rect 285618 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 286238 -1244
rect 285618 -1368 286238 -1300
rect 285618 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 286238 -1368
rect 285618 -1492 286238 -1424
rect 285618 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 286238 -1492
rect 285618 -1644 286238 -1548
rect 312618 4350 313238 21922
rect 314972 4978 315028 234602
rect 315196 234500 315252 234510
rect 315084 211258 315140 211268
rect 315084 48580 315140 211202
rect 315196 87668 315252 234444
rect 316338 226350 316958 241154
rect 317884 241108 317940 241118
rect 317884 240660 317940 241052
rect 317884 240594 317940 240604
rect 318556 240660 318612 241276
rect 318556 240594 318612 240604
rect 322588 240660 322644 241388
rect 322588 240594 322644 240604
rect 323260 240660 323316 242702
rect 334236 242038 334292 242048
rect 323260 240594 323316 240604
rect 334124 240996 334180 241006
rect 334124 240598 334180 240940
rect 334236 240772 334292 241982
rect 335804 241668 335860 253502
rect 335804 241602 335860 241612
rect 335916 241780 335972 241790
rect 334236 240706 334292 240716
rect 335916 240778 335972 241724
rect 335916 240712 335972 240722
rect 334124 240532 334180 240542
rect 320572 240238 320628 240250
rect 320572 240146 320628 240156
rect 319900 240100 319956 240110
rect 319900 239992 319956 240002
rect 316338 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 316958 226350
rect 316338 226226 316958 226294
rect 316338 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 316958 226226
rect 316338 226102 316958 226170
rect 316338 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 316958 226102
rect 316338 225978 316958 226046
rect 316338 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 316958 225978
rect 316338 208350 316958 225922
rect 316338 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 316958 208350
rect 316338 208226 316958 208294
rect 316338 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 316958 208226
rect 316338 208102 316958 208170
rect 316338 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 316958 208102
rect 316338 207978 316958 208046
rect 316338 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 316958 207978
rect 315196 87602 315252 87612
rect 315308 197652 315364 197662
rect 315308 50372 315364 197596
rect 316338 193230 316958 207922
rect 317436 239092 317492 239102
rect 317212 197876 317268 197886
rect 315468 184350 315788 184384
rect 315468 184294 315538 184350
rect 315594 184294 315662 184350
rect 315718 184294 315788 184350
rect 315468 184226 315788 184294
rect 315468 184170 315538 184226
rect 315594 184170 315662 184226
rect 315718 184170 315788 184226
rect 315468 184102 315788 184170
rect 315468 184046 315538 184102
rect 315594 184046 315662 184102
rect 315718 184046 315788 184102
rect 315468 183978 315788 184046
rect 315468 183922 315538 183978
rect 315594 183922 315662 183978
rect 315718 183922 315788 183978
rect 315468 183888 315788 183922
rect 317212 173068 317268 197820
rect 317100 173012 317268 173068
rect 317324 197764 317380 197774
rect 315468 166350 315788 166384
rect 315468 166294 315538 166350
rect 315594 166294 315662 166350
rect 315718 166294 315788 166350
rect 315468 166226 315788 166294
rect 315468 166170 315538 166226
rect 315594 166170 315662 166226
rect 315718 166170 315788 166226
rect 315468 166102 315788 166170
rect 315468 166046 315538 166102
rect 315594 166046 315662 166102
rect 315718 166046 315788 166102
rect 315468 165978 315788 166046
rect 315468 165922 315538 165978
rect 315594 165922 315662 165978
rect 315718 165922 315788 165978
rect 315468 165888 315788 165922
rect 316338 154350 316958 163170
rect 317100 157556 317156 173012
rect 317324 157780 317380 197708
rect 317436 160132 317492 239036
rect 321244 238532 321300 238542
rect 321244 237718 321300 238476
rect 321244 237652 321300 237662
rect 321916 238532 321972 238542
rect 321916 237538 321972 238476
rect 321916 237472 321972 237482
rect 320012 231252 320068 231262
rect 320012 230698 320068 231196
rect 320012 230632 320068 230642
rect 329196 231140 329252 231150
rect 329196 230338 329252 231084
rect 329196 230272 329252 230282
rect 336028 194740 336084 368702
rect 336700 304858 336756 304868
rect 336588 241678 336644 241688
rect 336588 224420 336644 241622
rect 336588 224354 336644 224364
rect 336700 197988 336756 304802
rect 336812 253018 336868 379484
rect 336924 308998 336980 380492
rect 338268 368758 338324 368768
rect 336924 308932 336980 308942
rect 338156 336358 338212 336368
rect 336812 252952 336868 252962
rect 336924 284698 336980 284708
rect 336812 241858 336868 241868
rect 336812 222852 336868 241802
rect 336924 240548 336980 284642
rect 337260 279658 337316 279668
rect 336924 240482 336980 240492
rect 337036 277318 337092 277328
rect 337036 239988 337092 277262
rect 337036 239922 337092 239932
rect 337148 267238 337204 267248
rect 337148 231588 337204 267182
rect 337260 253558 337316 279602
rect 337260 253492 337316 253502
rect 337372 257878 337428 257888
rect 337148 231522 337204 231532
rect 337260 244738 337316 244748
rect 337260 226324 337316 244682
rect 337372 231700 337428 257822
rect 337484 254818 337540 254828
rect 337484 234658 337540 254762
rect 337596 246358 337652 246368
rect 337596 240324 337652 246302
rect 337708 241668 337764 241678
rect 337708 240418 337764 241612
rect 337708 240352 337764 240362
rect 337596 240258 337652 240268
rect 337484 234592 337540 234602
rect 337372 231634 337428 231644
rect 337260 226258 337316 226268
rect 336812 222786 336868 222796
rect 336700 197922 336756 197932
rect 338156 197316 338212 336302
rect 338268 250348 338324 368702
rect 338492 325948 338548 385756
rect 339276 337708 339332 408940
rect 343338 400350 343958 410034
rect 343338 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 343958 400350
rect 343338 400226 343958 400294
rect 343338 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 343958 400226
rect 343338 400102 343958 400170
rect 343338 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 343958 400102
rect 343338 399978 343958 400046
rect 343338 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 343958 399978
rect 341964 392338 342020 392348
rect 340060 383236 340116 383246
rect 339164 337652 339332 337708
rect 339948 368004 340004 368014
rect 339164 337438 339220 337652
rect 339164 337382 339444 337438
rect 339276 337316 339332 337326
rect 339276 337078 339332 337260
rect 338940 337022 339332 337078
rect 338492 325892 338884 325948
rect 338828 313318 338884 325892
rect 338828 313252 338884 313262
rect 338940 267148 338996 337022
rect 339388 336718 339444 337382
rect 339276 336662 339444 336718
rect 339276 325948 339332 336662
rect 339388 336420 339444 336430
rect 339388 336358 339444 336364
rect 339388 336292 339444 336302
rect 339052 325892 339332 325948
rect 339052 309898 339108 325892
rect 339276 318500 339332 318510
rect 339276 310078 339332 318444
rect 339388 313348 339444 313358
rect 339388 313252 339444 313262
rect 339276 310022 339444 310078
rect 339052 309876 339332 309898
rect 339052 309842 339276 309876
rect 339276 309810 339332 309820
rect 339388 309358 339444 310022
rect 339164 309302 339444 309358
rect 339500 309876 339556 309886
rect 339164 302428 339220 309302
rect 339500 305788 339556 309820
rect 339276 305732 339556 305788
rect 339276 305218 339332 305732
rect 339276 305162 339444 305218
rect 339276 305060 339332 305070
rect 339276 304966 339332 304982
rect 339388 304858 339444 305162
rect 339052 302372 339220 302428
rect 339276 304802 339444 304858
rect 339052 285628 339108 302372
rect 339276 288932 339332 304802
rect 339276 288866 339332 288876
rect 339612 303268 339668 303278
rect 339052 285572 339332 285628
rect 339276 281818 339332 285572
rect 339388 284788 339444 284798
rect 339388 284698 339444 284732
rect 339388 284632 339444 284642
rect 339276 281762 339556 281818
rect 339276 281204 339332 281214
rect 339276 280738 339332 281148
rect 339500 280918 339556 281762
rect 338604 267092 338996 267148
rect 339052 280682 339332 280738
rect 339388 280862 339556 280918
rect 338604 262108 338660 267092
rect 339052 264538 339108 280682
rect 339388 280558 339444 280862
rect 339164 280502 339444 280558
rect 339164 270508 339220 280502
rect 339276 280196 339332 280206
rect 339276 277318 339332 280140
rect 339388 279658 339444 279668
rect 339388 279564 339444 279580
rect 339276 277252 339332 277262
rect 339164 270452 339556 270508
rect 339276 270116 339332 270126
rect 339332 270060 339444 270116
rect 339276 270050 339332 270060
rect 339276 267428 339332 267438
rect 339276 267334 339332 267362
rect 339052 264482 339332 264538
rect 338380 262052 338660 262108
rect 338716 264358 338772 264368
rect 338380 254638 338436 262052
rect 338604 258778 338660 258788
rect 338380 254572 338436 254582
rect 338492 258722 338604 258778
rect 338268 250292 338436 250348
rect 338268 248698 338324 248708
rect 338268 240548 338324 248642
rect 338268 240482 338324 240492
rect 338380 239988 338436 250292
rect 338380 239338 338436 239932
rect 338380 239272 338436 239282
rect 338492 238588 338548 258722
rect 338604 258712 338660 258722
rect 338716 256258 338772 264302
rect 339276 264178 339332 264482
rect 339388 264358 339444 270060
rect 339388 264292 339444 264302
rect 338828 264122 339332 264178
rect 338828 258748 338884 264122
rect 339500 260578 339556 270452
rect 339164 260522 339556 260578
rect 338828 258692 339108 258748
rect 338716 256202 338996 256258
rect 338828 255718 338884 255728
rect 338604 255662 338828 255718
rect 338604 250348 338660 255662
rect 338828 255652 338884 255662
rect 338940 250348 338996 256202
rect 338604 250292 338772 250348
rect 338380 238532 338548 238588
rect 338604 241892 338660 241902
rect 338380 226436 338436 238532
rect 338380 226370 338436 226380
rect 338604 219828 338660 241836
rect 338716 226212 338772 250292
rect 338716 226146 338772 226156
rect 338828 250292 338996 250348
rect 338604 219762 338660 219772
rect 338828 219716 338884 250292
rect 338940 248878 338996 248888
rect 338940 229572 338996 248822
rect 339052 248698 339108 258692
rect 339164 248698 339220 260522
rect 339276 260260 339332 260270
rect 339276 255718 339332 260204
rect 339276 255652 339332 255662
rect 339388 260036 339444 260046
rect 339276 254884 339332 254894
rect 339276 254818 339332 254828
rect 339276 254752 339332 254762
rect 339276 254638 339332 254648
rect 339276 252532 339332 254582
rect 339276 252466 339332 252476
rect 339276 250404 339332 250414
rect 339276 248878 339332 250348
rect 339388 250348 339444 259980
rect 339500 258804 339556 258814
rect 339500 258710 339556 258722
rect 339500 257908 339556 257918
rect 339500 257812 339556 257822
rect 339388 250292 339556 250348
rect 339276 248812 339332 248822
rect 339164 248642 339444 248698
rect 339052 248632 339108 248642
rect 339388 248338 339444 248642
rect 339164 248282 339444 248338
rect 339164 238588 339220 248282
rect 339276 247156 339332 247166
rect 339276 241892 339332 247100
rect 339388 246372 339444 246382
rect 339388 246278 339444 246302
rect 339276 241826 339332 241836
rect 339500 241858 339556 250292
rect 339500 241792 339556 241802
rect 339164 238532 339332 238588
rect 338940 229506 338996 229516
rect 338828 219650 338884 219660
rect 338156 197250 338212 197260
rect 336028 194674 336084 194684
rect 339276 193258 339332 238532
rect 339612 197092 339668 303212
rect 339724 275492 339780 275502
rect 339724 227638 339780 275436
rect 339836 274596 339892 274606
rect 339836 229348 339892 274540
rect 339836 229282 339892 229292
rect 339724 227572 339780 227582
rect 339612 197026 339668 197036
rect 339948 193978 340004 367948
rect 340060 197652 340116 383180
rect 340284 373798 340340 373808
rect 340172 359604 340228 359614
rect 340172 235172 340228 359548
rect 340172 235106 340228 235116
rect 340284 295764 340340 373742
rect 340284 231476 340340 295708
rect 341852 350756 341908 350766
rect 341292 287140 341348 287150
rect 341292 255892 341348 287084
rect 341180 255780 341236 255790
rect 340396 251300 340452 251310
rect 340396 241678 340452 251244
rect 341180 244738 341236 255724
rect 341180 244672 341236 244682
rect 340396 241612 340452 241622
rect 341292 239876 341348 255836
rect 341292 239810 341348 239820
rect 341404 278180 341460 278190
rect 341404 239698 341460 278124
rect 341740 277284 341796 277294
rect 341068 239652 341460 239698
rect 341124 239642 341460 239652
rect 341516 276388 341572 276398
rect 341068 238644 341124 239596
rect 341068 238578 341124 238588
rect 340284 231410 340340 231420
rect 341516 224218 341572 276332
rect 341516 224152 341572 224162
rect 341628 245924 341684 245934
rect 341628 222628 341684 245868
rect 341740 234298 341796 277228
rect 341740 234232 341796 234242
rect 341628 222562 341684 222572
rect 340060 197586 340116 197596
rect 339948 193912 340004 193922
rect 339276 193192 339332 193202
rect 341852 192538 341908 350700
rect 341964 237748 342020 392282
rect 342300 386036 342356 386046
rect 342076 373078 342132 373088
rect 342076 290724 342132 373022
rect 342300 325918 342356 385980
rect 343084 383908 343140 383918
rect 342972 379652 343028 379662
rect 342300 325852 342356 325862
rect 342860 378838 342916 378848
rect 342076 290658 342132 290668
rect 342188 314916 342244 314926
rect 342188 247828 342244 314860
rect 342412 297892 342468 297902
rect 342412 248500 342468 297836
rect 342748 292618 342804 292628
rect 342748 292516 342804 292562
rect 342748 292450 342804 292460
rect 342860 289828 342916 378782
rect 342972 344484 343028 379596
rect 342972 344418 343028 344428
rect 343084 290948 343140 383852
rect 343084 290882 343140 290892
rect 343338 382350 343958 399922
rect 347058 406350 347678 410034
rect 356188 408178 356244 408188
rect 356188 407428 356244 408122
rect 356188 407362 356244 407372
rect 357196 407092 357252 411002
rect 359884 410116 359940 410126
rect 358764 409978 358820 409988
rect 357196 406644 357252 407036
rect 357308 409618 357364 409628
rect 357308 407988 357364 409562
rect 358092 409438 358148 409448
rect 357308 406756 357364 407932
rect 357308 406690 357364 406700
rect 357644 409078 357700 409088
rect 357644 407638 357700 409022
rect 358092 408268 358148 409382
rect 357196 406578 357252 406588
rect 347058 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 347678 406350
rect 347058 406226 347678 406294
rect 347058 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 347678 406226
rect 347058 406102 347678 406170
rect 347058 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 347678 406102
rect 347058 405978 347678 406046
rect 347058 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 347678 405978
rect 343338 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 343958 382350
rect 343338 382226 343958 382294
rect 343338 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 343958 382226
rect 343338 382102 343958 382170
rect 343338 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 343958 382102
rect 343338 381978 343958 382046
rect 343338 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 343958 381978
rect 343338 364350 343958 381922
rect 344092 398278 344148 398288
rect 344092 373156 344148 398222
rect 345548 396658 345604 396668
rect 344092 373090 344148 373100
rect 344204 395398 344260 395408
rect 344204 372260 344260 395342
rect 344204 372194 344260 372204
rect 343338 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 343958 364350
rect 343338 364226 343958 364294
rect 343338 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 343958 364226
rect 343338 364102 343958 364170
rect 343338 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 343958 364102
rect 343338 363978 343958 364046
rect 343338 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 343958 363978
rect 343338 346350 343958 363922
rect 343338 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 343958 346350
rect 343338 346226 343958 346294
rect 343338 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 343958 346226
rect 343338 346102 343958 346170
rect 343338 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 343958 346102
rect 343338 345978 343958 346046
rect 343338 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 343958 345978
rect 343338 328350 343958 345922
rect 344428 366418 344484 366428
rect 344428 343588 344484 366362
rect 345324 363300 345380 363310
rect 344428 343522 344484 343532
rect 345212 353444 345268 353454
rect 343338 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 343958 328350
rect 343338 328226 343958 328294
rect 343338 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 343958 328226
rect 343338 328102 343958 328170
rect 343338 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 343958 328102
rect 343338 327978 343958 328046
rect 343338 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 343958 327978
rect 343338 310350 343958 327922
rect 343338 310294 343434 310350
rect 343490 310294 343558 310350
rect 343614 310294 343682 310350
rect 343738 310294 343806 310350
rect 343862 310294 343958 310350
rect 343338 310226 343958 310294
rect 343338 310170 343434 310226
rect 343490 310170 343558 310226
rect 343614 310170 343682 310226
rect 343738 310170 343806 310226
rect 343862 310170 343958 310226
rect 343338 310102 343958 310170
rect 343338 310046 343434 310102
rect 343490 310046 343558 310102
rect 343614 310046 343682 310102
rect 343738 310046 343806 310102
rect 343862 310046 343958 310102
rect 343338 309978 343958 310046
rect 343338 309922 343434 309978
rect 343490 309922 343558 309978
rect 343614 309922 343682 309978
rect 343738 309922 343806 309978
rect 343862 309922 343958 309978
rect 343338 292350 343958 309922
rect 343338 292294 343434 292350
rect 343490 292294 343558 292350
rect 343614 292294 343682 292350
rect 343738 292294 343806 292350
rect 343862 292294 343958 292350
rect 343338 292226 343958 292294
rect 343338 292170 343434 292226
rect 343490 292170 343558 292226
rect 343614 292170 343682 292226
rect 343738 292170 343806 292226
rect 343862 292170 343958 292226
rect 343338 292102 343958 292170
rect 343338 292046 343434 292102
rect 343490 292046 343558 292102
rect 343614 292046 343682 292102
rect 343738 292046 343806 292102
rect 343862 292046 343958 292102
rect 343338 291978 343958 292046
rect 343338 291922 343434 291978
rect 343490 291922 343558 291978
rect 343614 291922 343682 291978
rect 343738 291922 343806 291978
rect 343862 291922 343958 291978
rect 342860 289762 342916 289772
rect 342860 288932 342916 288942
rect 342748 288036 342804 288046
rect 342748 287398 342804 287980
rect 342748 287332 342804 287342
rect 342748 284788 342804 284798
rect 342748 284004 342804 284732
rect 342748 283938 342804 283948
rect 342748 279076 342804 279086
rect 342748 275604 342804 279020
rect 342860 278852 342916 288876
rect 342860 278786 342916 278796
rect 342748 275538 342804 275548
rect 343338 274350 343958 291922
rect 343338 274294 343434 274350
rect 343490 274294 343558 274350
rect 343614 274294 343682 274350
rect 343738 274294 343806 274350
rect 343862 274294 343958 274350
rect 343338 274226 343958 274294
rect 343338 274170 343434 274226
rect 343490 274170 343558 274226
rect 343614 274170 343682 274226
rect 343738 274170 343806 274226
rect 343862 274170 343958 274226
rect 343338 274102 343958 274170
rect 343338 274046 343434 274102
rect 343490 274046 343558 274102
rect 343614 274046 343682 274102
rect 343738 274046 343806 274102
rect 343862 274046 343958 274102
rect 343338 273978 343958 274046
rect 343338 273922 343434 273978
rect 343490 273922 343558 273978
rect 343614 273922 343682 273978
rect 343738 273922 343806 273978
rect 343862 273922 343958 273978
rect 342860 271012 342916 271022
rect 342412 248434 342468 248444
rect 342748 253988 342804 253998
rect 342188 247762 342244 247772
rect 342748 247078 342804 253932
rect 341964 237682 342020 237692
rect 342636 247022 342804 247078
rect 342636 231058 342692 247022
rect 342860 236098 342916 270956
rect 342860 236032 342916 236042
rect 342972 269220 343028 269230
rect 342972 234478 343028 269164
rect 343338 256350 343958 273922
rect 343338 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 343958 256350
rect 343338 256226 343958 256294
rect 343338 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 343958 256226
rect 343338 256102 343958 256170
rect 343338 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 343958 256102
rect 343338 255978 343958 256046
rect 343338 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 343958 255978
rect 343084 248612 343140 248622
rect 343084 241138 343140 248556
rect 343084 241072 343140 241082
rect 342972 234412 343028 234422
rect 343338 238350 343958 255922
rect 343338 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 343958 238350
rect 343338 238226 343958 238294
rect 343338 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 343958 238226
rect 343338 238102 343958 238170
rect 343338 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 343958 238102
rect 343338 237978 343958 238046
rect 343338 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 343958 237978
rect 342636 230992 342692 231002
rect 343338 220350 343958 237922
rect 343338 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 343958 220350
rect 343338 220226 343958 220294
rect 343338 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 343958 220226
rect 343338 220102 343958 220170
rect 343338 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 343958 220102
rect 343338 219978 343958 220046
rect 343338 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 343958 219978
rect 342972 211078 343028 211088
rect 342972 201572 343028 211022
rect 342972 201506 343028 201516
rect 343338 202350 343958 219922
rect 343338 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 343958 202350
rect 343338 202226 343958 202294
rect 343338 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 343958 202226
rect 343338 202102 343958 202170
rect 343338 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 343958 202102
rect 343338 201978 343958 202046
rect 343338 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 343958 201978
rect 343338 193230 343958 201922
rect 344092 341796 344148 341806
rect 341852 192472 341908 192482
rect 344092 191638 344148 341740
rect 344316 340004 344372 340014
rect 344204 196196 344260 196206
rect 344204 195748 344260 196140
rect 344204 195682 344260 195692
rect 344316 192718 344372 339948
rect 344428 334628 344484 334638
rect 344428 252084 344484 334572
rect 344540 319396 344596 319406
rect 344540 272132 344596 319340
rect 344540 272066 344596 272076
rect 344652 275604 344708 275614
rect 344652 255388 344708 275548
rect 344652 255332 345044 255388
rect 344428 252018 344484 252028
rect 344316 192652 344372 192662
rect 344876 240324 344932 240334
rect 344876 191818 344932 240268
rect 344988 239764 345044 255332
rect 344988 197540 345044 239708
rect 344988 197474 345044 197484
rect 345100 253018 345156 253028
rect 345100 194964 345156 252962
rect 345100 194898 345156 194908
rect 344876 191752 344932 191762
rect 344092 191572 344148 191582
rect 319752 190350 320072 190384
rect 319752 190294 319822 190350
rect 319878 190294 319946 190350
rect 320002 190294 320072 190350
rect 319752 190226 320072 190294
rect 319752 190170 319822 190226
rect 319878 190170 319946 190226
rect 320002 190170 320072 190226
rect 319752 190102 320072 190170
rect 319752 190046 319822 190102
rect 319878 190046 319946 190102
rect 320002 190046 320072 190102
rect 319752 189978 320072 190046
rect 319752 189922 319822 189978
rect 319878 189922 319946 189978
rect 320002 189922 320072 189978
rect 319752 189888 320072 189922
rect 328320 190350 328640 190384
rect 328320 190294 328390 190350
rect 328446 190294 328514 190350
rect 328570 190294 328640 190350
rect 328320 190226 328640 190294
rect 328320 190170 328390 190226
rect 328446 190170 328514 190226
rect 328570 190170 328640 190226
rect 328320 190102 328640 190170
rect 328320 190046 328390 190102
rect 328446 190046 328514 190102
rect 328570 190046 328640 190102
rect 328320 189978 328640 190046
rect 328320 189922 328390 189978
rect 328446 189922 328514 189978
rect 328570 189922 328640 189978
rect 328320 189888 328640 189922
rect 336888 190350 337208 190384
rect 336888 190294 336958 190350
rect 337014 190294 337082 190350
rect 337138 190294 337208 190350
rect 336888 190226 337208 190294
rect 336888 190170 336958 190226
rect 337014 190170 337082 190226
rect 337138 190170 337208 190226
rect 336888 190102 337208 190170
rect 336888 190046 336958 190102
rect 337014 190046 337082 190102
rect 337138 190046 337208 190102
rect 336888 189978 337208 190046
rect 336888 189922 336958 189978
rect 337014 189922 337082 189978
rect 337138 189922 337208 189978
rect 336888 189888 337208 189922
rect 324036 184350 324356 184384
rect 324036 184294 324106 184350
rect 324162 184294 324230 184350
rect 324286 184294 324356 184350
rect 324036 184226 324356 184294
rect 324036 184170 324106 184226
rect 324162 184170 324230 184226
rect 324286 184170 324356 184226
rect 324036 184102 324356 184170
rect 324036 184046 324106 184102
rect 324162 184046 324230 184102
rect 324286 184046 324356 184102
rect 324036 183978 324356 184046
rect 324036 183922 324106 183978
rect 324162 183922 324230 183978
rect 324286 183922 324356 183978
rect 324036 183888 324356 183922
rect 332604 184350 332924 184384
rect 332604 184294 332674 184350
rect 332730 184294 332798 184350
rect 332854 184294 332924 184350
rect 332604 184226 332924 184294
rect 332604 184170 332674 184226
rect 332730 184170 332798 184226
rect 332854 184170 332924 184226
rect 332604 184102 332924 184170
rect 332604 184046 332674 184102
rect 332730 184046 332798 184102
rect 332854 184046 332924 184102
rect 332604 183978 332924 184046
rect 332604 183922 332674 183978
rect 332730 183922 332798 183978
rect 332854 183922 332924 183978
rect 332604 183888 332924 183922
rect 341172 184350 341492 184384
rect 341172 184294 341242 184350
rect 341298 184294 341366 184350
rect 341422 184294 341492 184350
rect 341172 184226 341492 184294
rect 341172 184170 341242 184226
rect 341298 184170 341366 184226
rect 341422 184170 341492 184226
rect 341172 184102 341492 184170
rect 341172 184046 341242 184102
rect 341298 184046 341366 184102
rect 341422 184046 341492 184102
rect 341172 183978 341492 184046
rect 341172 183922 341242 183978
rect 341298 183922 341366 183978
rect 341422 183922 341492 183978
rect 341172 183888 341492 183922
rect 345212 173998 345268 353388
rect 345324 192358 345380 363244
rect 345436 360612 345492 360622
rect 345436 195778 345492 360556
rect 345548 241444 345604 396602
rect 347058 388350 347678 405922
rect 357644 404578 357700 407582
rect 357084 404522 357700 404578
rect 357756 408212 358148 408268
rect 357756 406918 357812 408212
rect 347058 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 347678 388350
rect 347058 388226 347678 388294
rect 347058 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 347678 388226
rect 347058 388102 347678 388170
rect 347058 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 347678 388102
rect 347058 387978 347678 388046
rect 347058 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 347678 387978
rect 346108 380100 346164 380110
rect 345884 347172 345940 347182
rect 345548 241378 345604 241388
rect 345660 298788 345716 298798
rect 345660 196756 345716 298732
rect 345660 196690 345716 196700
rect 345772 238644 345828 238654
rect 345548 196644 345604 196654
rect 345548 195972 345604 196588
rect 345548 195906 345604 195916
rect 345436 195712 345492 195722
rect 345772 194852 345828 238588
rect 345772 194786 345828 194796
rect 345324 192292 345380 192302
rect 345456 190350 345776 190384
rect 345456 190294 345526 190350
rect 345582 190294 345650 190350
rect 345706 190294 345776 190350
rect 345456 190226 345776 190294
rect 345456 190170 345526 190226
rect 345582 190170 345650 190226
rect 345706 190170 345776 190226
rect 345456 190102 345776 190170
rect 345456 190046 345526 190102
rect 345582 190046 345650 190102
rect 345706 190046 345776 190102
rect 345456 189978 345776 190046
rect 345456 189922 345526 189978
rect 345582 189922 345650 189978
rect 345706 189922 345776 189978
rect 345456 189888 345776 189922
rect 345884 175258 345940 347116
rect 345996 198212 346052 198222
rect 345996 196678 346052 198156
rect 345996 196612 346052 196622
rect 345884 175192 345940 175202
rect 345212 173932 345268 173942
rect 319752 172350 320072 172384
rect 319752 172294 319822 172350
rect 319878 172294 319946 172350
rect 320002 172294 320072 172350
rect 319752 172226 320072 172294
rect 319752 172170 319822 172226
rect 319878 172170 319946 172226
rect 320002 172170 320072 172226
rect 319752 172102 320072 172170
rect 319752 172046 319822 172102
rect 319878 172046 319946 172102
rect 320002 172046 320072 172102
rect 319752 171978 320072 172046
rect 319752 171922 319822 171978
rect 319878 171922 319946 171978
rect 320002 171922 320072 171978
rect 319752 171888 320072 171922
rect 328320 172350 328640 172384
rect 328320 172294 328390 172350
rect 328446 172294 328514 172350
rect 328570 172294 328640 172350
rect 328320 172226 328640 172294
rect 328320 172170 328390 172226
rect 328446 172170 328514 172226
rect 328570 172170 328640 172226
rect 328320 172102 328640 172170
rect 328320 172046 328390 172102
rect 328446 172046 328514 172102
rect 328570 172046 328640 172102
rect 328320 171978 328640 172046
rect 328320 171922 328390 171978
rect 328446 171922 328514 171978
rect 328570 171922 328640 171978
rect 328320 171888 328640 171922
rect 336888 172350 337208 172384
rect 336888 172294 336958 172350
rect 337014 172294 337082 172350
rect 337138 172294 337208 172350
rect 336888 172226 337208 172294
rect 336888 172170 336958 172226
rect 337014 172170 337082 172226
rect 337138 172170 337208 172226
rect 336888 172102 337208 172170
rect 336888 172046 336958 172102
rect 337014 172046 337082 172102
rect 337138 172046 337208 172102
rect 336888 171978 337208 172046
rect 336888 171922 336958 171978
rect 337014 171922 337082 171978
rect 337138 171922 337208 171978
rect 336888 171888 337208 171922
rect 345456 172350 345776 172384
rect 345456 172294 345526 172350
rect 345582 172294 345650 172350
rect 345706 172294 345776 172350
rect 345456 172226 345776 172294
rect 345456 172170 345526 172226
rect 345582 172170 345650 172226
rect 345706 172170 345776 172226
rect 345456 172102 345776 172170
rect 345456 172046 345526 172102
rect 345582 172046 345650 172102
rect 345706 172046 345776 172102
rect 345456 171978 345776 172046
rect 345456 171922 345526 171978
rect 345582 171922 345650 171978
rect 345706 171922 345776 171978
rect 345456 171888 345776 171922
rect 324036 166350 324356 166384
rect 324036 166294 324106 166350
rect 324162 166294 324230 166350
rect 324286 166294 324356 166350
rect 324036 166226 324356 166294
rect 324036 166170 324106 166226
rect 324162 166170 324230 166226
rect 324286 166170 324356 166226
rect 324036 166102 324356 166170
rect 324036 166046 324106 166102
rect 324162 166046 324230 166102
rect 324286 166046 324356 166102
rect 324036 165978 324356 166046
rect 324036 165922 324106 165978
rect 324162 165922 324230 165978
rect 324286 165922 324356 165978
rect 324036 165888 324356 165922
rect 332604 166350 332924 166384
rect 332604 166294 332674 166350
rect 332730 166294 332798 166350
rect 332854 166294 332924 166350
rect 332604 166226 332924 166294
rect 332604 166170 332674 166226
rect 332730 166170 332798 166226
rect 332854 166170 332924 166226
rect 332604 166102 332924 166170
rect 332604 166046 332674 166102
rect 332730 166046 332798 166102
rect 332854 166046 332924 166102
rect 332604 165978 332924 166046
rect 332604 165922 332674 165978
rect 332730 165922 332798 165978
rect 332854 165922 332924 165978
rect 332604 165888 332924 165922
rect 341172 166350 341492 166384
rect 341172 166294 341242 166350
rect 341298 166294 341366 166350
rect 341422 166294 341492 166350
rect 341172 166226 341492 166294
rect 341172 166170 341242 166226
rect 341298 166170 341366 166226
rect 341422 166170 341492 166226
rect 341172 166102 341492 166170
rect 341172 166046 341242 166102
rect 341298 166046 341366 166102
rect 341422 166046 341492 166102
rect 341172 165978 341492 166046
rect 341172 165922 341242 165978
rect 341298 165922 341366 165978
rect 341422 165922 341492 165978
rect 341172 165888 341492 165922
rect 317436 160066 317492 160076
rect 324380 157892 324436 157902
rect 324380 157798 324436 157836
rect 324380 157732 324436 157742
rect 330652 157892 330708 157902
rect 317324 157714 317380 157724
rect 330652 157618 330708 157836
rect 330652 157552 330708 157562
rect 332220 157892 332276 157902
rect 317100 157490 317156 157500
rect 332220 157438 332276 157836
rect 332220 157372 332276 157382
rect 316338 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 316958 154350
rect 316338 154226 316958 154294
rect 316338 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 316958 154226
rect 316338 154102 316958 154170
rect 316338 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 316958 154102
rect 316338 153978 316958 154046
rect 316338 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 316958 153978
rect 316338 136350 316958 153922
rect 343338 148350 343958 163170
rect 346108 157618 346164 380044
rect 347058 370350 347678 387922
rect 348908 401716 348964 401726
rect 347058 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 347678 370350
rect 347058 370226 347678 370294
rect 347058 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 347678 370226
rect 347058 370102 347678 370170
rect 347058 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 347678 370102
rect 347058 369978 347678 370046
rect 347058 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 347678 369978
rect 347058 352350 347678 369922
rect 347058 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 347678 352350
rect 347058 352226 347678 352294
rect 347058 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 347678 352226
rect 347058 352102 347678 352170
rect 347058 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 347678 352102
rect 347058 351978 347678 352046
rect 347058 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 347678 351978
rect 347058 334350 347678 351922
rect 347058 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 347678 334350
rect 347058 334226 347678 334294
rect 347058 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 347678 334226
rect 347058 334102 347678 334170
rect 347058 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 347678 334102
rect 347058 333978 347678 334046
rect 347058 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 347678 333978
rect 346780 330148 346836 330158
rect 346668 329252 346724 329262
rect 346220 315812 346276 315822
rect 346220 284788 346276 315756
rect 346332 310436 346388 310446
rect 346332 296548 346388 310380
rect 346332 296482 346388 296492
rect 346220 284722 346276 284732
rect 346220 284116 346276 284126
rect 346220 243118 346276 284060
rect 346220 243052 346276 243062
rect 346556 214564 346612 214574
rect 346444 194964 346500 194974
rect 346332 193258 346388 193268
rect 346108 157552 346164 157562
rect 346220 191638 346276 191648
rect 346220 159796 346276 191582
rect 346332 184828 346388 193202
rect 346444 192500 346500 194908
rect 346444 192434 346500 192444
rect 346332 184772 346500 184828
rect 346444 163940 346500 184772
rect 346556 175476 346612 214508
rect 346556 175410 346612 175420
rect 346668 167076 346724 329196
rect 346668 167010 346724 167020
rect 346444 163874 346500 163884
rect 346780 163828 346836 330092
rect 347058 316350 347678 333922
rect 347058 316294 347154 316350
rect 347210 316294 347278 316350
rect 347334 316294 347402 316350
rect 347458 316294 347526 316350
rect 347582 316294 347678 316350
rect 347058 316226 347678 316294
rect 347058 316170 347154 316226
rect 347210 316170 347278 316226
rect 347334 316170 347402 316226
rect 347458 316170 347526 316226
rect 347582 316170 347678 316226
rect 347058 316102 347678 316170
rect 347058 316046 347154 316102
rect 347210 316046 347278 316102
rect 347334 316046 347402 316102
rect 347458 316046 347526 316102
rect 347582 316046 347678 316102
rect 347058 315978 347678 316046
rect 347058 315922 347154 315978
rect 347210 315922 347278 315978
rect 347334 315922 347402 315978
rect 347458 315922 347526 315978
rect 347582 315922 347678 315978
rect 347058 298350 347678 315922
rect 347058 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 347678 298350
rect 347058 298226 347678 298294
rect 347058 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 347678 298226
rect 347058 298102 347678 298170
rect 347058 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 347678 298102
rect 347058 297978 347678 298046
rect 347058 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 347678 297978
rect 346780 163762 346836 163772
rect 346892 296996 346948 297006
rect 346220 157108 346276 159740
rect 346220 157042 346276 157052
rect 343338 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 343958 148350
rect 343338 148226 343958 148294
rect 343338 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 343958 148226
rect 343338 148102 343958 148170
rect 343338 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 343958 148102
rect 343338 147978 343958 148046
rect 343338 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 343958 147978
rect 316338 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 316958 136350
rect 316338 136226 316958 136294
rect 316338 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 316958 136226
rect 316338 136102 316958 136170
rect 316338 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 316958 136102
rect 316338 135978 316958 136046
rect 316338 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 316958 135978
rect 316338 118350 316958 135922
rect 316338 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 316958 118350
rect 316338 118226 316958 118294
rect 316338 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 316958 118226
rect 316338 118102 316958 118170
rect 316338 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 316958 118102
rect 316338 117978 316958 118046
rect 316338 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 316958 117978
rect 316338 100350 316958 117922
rect 316338 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 316958 100350
rect 316338 100226 316958 100294
rect 316338 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 316958 100226
rect 316338 100102 316958 100170
rect 316338 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 316958 100102
rect 316338 99978 316958 100046
rect 316338 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 316958 99978
rect 316338 84316 316958 99922
rect 330092 146998 330148 147008
rect 330092 84756 330148 146942
rect 330092 84690 330148 84700
rect 343338 130350 343958 147922
rect 343338 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 343958 130350
rect 343338 130226 343958 130294
rect 343338 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 343958 130226
rect 343338 130102 343958 130170
rect 343338 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 343958 130102
rect 343338 129978 343958 130046
rect 343338 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 343958 129978
rect 343338 112350 343958 129922
rect 346892 121940 346948 296940
rect 347058 280350 347678 297922
rect 347058 280294 347154 280350
rect 347210 280294 347278 280350
rect 347334 280294 347402 280350
rect 347458 280294 347526 280350
rect 347582 280294 347678 280350
rect 347058 280226 347678 280294
rect 347058 280170 347154 280226
rect 347210 280170 347278 280226
rect 347334 280170 347402 280226
rect 347458 280170 347526 280226
rect 347582 280170 347678 280226
rect 347058 280102 347678 280170
rect 347058 280046 347154 280102
rect 347210 280046 347278 280102
rect 347334 280046 347402 280102
rect 347458 280046 347526 280102
rect 347582 280046 347678 280102
rect 347058 279978 347678 280046
rect 347058 279922 347154 279978
rect 347210 279922 347278 279978
rect 347334 279922 347402 279978
rect 347458 279922 347526 279978
rect 347582 279922 347678 279978
rect 347058 262350 347678 279922
rect 347058 262294 347154 262350
rect 347210 262294 347278 262350
rect 347334 262294 347402 262350
rect 347458 262294 347526 262350
rect 347582 262294 347678 262350
rect 347058 262226 347678 262294
rect 347058 262170 347154 262226
rect 347210 262170 347278 262226
rect 347334 262170 347402 262226
rect 347458 262170 347526 262226
rect 347582 262170 347678 262226
rect 347058 262102 347678 262170
rect 347058 262046 347154 262102
rect 347210 262046 347278 262102
rect 347334 262046 347402 262102
rect 347458 262046 347526 262102
rect 347582 262046 347678 262102
rect 347058 261978 347678 262046
rect 347058 261922 347154 261978
rect 347210 261922 347278 261978
rect 347334 261922 347402 261978
rect 347458 261922 347526 261978
rect 347582 261922 347678 261978
rect 347058 244350 347678 261922
rect 347058 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 347678 244350
rect 347058 244226 347678 244294
rect 347058 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 347678 244226
rect 347058 244102 347678 244170
rect 347058 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 347678 244102
rect 347058 243978 347678 244046
rect 347058 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 347678 243978
rect 347058 226350 347678 243922
rect 347058 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 347678 226350
rect 347058 226226 347678 226294
rect 347058 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 347678 226226
rect 347058 226102 347678 226170
rect 347058 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 347678 226102
rect 347058 225978 347678 226046
rect 347058 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 347678 225978
rect 347058 208350 347678 225922
rect 347058 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 347678 208350
rect 347058 208226 347678 208294
rect 347058 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 347678 208226
rect 347058 208102 347678 208170
rect 347058 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 347678 208102
rect 347058 207978 347678 208046
rect 347058 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 347678 207978
rect 347058 193230 347678 207922
rect 347788 379988 347844 379998
rect 347004 191818 347060 191828
rect 347004 173818 347060 191762
rect 347004 173752 347060 173762
rect 346892 121874 346948 121884
rect 347058 154350 347678 163170
rect 347788 157438 347844 379932
rect 348572 375418 348628 375428
rect 348572 343140 348628 375362
rect 348572 343074 348628 343084
rect 348572 331044 348628 331054
rect 347900 324772 347956 324782
rect 347900 248612 347956 324716
rect 348012 321188 348068 321198
rect 348012 283892 348068 321132
rect 348012 283826 348068 283836
rect 348124 320292 348180 320302
rect 348124 283780 348180 320236
rect 348124 283714 348180 283724
rect 348236 283556 348292 283566
rect 348236 255388 348292 283500
rect 348236 255332 348516 255388
rect 347900 248546 347956 248556
rect 347788 157372 347844 157382
rect 348460 242038 348516 255332
rect 347058 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 347678 154350
rect 347058 154226 347678 154294
rect 347058 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 347678 154226
rect 347058 154102 347678 154170
rect 347058 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 347678 154102
rect 347058 153978 347678 154046
rect 347058 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 347678 153978
rect 347058 136350 347678 153922
rect 347058 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 347678 136350
rect 347058 136226 347678 136294
rect 347058 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 347678 136226
rect 347058 136102 347678 136170
rect 347058 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 347678 136102
rect 347058 135978 347678 136046
rect 347058 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 347678 135978
rect 343338 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 343958 112350
rect 343338 112226 343958 112294
rect 343338 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 343958 112226
rect 343338 112102 343958 112170
rect 343338 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 343958 112102
rect 343338 111978 343958 112046
rect 343338 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 343958 111978
rect 343338 94350 343958 111922
rect 343338 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 343958 94350
rect 343338 94226 343958 94294
rect 343338 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 343958 94226
rect 343338 94102 343958 94170
rect 343338 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 343958 94102
rect 343338 93978 343958 94046
rect 343338 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 343958 93978
rect 316132 82147 316452 82204
rect 316132 82091 316160 82147
rect 316216 82091 316264 82147
rect 316320 82091 316368 82147
rect 316424 82091 316452 82147
rect 316132 82043 316452 82091
rect 316132 81987 316160 82043
rect 316216 81987 316264 82043
rect 316320 81987 316368 82043
rect 316424 81987 316452 82043
rect 316132 81939 316452 81987
rect 316132 81883 316160 81939
rect 316216 81883 316264 81939
rect 316320 81883 316368 81939
rect 316424 81883 316452 81939
rect 316132 81826 316452 81883
rect 324448 82147 324768 82204
rect 324448 82091 324476 82147
rect 324532 82091 324580 82147
rect 324636 82091 324684 82147
rect 324740 82091 324768 82147
rect 324448 82043 324768 82091
rect 324448 81987 324476 82043
rect 324532 81987 324580 82043
rect 324636 81987 324684 82043
rect 324740 81987 324768 82043
rect 324448 81939 324768 81987
rect 324448 81883 324476 81939
rect 324532 81883 324580 81939
rect 324636 81883 324684 81939
rect 324740 81883 324768 81939
rect 324448 81826 324768 81883
rect 320290 76350 320610 76384
rect 320290 76294 320360 76350
rect 320416 76294 320484 76350
rect 320540 76294 320610 76350
rect 320290 76226 320610 76294
rect 320290 76170 320360 76226
rect 320416 76170 320484 76226
rect 320540 76170 320610 76226
rect 320290 76102 320610 76170
rect 320290 76046 320360 76102
rect 320416 76046 320484 76102
rect 320540 76046 320610 76102
rect 320290 75978 320610 76046
rect 320290 75922 320360 75978
rect 320416 75922 320484 75978
rect 320540 75922 320610 75978
rect 320290 75888 320610 75922
rect 343338 76350 343958 93922
rect 343338 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 343958 76350
rect 343338 76226 343958 76294
rect 343338 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 343958 76226
rect 343338 76102 343958 76170
rect 343338 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 343958 76102
rect 343338 75978 343958 76046
rect 343338 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 343958 75978
rect 316132 64350 316452 64384
rect 316132 64294 316202 64350
rect 316258 64294 316326 64350
rect 316382 64294 316452 64350
rect 316132 64226 316452 64294
rect 316132 64170 316202 64226
rect 316258 64170 316326 64226
rect 316382 64170 316452 64226
rect 316132 64102 316452 64170
rect 316132 64046 316202 64102
rect 316258 64046 316326 64102
rect 316382 64046 316452 64102
rect 316132 63978 316452 64046
rect 316132 63922 316202 63978
rect 316258 63922 316326 63978
rect 316382 63922 316452 63978
rect 316132 63888 316452 63922
rect 324448 64350 324768 64384
rect 324448 64294 324518 64350
rect 324574 64294 324642 64350
rect 324698 64294 324768 64350
rect 324448 64226 324768 64294
rect 324448 64170 324518 64226
rect 324574 64170 324642 64226
rect 324698 64170 324768 64226
rect 324448 64102 324768 64170
rect 324448 64046 324518 64102
rect 324574 64046 324642 64102
rect 324698 64046 324768 64102
rect 324448 63978 324768 64046
rect 324448 63922 324518 63978
rect 324574 63922 324642 63978
rect 324698 63922 324768 63978
rect 324448 63888 324768 63922
rect 320290 58350 320610 58384
rect 320290 58294 320360 58350
rect 320416 58294 320484 58350
rect 320540 58294 320610 58350
rect 320290 58226 320610 58294
rect 320290 58170 320360 58226
rect 320416 58170 320484 58226
rect 320540 58170 320610 58226
rect 320290 58102 320610 58170
rect 320290 58046 320360 58102
rect 320416 58046 320484 58102
rect 320540 58046 320610 58102
rect 320290 57978 320610 58046
rect 320290 57922 320360 57978
rect 320416 57922 320484 57978
rect 320540 57922 320610 57978
rect 320290 57888 320610 57922
rect 343338 58350 343958 75922
rect 343338 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 343958 58350
rect 343338 58226 343958 58294
rect 343338 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 343958 58226
rect 343338 58102 343958 58170
rect 343338 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 343958 58102
rect 343338 57978 343958 58046
rect 343338 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 343958 57978
rect 315308 50306 315364 50316
rect 315084 48514 315140 48524
rect 314972 4912 315028 4922
rect 316338 46350 316958 50964
rect 316338 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 316958 46350
rect 316338 46226 316958 46294
rect 316338 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 316958 46226
rect 316338 46102 316958 46170
rect 316338 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 316958 46102
rect 316338 45978 316958 46046
rect 316338 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 316958 45978
rect 316338 28350 316958 45922
rect 316338 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 316958 28350
rect 316338 28226 316958 28294
rect 316338 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 316958 28226
rect 316338 28102 316958 28170
rect 316338 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 316958 28102
rect 316338 27978 316958 28046
rect 316338 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 316958 27978
rect 316338 10350 316958 27922
rect 316338 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 316958 10350
rect 316338 10226 316958 10294
rect 316338 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 316958 10226
rect 316338 10102 316958 10170
rect 316338 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 316958 10102
rect 316338 9978 316958 10046
rect 316338 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 316958 9978
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 312618 4102 313238 4170
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 316338 -1120 316958 9922
rect 316338 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 316958 -1120
rect 316338 -1244 316958 -1176
rect 316338 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 316958 -1244
rect 316338 -1368 316958 -1300
rect 316338 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 316958 -1368
rect 316338 -1492 316958 -1424
rect 316338 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 316958 -1492
rect 316338 -1644 316958 -1548
rect 343338 40350 343958 57922
rect 343338 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 343958 40350
rect 343338 40226 343958 40294
rect 343338 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 343958 40226
rect 343338 40102 343958 40170
rect 343338 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 343958 40102
rect 343338 39978 343958 40046
rect 343338 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 343958 39978
rect 343338 22350 343958 39922
rect 343338 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 343958 22350
rect 343338 22226 343958 22294
rect 343338 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 343958 22226
rect 343338 22102 343958 22170
rect 343338 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 343958 22102
rect 343338 21978 343958 22046
rect 343338 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 343958 21978
rect 343338 4350 343958 21922
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 343338 4102 343958 4170
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 347058 118350 347678 135922
rect 348460 128548 348516 241982
rect 348572 152628 348628 330988
rect 348572 152562 348628 152572
rect 348684 326564 348740 326574
rect 348684 150500 348740 326508
rect 348684 150434 348740 150444
rect 348796 323876 348852 323886
rect 348796 148820 348852 323820
rect 348908 237538 348964 401660
rect 349020 397198 349076 397208
rect 349020 240058 349076 397142
rect 353500 397018 353556 397028
rect 349468 383124 349524 383134
rect 349020 239992 349076 240002
rect 349132 248500 349188 248510
rect 348908 237472 348964 237482
rect 348796 148754 348852 148764
rect 348460 128482 348516 128492
rect 349132 121828 349188 248444
rect 349356 242004 349412 242014
rect 349132 121762 349188 121772
rect 349244 238644 349300 238654
rect 347058 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 347678 118350
rect 347058 118226 347678 118294
rect 347058 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 347678 118226
rect 347058 118102 347678 118170
rect 347058 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 347678 118102
rect 347058 117978 347678 118046
rect 347058 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 347678 117978
rect 347058 100350 347678 117922
rect 347058 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 347678 100350
rect 347058 100226 347678 100294
rect 347058 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 347678 100226
rect 347058 100102 347678 100170
rect 347058 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 347678 100102
rect 347058 99978 347678 100046
rect 347058 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 347678 99978
rect 347058 82350 347678 99922
rect 347058 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 347678 82350
rect 347058 82226 347678 82294
rect 347058 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 347678 82226
rect 347058 82102 347678 82170
rect 347058 82046 347154 82102
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 347678 82102
rect 347058 81978 347678 82046
rect 347058 81922 347154 81978
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 347678 81978
rect 347058 64350 347678 81922
rect 347058 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 347678 64350
rect 347058 64226 347678 64294
rect 347058 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 347678 64226
rect 347058 64102 347678 64170
rect 347058 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 347678 64102
rect 347058 63978 347678 64046
rect 347058 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 347678 63978
rect 347058 46350 347678 63922
rect 349244 48020 349300 238588
rect 349244 47954 349300 47964
rect 347058 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 347678 46350
rect 347058 46226 347678 46294
rect 347058 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 347678 46226
rect 347058 46102 347678 46170
rect 347058 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 347678 46102
rect 347058 45978 347678 46046
rect 347058 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 347678 45978
rect 347058 28350 347678 45922
rect 349356 45332 349412 241948
rect 349468 157798 349524 383068
rect 350252 379738 350308 379748
rect 349580 314020 349636 314030
rect 349580 193284 349636 313964
rect 349692 306852 349748 306862
rect 349692 209972 349748 306796
rect 349692 209906 349748 209916
rect 349804 209412 349860 209422
rect 349804 196588 349860 209356
rect 349580 193218 349636 193228
rect 349692 196532 349860 196588
rect 349692 165060 349748 196532
rect 349692 164994 349748 165004
rect 349468 157732 349524 157742
rect 350252 84980 350308 379682
rect 350588 372178 350644 372188
rect 350364 332836 350420 332846
rect 350364 162260 350420 332780
rect 350476 327460 350532 327470
rect 350476 167300 350532 327404
rect 350588 302260 350644 372122
rect 352268 331940 352324 331950
rect 350588 302194 350644 302204
rect 350700 322980 350756 322990
rect 350476 167234 350532 167244
rect 350588 240660 350644 240670
rect 350364 162194 350420 162204
rect 350588 126868 350644 240604
rect 350700 178052 350756 322924
rect 351932 312228 351988 312238
rect 351148 308644 351204 308654
rect 350812 302260 350868 302270
rect 350812 205940 350868 302204
rect 350812 205874 350868 205884
rect 350700 177986 350756 177996
rect 350812 196678 350868 196688
rect 350812 170578 350868 196622
rect 351036 194628 351092 194638
rect 351036 191828 351092 194572
rect 351036 191762 351092 191772
rect 351148 191716 351204 308588
rect 351148 191650 351204 191660
rect 351260 295204 351316 295214
rect 351260 191604 351316 295148
rect 351372 256676 351428 256686
rect 351372 225988 351428 256620
rect 351372 225922 351428 225932
rect 351260 191538 351316 191548
rect 351372 192718 351428 192728
rect 350812 170512 350868 170522
rect 351372 159572 351428 192662
rect 351372 159506 351428 159516
rect 350588 126802 350644 126812
rect 350252 84914 350308 84924
rect 351932 50148 351988 312172
rect 352156 301476 352212 301486
rect 352044 290836 352100 290846
rect 352044 120148 352100 290780
rect 352156 133476 352212 301420
rect 352268 165620 352324 331884
rect 352380 325668 352436 325678
rect 352380 168980 352436 325612
rect 352828 313124 352884 313134
rect 352380 168914 352436 168924
rect 352492 305956 352548 305966
rect 352268 165554 352324 165564
rect 352492 162484 352548 305900
rect 352828 282212 352884 313068
rect 352828 282146 352884 282156
rect 353500 240238 353556 396962
rect 355852 396838 355908 396848
rect 354396 394858 354452 394868
rect 354284 376292 354340 376302
rect 354284 368758 354340 376236
rect 354284 368692 354340 368702
rect 354060 335524 354116 335534
rect 353948 328356 354004 328366
rect 353500 240172 353556 240182
rect 353612 322084 353668 322094
rect 352492 162418 352548 162428
rect 352604 196644 352660 196654
rect 352156 133410 352212 133420
rect 352604 124740 352660 196588
rect 352716 192538 352772 192548
rect 352716 175140 352772 192482
rect 352716 175074 352772 175084
rect 352940 151172 352996 151182
rect 352940 150598 352996 151116
rect 352940 150532 352996 150542
rect 352604 124674 352660 124684
rect 352044 120082 352100 120092
rect 351932 50082 351988 50092
rect 349356 45266 349412 45276
rect 353612 45220 353668 322028
rect 353724 316708 353780 316718
rect 353724 50036 353780 316652
rect 353836 280756 353892 280766
rect 353836 51492 353892 280700
rect 353948 152740 354004 328300
rect 354060 168868 354116 335468
rect 354284 304164 354340 304174
rect 354060 168802 354116 168812
rect 354172 302372 354228 302382
rect 353948 152674 354004 152684
rect 354172 136388 354228 302316
rect 354284 142212 354340 304108
rect 354396 237718 354452 394802
rect 355404 366598 355460 366608
rect 355292 311332 355348 311342
rect 354620 307748 354676 307758
rect 354396 237652 354452 237662
rect 354508 285796 354564 285806
rect 354508 235198 354564 285740
rect 354620 280420 354676 307692
rect 354732 293188 354788 293198
rect 354732 280532 354788 293132
rect 354732 280466 354788 280476
rect 354620 280354 354676 280364
rect 354508 235132 354564 235142
rect 354396 214318 354452 214328
rect 354396 167972 354452 214262
rect 355180 210898 355236 210908
rect 355180 173572 355236 210842
rect 355180 173506 355236 173516
rect 354396 167906 354452 167916
rect 354284 142146 354340 142156
rect 354172 136322 354228 136332
rect 353836 51426 353892 51436
rect 353724 49970 353780 49980
rect 355292 48132 355348 311276
rect 355404 284900 355460 366542
rect 355628 333732 355684 333742
rect 355404 284834 355460 284844
rect 355516 289828 355572 289838
rect 355404 278964 355460 278974
rect 355404 52948 355460 278908
rect 355516 118468 355572 289772
rect 355628 164052 355684 333676
rect 355628 163986 355684 163996
rect 355740 300580 355796 300590
rect 355740 131908 355796 300524
rect 355852 242758 355908 396782
rect 357084 384748 357140 404522
rect 357196 404404 357252 404414
rect 357196 401698 357252 404348
rect 357196 401642 357476 401698
rect 356972 384692 357140 384748
rect 356524 356158 356580 356168
rect 356524 354788 356580 356102
rect 356524 354722 356580 354732
rect 356188 325918 356244 325928
rect 356188 325668 356244 325862
rect 356188 325602 356244 325612
rect 356524 299572 356580 299582
rect 356524 296758 356580 299516
rect 356524 296692 356580 296702
rect 355852 242692 355908 242702
rect 355964 284004 356020 284014
rect 355852 235198 355908 235208
rect 355852 169316 355908 235142
rect 355964 170772 356020 283948
rect 356748 273140 356804 273150
rect 356748 235172 356804 273084
rect 356860 273028 356916 273038
rect 356860 255388 356916 272972
rect 356972 257012 357028 384692
rect 357084 369118 357140 369128
rect 357084 348852 357140 369062
rect 357084 347844 357140 348796
rect 357084 347778 357140 347788
rect 357196 367108 357252 367118
rect 356972 256946 357028 256956
rect 356860 255332 357140 255388
rect 356972 249844 357028 249854
rect 356972 243628 357028 249788
rect 357084 249508 357140 255332
rect 357084 249442 357140 249452
rect 356972 243572 357140 243628
rect 356748 234500 356804 235116
rect 356748 234434 356804 234444
rect 356972 238196 357028 238206
rect 356860 220724 356916 220734
rect 355964 170706 356020 170716
rect 356076 197092 356132 197102
rect 355852 169250 355908 169260
rect 356076 139300 356132 197036
rect 356748 181412 356804 181422
rect 356188 154532 356244 154542
rect 356188 153478 356244 154476
rect 356188 153412 356244 153422
rect 356076 139234 356132 139244
rect 355740 131842 355796 131852
rect 356748 127652 356804 181356
rect 356860 179788 356916 220668
rect 356972 183876 357028 238140
rect 356972 183810 357028 183820
rect 356972 181188 357028 181198
rect 356972 181018 357028 181132
rect 356972 180952 357028 180962
rect 356860 179732 357028 179788
rect 356972 175812 357028 179732
rect 356972 175364 357028 175756
rect 356972 175298 357028 175308
rect 357084 164948 357140 243572
rect 356972 164612 357028 164622
rect 356972 163156 357028 164556
rect 356972 141988 357028 163100
rect 356972 141922 357028 141932
rect 357084 138628 357140 164892
rect 357196 154532 357252 367052
rect 357308 308998 357364 309008
rect 357308 308084 357364 308942
rect 357308 308018 357364 308028
rect 357420 273140 357476 401642
rect 357756 384748 357812 406862
rect 357420 273074 357476 273084
rect 357532 384692 357812 384748
rect 357420 268772 357476 268782
rect 357420 267428 357476 268716
rect 357196 154466 357252 154476
rect 357308 257012 357364 257022
rect 357308 255780 357364 256956
rect 357308 164836 357364 255724
rect 357084 138562 357140 138572
rect 357308 132020 357364 164780
rect 357420 147718 357476 267372
rect 357532 261380 357588 384692
rect 357868 383158 357924 383168
rect 357868 376292 357924 383102
rect 357868 376226 357924 376236
rect 357756 347844 357812 347854
rect 357532 164612 357588 261324
rect 357532 164546 357588 164556
rect 357644 343140 357700 343150
rect 357644 166404 357700 343084
rect 357420 146998 357476 147662
rect 357644 147028 357700 166348
rect 357756 163044 357812 347788
rect 357868 325668 357924 325678
rect 357868 230338 357924 325612
rect 357868 230272 357924 230282
rect 357980 307972 358036 307982
rect 357980 230244 358036 307916
rect 357980 230178 358036 230188
rect 358652 280644 358708 280654
rect 358540 192358 358596 192368
rect 358428 174692 358484 174702
rect 358428 173098 358484 174636
rect 358428 173032 358484 173042
rect 358540 171220 358596 192302
rect 358540 171154 358596 171164
rect 357756 153860 357812 162988
rect 357756 153794 357812 153804
rect 357644 146962 357700 146972
rect 357420 146932 357476 146942
rect 357308 131954 357364 131964
rect 356748 127586 356804 127596
rect 355516 118402 355572 118412
rect 355404 52882 355460 52892
rect 358652 52724 358708 280588
rect 358764 239540 358820 409922
rect 359548 408436 359604 408446
rect 358988 406918 359044 406928
rect 358988 390964 359044 406862
rect 358988 390898 359044 390908
rect 359548 389396 359604 408380
rect 359772 404964 359828 404974
rect 359548 389330 359604 389340
rect 359660 396676 359716 396686
rect 359436 331044 359492 331054
rect 358988 313348 359044 313358
rect 358764 239474 358820 239484
rect 358876 284116 358932 284126
rect 358764 230244 358820 230254
rect 358764 168778 358820 230188
rect 358764 168712 358820 168722
rect 358876 126980 358932 284060
rect 358988 240324 359044 313292
rect 359324 255892 359380 255902
rect 359324 255718 359380 255836
rect 359324 255652 359380 255662
rect 358988 240258 359044 240268
rect 359100 230338 359156 230348
rect 358988 197988 359044 197998
rect 358988 145124 359044 197932
rect 359100 170548 359156 230282
rect 359212 214138 359268 214148
rect 359212 176338 359268 214082
rect 359212 176272 359268 176282
rect 359324 197540 359380 197550
rect 359100 170482 359156 170492
rect 358988 145058 359044 145068
rect 358876 126914 358932 126924
rect 359324 120484 359380 197484
rect 359436 174020 359492 330988
rect 359436 173954 359492 173964
rect 359548 264628 359604 264638
rect 359324 120418 359380 120428
rect 359548 117012 359604 264572
rect 359660 241108 359716 396620
rect 359660 241042 359716 241052
rect 359772 240212 359828 404908
rect 359884 389956 359940 410060
rect 362012 407428 362068 407438
rect 360444 407098 360500 407108
rect 359996 403508 360052 403518
rect 359996 396478 360052 403452
rect 359996 396422 360276 396478
rect 359884 389890 359940 389900
rect 360220 389638 360276 396422
rect 360444 392644 360500 407042
rect 361900 400036 361956 400046
rect 360444 392578 360500 392588
rect 360556 399924 360612 399934
rect 359884 389582 360276 389638
rect 359884 389508 359940 389582
rect 359884 389442 359940 389452
rect 359884 388948 359940 388958
rect 360556 388918 360612 399868
rect 361900 396508 361956 399980
rect 361676 396452 361956 396508
rect 361676 391438 361732 396452
rect 362012 395758 362068 407372
rect 511308 404404 511364 590604
rect 514892 590212 514948 590222
rect 511308 404338 511364 404348
rect 511420 567028 511476 567038
rect 471996 398244 472052 398254
rect 361788 395702 362068 395758
rect 375452 397348 375508 397358
rect 361788 392420 361844 395702
rect 362124 395578 362180 395588
rect 362012 395522 362124 395578
rect 361788 392354 361844 392364
rect 361900 392644 361956 392654
rect 361900 391978 361956 392588
rect 361900 391912 361956 391922
rect 361676 391372 361732 391382
rect 359940 388892 360612 388918
rect 359884 388862 360612 388892
rect 362012 384748 362068 395522
rect 362124 395512 362180 395522
rect 375452 395578 375508 397292
rect 375452 395512 375508 395522
rect 362908 395108 362964 395118
rect 362908 392756 362964 395052
rect 362908 392690 362964 392700
rect 405468 394548 405524 394558
rect 405468 392532 405524 394492
rect 441756 394548 441812 394558
rect 438508 394212 438564 394222
rect 438508 393988 438564 394156
rect 438508 393922 438564 393932
rect 405468 392466 405524 392476
rect 441756 392338 441812 394492
rect 471996 392420 472052 398188
rect 511420 397348 511476 566972
rect 514892 409618 514948 590156
rect 527658 580350 528278 596784
rect 527658 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 528278 580350
rect 527658 580226 528278 580294
rect 527658 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 528278 580226
rect 527658 580102 528278 580170
rect 527658 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 528278 580102
rect 527658 579978 528278 580046
rect 527658 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 528278 579978
rect 527658 562350 528278 579922
rect 527658 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 528278 562350
rect 527658 562226 528278 562294
rect 527658 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 528278 562226
rect 527658 562102 528278 562170
rect 527658 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 528278 562102
rect 527658 561978 528278 562046
rect 527658 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 528278 561978
rect 517008 550350 517328 550384
rect 517008 550294 517078 550350
rect 517134 550294 517202 550350
rect 517258 550294 517328 550350
rect 517008 550226 517328 550294
rect 517008 550170 517078 550226
rect 517134 550170 517202 550226
rect 517258 550170 517328 550226
rect 517008 550102 517328 550170
rect 517008 550046 517078 550102
rect 517134 550046 517202 550102
rect 517258 550046 517328 550102
rect 517008 549978 517328 550046
rect 517008 549922 517078 549978
rect 517134 549922 517202 549978
rect 517258 549922 517328 549978
rect 517008 549888 517328 549922
rect 527658 544350 528278 561922
rect 527658 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 528278 544350
rect 527658 544226 528278 544294
rect 527658 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 528278 544226
rect 527658 544102 528278 544170
rect 527658 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 528278 544102
rect 527658 543978 528278 544046
rect 527658 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 528278 543978
rect 517008 532350 517328 532384
rect 517008 532294 517078 532350
rect 517134 532294 517202 532350
rect 517258 532294 517328 532350
rect 517008 532226 517328 532294
rect 517008 532170 517078 532226
rect 517134 532170 517202 532226
rect 517258 532170 517328 532226
rect 517008 532102 517328 532170
rect 517008 532046 517078 532102
rect 517134 532046 517202 532102
rect 517258 532046 517328 532102
rect 517008 531978 517328 532046
rect 517008 531922 517078 531978
rect 517134 531922 517202 531978
rect 517258 531922 517328 531978
rect 517008 531888 517328 531922
rect 527658 526350 528278 543922
rect 527658 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 528278 526350
rect 527658 526226 528278 526294
rect 527658 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 528278 526226
rect 527658 526102 528278 526170
rect 527658 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 528278 526102
rect 527658 525978 528278 526046
rect 527658 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 528278 525978
rect 517008 514350 517328 514384
rect 517008 514294 517078 514350
rect 517134 514294 517202 514350
rect 517258 514294 517328 514350
rect 517008 514226 517328 514294
rect 517008 514170 517078 514226
rect 517134 514170 517202 514226
rect 517258 514170 517328 514226
rect 517008 514102 517328 514170
rect 517008 514046 517078 514102
rect 517134 514046 517202 514102
rect 517258 514046 517328 514102
rect 517008 513978 517328 514046
rect 517008 513922 517078 513978
rect 517134 513922 517202 513978
rect 517258 513922 517328 513978
rect 517008 513888 517328 513922
rect 527658 508350 528278 525922
rect 527658 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 528278 508350
rect 527658 508226 528278 508294
rect 527658 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 528278 508226
rect 527658 508102 528278 508170
rect 527658 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 528278 508102
rect 527658 507978 528278 508046
rect 527658 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 528278 507978
rect 517008 496350 517328 496384
rect 517008 496294 517078 496350
rect 517134 496294 517202 496350
rect 517258 496294 517328 496350
rect 517008 496226 517328 496294
rect 517008 496170 517078 496226
rect 517134 496170 517202 496226
rect 517258 496170 517328 496226
rect 517008 496102 517328 496170
rect 517008 496046 517078 496102
rect 517134 496046 517202 496102
rect 517258 496046 517328 496102
rect 517008 495978 517328 496046
rect 517008 495922 517078 495978
rect 517134 495922 517202 495978
rect 517258 495922 517328 495978
rect 517008 495888 517328 495922
rect 527658 490350 528278 507922
rect 527658 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 528278 490350
rect 527658 490226 528278 490294
rect 527658 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 528278 490226
rect 527658 490102 528278 490170
rect 527658 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 528278 490102
rect 527658 489978 528278 490046
rect 527658 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 528278 489978
rect 517008 478350 517328 478384
rect 517008 478294 517078 478350
rect 517134 478294 517202 478350
rect 517258 478294 517328 478350
rect 517008 478226 517328 478294
rect 517008 478170 517078 478226
rect 517134 478170 517202 478226
rect 517258 478170 517328 478226
rect 517008 478102 517328 478170
rect 517008 478046 517078 478102
rect 517134 478046 517202 478102
rect 517258 478046 517328 478102
rect 517008 477978 517328 478046
rect 517008 477922 517078 477978
rect 517134 477922 517202 477978
rect 517258 477922 517328 477978
rect 517008 477888 517328 477922
rect 527658 472350 528278 489922
rect 527658 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 528278 472350
rect 527658 472226 528278 472294
rect 527658 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 528278 472226
rect 527658 472102 528278 472170
rect 527658 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 528278 472102
rect 527658 471978 528278 472046
rect 527658 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 528278 471978
rect 517008 460350 517328 460384
rect 517008 460294 517078 460350
rect 517134 460294 517202 460350
rect 517258 460294 517328 460350
rect 517008 460226 517328 460294
rect 517008 460170 517078 460226
rect 517134 460170 517202 460226
rect 517258 460170 517328 460226
rect 517008 460102 517328 460170
rect 517008 460046 517078 460102
rect 517134 460046 517202 460102
rect 517258 460046 517328 460102
rect 517008 459978 517328 460046
rect 517008 459922 517078 459978
rect 517134 459922 517202 459978
rect 517258 459922 517328 459978
rect 517008 459888 517328 459922
rect 527658 454350 528278 471922
rect 527658 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 528278 454350
rect 527658 454226 528278 454294
rect 527658 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 528278 454226
rect 527658 454102 528278 454170
rect 527658 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 528278 454102
rect 527658 453978 528278 454046
rect 527658 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 528278 453978
rect 517008 442350 517328 442384
rect 517008 442294 517078 442350
rect 517134 442294 517202 442350
rect 517258 442294 517328 442350
rect 517008 442226 517328 442294
rect 517008 442170 517078 442226
rect 517134 442170 517202 442226
rect 517258 442170 517328 442226
rect 517008 442102 517328 442170
rect 517008 442046 517078 442102
rect 517134 442046 517202 442102
rect 517258 442046 517328 442102
rect 517008 441978 517328 442046
rect 517008 441922 517078 441978
rect 517134 441922 517202 441978
rect 517258 441922 517328 441978
rect 517008 441888 517328 441922
rect 527658 436350 528278 453922
rect 527658 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 528278 436350
rect 527658 436226 528278 436294
rect 527658 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 528278 436226
rect 527658 436102 528278 436170
rect 527658 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 528278 436102
rect 527658 435978 528278 436046
rect 527658 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 528278 435978
rect 517008 424350 517328 424384
rect 517008 424294 517078 424350
rect 517134 424294 517202 424350
rect 517258 424294 517328 424350
rect 517008 424226 517328 424294
rect 517008 424170 517078 424226
rect 517134 424170 517202 424226
rect 517258 424170 517328 424226
rect 517008 424102 517328 424170
rect 517008 424046 517078 424102
rect 517134 424046 517202 424102
rect 517258 424046 517328 424102
rect 517008 423978 517328 424046
rect 517008 423922 517078 423978
rect 517134 423922 517202 423978
rect 517258 423922 517328 423978
rect 517008 423888 517328 423922
rect 527658 418350 528278 435922
rect 527658 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 528278 418350
rect 527658 418226 528278 418294
rect 527658 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 528278 418226
rect 527658 418102 528278 418170
rect 527658 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 528278 418102
rect 527658 417978 528278 418046
rect 527658 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 528278 417978
rect 514892 409552 514948 409562
rect 519148 409978 519204 409988
rect 519148 398132 519204 409922
rect 519148 398066 519204 398076
rect 527658 400350 528278 417922
rect 527658 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 528278 400350
rect 527658 400226 528278 400294
rect 527658 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 528278 400226
rect 527658 400102 528278 400170
rect 527658 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 528278 400102
rect 527658 399978 528278 400046
rect 527658 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 528278 399978
rect 511420 397282 511476 397292
rect 526428 397198 526484 397208
rect 526428 396900 526484 397142
rect 526428 396834 526484 396844
rect 527658 394038 528278 399922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 531378 568350 531998 585922
rect 531378 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 531998 568350
rect 531378 568226 531998 568294
rect 531378 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 531998 568226
rect 531378 568102 531998 568170
rect 531378 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 531998 568102
rect 531378 567978 531998 568046
rect 531378 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 531998 567978
rect 531378 550350 531998 567922
rect 558378 597212 558998 598268
rect 558378 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 558998 597212
rect 558378 597088 558998 597156
rect 558378 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 558998 597088
rect 558378 596964 558998 597032
rect 558378 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 558998 596964
rect 558378 596840 558998 596908
rect 558378 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 558998 596840
rect 558378 580350 558998 596784
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 558378 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 558998 580350
rect 558378 580226 558998 580294
rect 558378 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 558998 580226
rect 558378 580102 558998 580170
rect 558378 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 558998 580102
rect 558378 579978 558998 580046
rect 558378 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 558998 579978
rect 556108 565124 556164 565134
rect 532368 562350 532688 562384
rect 532368 562294 532438 562350
rect 532494 562294 532562 562350
rect 532618 562294 532688 562350
rect 532368 562226 532688 562294
rect 532368 562170 532438 562226
rect 532494 562170 532562 562226
rect 532618 562170 532688 562226
rect 532368 562102 532688 562170
rect 532368 562046 532438 562102
rect 532494 562046 532562 562102
rect 532618 562046 532688 562102
rect 532368 561978 532688 562046
rect 532368 561922 532438 561978
rect 532494 561922 532562 561978
rect 532618 561922 532688 561978
rect 532368 561888 532688 561922
rect 552748 555716 552804 555726
rect 531378 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 531998 550350
rect 531378 550226 531998 550294
rect 531378 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 531998 550226
rect 531378 550102 531998 550170
rect 531378 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 531998 550102
rect 531378 549978 531998 550046
rect 531378 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 531998 549978
rect 531378 532350 531998 549922
rect 547728 550350 548048 550384
rect 547728 550294 547798 550350
rect 547854 550294 547922 550350
rect 547978 550294 548048 550350
rect 547728 550226 548048 550294
rect 547728 550170 547798 550226
rect 547854 550170 547922 550226
rect 547978 550170 548048 550226
rect 547728 550102 548048 550170
rect 547728 550046 547798 550102
rect 547854 550046 547922 550102
rect 547978 550046 548048 550102
rect 547728 549978 548048 550046
rect 547728 549922 547798 549978
rect 547854 549922 547922 549978
rect 547978 549922 548048 549978
rect 547728 549888 548048 549922
rect 532368 544350 532688 544384
rect 532368 544294 532438 544350
rect 532494 544294 532562 544350
rect 532618 544294 532688 544350
rect 532368 544226 532688 544294
rect 532368 544170 532438 544226
rect 532494 544170 532562 544226
rect 532618 544170 532688 544226
rect 532368 544102 532688 544170
rect 532368 544046 532438 544102
rect 532494 544046 532562 544102
rect 532618 544046 532688 544102
rect 532368 543978 532688 544046
rect 532368 543922 532438 543978
rect 532494 543922 532562 543978
rect 532618 543922 532688 543978
rect 532368 543888 532688 543922
rect 531378 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 531998 532350
rect 531378 532226 531998 532294
rect 531378 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 531998 532226
rect 531378 532102 531998 532170
rect 531378 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 531998 532102
rect 531378 531978 531998 532046
rect 531378 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 531998 531978
rect 531378 514350 531998 531922
rect 547728 532350 548048 532384
rect 547728 532294 547798 532350
rect 547854 532294 547922 532350
rect 547978 532294 548048 532350
rect 547728 532226 548048 532294
rect 547728 532170 547798 532226
rect 547854 532170 547922 532226
rect 547978 532170 548048 532226
rect 547728 532102 548048 532170
rect 547728 532046 547798 532102
rect 547854 532046 547922 532102
rect 547978 532046 548048 532102
rect 547728 531978 548048 532046
rect 547728 531922 547798 531978
rect 547854 531922 547922 531978
rect 547978 531922 548048 531978
rect 547728 531888 548048 531922
rect 532368 526350 532688 526384
rect 532368 526294 532438 526350
rect 532494 526294 532562 526350
rect 532618 526294 532688 526350
rect 532368 526226 532688 526294
rect 532368 526170 532438 526226
rect 532494 526170 532562 526226
rect 532618 526170 532688 526226
rect 532368 526102 532688 526170
rect 532368 526046 532438 526102
rect 532494 526046 532562 526102
rect 532618 526046 532688 526102
rect 532368 525978 532688 526046
rect 532368 525922 532438 525978
rect 532494 525922 532562 525978
rect 532618 525922 532688 525978
rect 532368 525888 532688 525922
rect 549388 522788 549444 522798
rect 531378 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 531998 514350
rect 531378 514226 531998 514294
rect 531378 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 531998 514226
rect 531378 514102 531998 514170
rect 531378 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 531998 514102
rect 531378 513978 531998 514046
rect 531378 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 531998 513978
rect 531378 496350 531998 513922
rect 547728 514350 548048 514384
rect 547728 514294 547798 514350
rect 547854 514294 547922 514350
rect 547978 514294 548048 514350
rect 547728 514226 548048 514294
rect 547728 514170 547798 514226
rect 547854 514170 547922 514226
rect 547978 514170 548048 514226
rect 547728 514102 548048 514170
rect 547728 514046 547798 514102
rect 547854 514046 547922 514102
rect 547978 514046 548048 514102
rect 547728 513978 548048 514046
rect 547728 513922 547798 513978
rect 547854 513922 547922 513978
rect 547978 513922 548048 513978
rect 547728 513888 548048 513922
rect 532368 508350 532688 508384
rect 532368 508294 532438 508350
rect 532494 508294 532562 508350
rect 532618 508294 532688 508350
rect 532368 508226 532688 508294
rect 532368 508170 532438 508226
rect 532494 508170 532562 508226
rect 532618 508170 532688 508226
rect 532368 508102 532688 508170
rect 532368 508046 532438 508102
rect 532494 508046 532562 508102
rect 532618 508046 532688 508102
rect 532368 507978 532688 508046
rect 532368 507922 532438 507978
rect 532494 507922 532562 507978
rect 532618 507922 532688 507978
rect 532368 507888 532688 507922
rect 531378 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 531998 496350
rect 531378 496226 531998 496294
rect 531378 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 531998 496226
rect 531378 496102 531998 496170
rect 531378 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 531998 496102
rect 531378 495978 531998 496046
rect 531378 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 531998 495978
rect 531378 478350 531998 495922
rect 547728 496350 548048 496384
rect 547728 496294 547798 496350
rect 547854 496294 547922 496350
rect 547978 496294 548048 496350
rect 547728 496226 548048 496294
rect 547728 496170 547798 496226
rect 547854 496170 547922 496226
rect 547978 496170 548048 496226
rect 547728 496102 548048 496170
rect 547728 496046 547798 496102
rect 547854 496046 547922 496102
rect 547978 496046 548048 496102
rect 547728 495978 548048 496046
rect 547728 495922 547798 495978
rect 547854 495922 547922 495978
rect 547978 495922 548048 495978
rect 547728 495888 548048 495922
rect 532368 490350 532688 490384
rect 532368 490294 532438 490350
rect 532494 490294 532562 490350
rect 532618 490294 532688 490350
rect 532368 490226 532688 490294
rect 532368 490170 532438 490226
rect 532494 490170 532562 490226
rect 532618 490170 532688 490226
rect 532368 490102 532688 490170
rect 532368 490046 532438 490102
rect 532494 490046 532562 490102
rect 532618 490046 532688 490102
rect 532368 489978 532688 490046
rect 532368 489922 532438 489978
rect 532494 489922 532562 489978
rect 532618 489922 532688 489978
rect 532368 489888 532688 489922
rect 531378 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 531998 478350
rect 531378 478226 531998 478294
rect 531378 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 531998 478226
rect 531378 478102 531998 478170
rect 531378 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 531998 478102
rect 531378 477978 531998 478046
rect 531378 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 531998 477978
rect 531378 460350 531998 477922
rect 547728 478350 548048 478384
rect 547728 478294 547798 478350
rect 547854 478294 547922 478350
rect 547978 478294 548048 478350
rect 547728 478226 548048 478294
rect 547728 478170 547798 478226
rect 547854 478170 547922 478226
rect 547978 478170 548048 478226
rect 547728 478102 548048 478170
rect 547728 478046 547798 478102
rect 547854 478046 547922 478102
rect 547978 478046 548048 478102
rect 547728 477978 548048 478046
rect 547728 477922 547798 477978
rect 547854 477922 547922 477978
rect 547978 477922 548048 477978
rect 547728 477888 548048 477922
rect 532368 472350 532688 472384
rect 532368 472294 532438 472350
rect 532494 472294 532562 472350
rect 532618 472294 532688 472350
rect 532368 472226 532688 472294
rect 532368 472170 532438 472226
rect 532494 472170 532562 472226
rect 532618 472170 532688 472226
rect 532368 472102 532688 472170
rect 532368 472046 532438 472102
rect 532494 472046 532562 472102
rect 532618 472046 532688 472102
rect 532368 471978 532688 472046
rect 532368 471922 532438 471978
rect 532494 471922 532562 471978
rect 532618 471922 532688 471978
rect 532368 471888 532688 471922
rect 531378 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 531998 460350
rect 531378 460226 531998 460294
rect 531378 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 531998 460226
rect 531378 460102 531998 460170
rect 531378 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 531998 460102
rect 531378 459978 531998 460046
rect 531378 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 531998 459978
rect 531378 442350 531998 459922
rect 547728 460350 548048 460384
rect 547728 460294 547798 460350
rect 547854 460294 547922 460350
rect 547978 460294 548048 460350
rect 547728 460226 548048 460294
rect 547728 460170 547798 460226
rect 547854 460170 547922 460226
rect 547978 460170 548048 460226
rect 547728 460102 548048 460170
rect 547728 460046 547798 460102
rect 547854 460046 547922 460102
rect 547978 460046 548048 460102
rect 547728 459978 548048 460046
rect 547728 459922 547798 459978
rect 547854 459922 547922 459978
rect 547978 459922 548048 459978
rect 547728 459888 548048 459922
rect 532368 454350 532688 454384
rect 532368 454294 532438 454350
rect 532494 454294 532562 454350
rect 532618 454294 532688 454350
rect 532368 454226 532688 454294
rect 532368 454170 532438 454226
rect 532494 454170 532562 454226
rect 532618 454170 532688 454226
rect 532368 454102 532688 454170
rect 532368 454046 532438 454102
rect 532494 454046 532562 454102
rect 532618 454046 532688 454102
rect 532368 453978 532688 454046
rect 532368 453922 532438 453978
rect 532494 453922 532562 453978
rect 532618 453922 532688 453978
rect 532368 453888 532688 453922
rect 531378 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 531998 442350
rect 531378 442226 531998 442294
rect 531378 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 531998 442226
rect 531378 442102 531998 442170
rect 531378 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 531998 442102
rect 531378 441978 531998 442046
rect 531378 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 531998 441978
rect 531378 424350 531998 441922
rect 547728 442350 548048 442384
rect 547728 442294 547798 442350
rect 547854 442294 547922 442350
rect 547978 442294 548048 442350
rect 547728 442226 548048 442294
rect 547728 442170 547798 442226
rect 547854 442170 547922 442226
rect 547978 442170 548048 442226
rect 547728 442102 548048 442170
rect 547728 442046 547798 442102
rect 547854 442046 547922 442102
rect 547978 442046 548048 442102
rect 547728 441978 548048 442046
rect 547728 441922 547798 441978
rect 547854 441922 547922 441978
rect 547978 441922 548048 441978
rect 547728 441888 548048 441922
rect 532368 436350 532688 436384
rect 532368 436294 532438 436350
rect 532494 436294 532562 436350
rect 532618 436294 532688 436350
rect 532368 436226 532688 436294
rect 532368 436170 532438 436226
rect 532494 436170 532562 436226
rect 532618 436170 532688 436226
rect 532368 436102 532688 436170
rect 532368 436046 532438 436102
rect 532494 436046 532562 436102
rect 532618 436046 532688 436102
rect 532368 435978 532688 436046
rect 532368 435922 532438 435978
rect 532494 435922 532562 435978
rect 532618 435922 532688 435978
rect 532368 435888 532688 435922
rect 531378 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 531998 424350
rect 531378 424226 531998 424294
rect 531378 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 531998 424226
rect 531378 424102 531998 424170
rect 531378 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 531998 424102
rect 531378 423978 531998 424046
rect 531378 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 531998 423978
rect 531378 406350 531998 423922
rect 547728 424350 548048 424384
rect 547728 424294 547798 424350
rect 547854 424294 547922 424350
rect 547978 424294 548048 424350
rect 547728 424226 548048 424294
rect 547728 424170 547798 424226
rect 547854 424170 547922 424226
rect 547978 424170 548048 424226
rect 547728 424102 548048 424170
rect 547728 424046 547798 424102
rect 547854 424046 547922 424102
rect 547978 424046 548048 424102
rect 547728 423978 548048 424046
rect 547728 423922 547798 423978
rect 547854 423922 547922 423978
rect 547978 423922 548048 423978
rect 547728 423888 548048 423922
rect 532368 418350 532688 418384
rect 532368 418294 532438 418350
rect 532494 418294 532562 418350
rect 532618 418294 532688 418350
rect 532368 418226 532688 418294
rect 532368 418170 532438 418226
rect 532494 418170 532562 418226
rect 532618 418170 532688 418226
rect 532368 418102 532688 418170
rect 532368 418046 532438 418102
rect 532494 418046 532562 418102
rect 532618 418046 532688 418102
rect 532368 417978 532688 418046
rect 532368 417922 532438 417978
rect 532494 417922 532562 417978
rect 532618 417922 532688 417978
rect 532368 417888 532688 417922
rect 533820 407652 533876 407662
rect 533820 407098 533876 407596
rect 533820 407032 533876 407042
rect 539196 407652 539252 407662
rect 539196 406918 539252 407596
rect 539196 406852 539252 406862
rect 531378 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 531998 406350
rect 531378 406226 531998 406294
rect 531378 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 531998 406226
rect 531378 406102 531998 406170
rect 531378 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 531998 406102
rect 531378 405978 531998 406046
rect 531378 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 531998 405978
rect 531378 394038 531998 405922
rect 549388 400618 549444 522732
rect 551068 494564 551124 494574
rect 549388 400552 549444 400562
rect 549500 489860 549556 489870
rect 549500 398998 549556 489804
rect 551068 399178 551124 494508
rect 551180 414596 551236 414606
rect 551180 407458 551236 414540
rect 551180 407392 551236 407402
rect 552748 405658 552804 555660
rect 556108 410878 556164 565068
rect 558378 562350 558998 579922
rect 558378 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 558998 562350
rect 558378 562226 558998 562294
rect 558378 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 558998 562226
rect 558378 562102 558998 562170
rect 558378 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 558998 562102
rect 558378 561978 558998 562046
rect 558378 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 558998 561978
rect 556108 410812 556164 410822
rect 556220 551012 556276 551022
rect 556220 409258 556276 550956
rect 558378 544350 558998 561922
rect 558378 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 558998 544350
rect 558378 544226 558998 544294
rect 558378 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 558998 544226
rect 558378 544102 558998 544170
rect 558378 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 558998 544102
rect 558378 543978 558998 544046
rect 558378 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 558998 543978
rect 556444 536900 556500 536910
rect 556220 409192 556276 409202
rect 556332 527492 556388 527502
rect 552748 405592 552804 405602
rect 556332 399358 556388 527436
rect 556444 410698 556500 536844
rect 556444 410632 556500 410642
rect 558378 526350 558998 543922
rect 558378 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 558998 526350
rect 558378 526226 558998 526294
rect 558378 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 558998 526226
rect 558378 526102 558998 526170
rect 558378 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 558998 526102
rect 558378 525978 558998 526046
rect 558378 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 558998 525978
rect 558378 508350 558998 525922
rect 558378 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 558998 508350
rect 558378 508226 558998 508294
rect 558378 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 558998 508226
rect 558378 508102 558998 508170
rect 558378 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 558998 508102
rect 558378 507978 558998 508046
rect 558378 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 558998 507978
rect 558378 490350 558998 507922
rect 558378 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 558998 490350
rect 558378 490226 558998 490294
rect 558378 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 558998 490226
rect 558378 490102 558998 490170
rect 558378 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 558998 490102
rect 558378 489978 558998 490046
rect 558378 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 558998 489978
rect 558378 472350 558998 489922
rect 558378 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 558998 472350
rect 558378 472226 558998 472294
rect 558378 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 558998 472226
rect 558378 472102 558998 472170
rect 558378 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 558998 472102
rect 558378 471978 558998 472046
rect 558378 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 558998 471978
rect 558378 454350 558998 471922
rect 558378 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 558998 454350
rect 558378 454226 558998 454294
rect 558378 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 558998 454226
rect 558378 454102 558998 454170
rect 558378 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 558998 454102
rect 558378 453978 558998 454046
rect 558378 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 558998 453978
rect 558378 436350 558998 453922
rect 558378 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 558998 436350
rect 558378 436226 558998 436294
rect 558378 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 558998 436226
rect 558378 436102 558998 436170
rect 558378 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 558998 436102
rect 558378 435978 558998 436046
rect 558378 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 558998 435978
rect 558378 418350 558998 435922
rect 558378 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 558998 418350
rect 558378 418226 558998 418294
rect 558378 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 558998 418226
rect 558378 418102 558998 418170
rect 558378 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 558998 418102
rect 558378 417978 558998 418046
rect 558378 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 558998 417978
rect 557788 407428 557844 407438
rect 557788 406738 557844 407372
rect 557788 406672 557844 406682
rect 556332 399292 556388 399302
rect 558378 400350 558998 417922
rect 560252 591332 560308 591342
rect 560252 404578 560308 591276
rect 560252 404512 560308 404522
rect 562098 586350 562718 597744
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 568350 562718 585922
rect 562098 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 562718 568350
rect 562098 568226 562718 568294
rect 562098 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 562718 568226
rect 562098 568102 562718 568170
rect 562098 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 562718 568102
rect 562098 567978 562718 568046
rect 562098 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 562718 567978
rect 562098 550350 562718 567922
rect 562098 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 562718 550350
rect 562098 550226 562718 550294
rect 562098 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 562718 550226
rect 562098 550102 562718 550170
rect 562098 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 562718 550102
rect 562098 549978 562718 550046
rect 562098 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 562718 549978
rect 562098 532350 562718 549922
rect 584668 590212 584724 590222
rect 562098 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 562718 532350
rect 562098 532226 562718 532294
rect 562098 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 562718 532226
rect 562098 532102 562718 532170
rect 562098 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 562718 532102
rect 562098 531978 562718 532046
rect 562098 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 562718 531978
rect 562098 514350 562718 531922
rect 562098 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 562718 514350
rect 562098 514226 562718 514294
rect 562098 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 562718 514226
rect 562098 514102 562718 514170
rect 562098 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 562718 514102
rect 562098 513978 562718 514046
rect 562098 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 562718 513978
rect 562098 496350 562718 513922
rect 562098 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 562718 496350
rect 562098 496226 562718 496294
rect 562098 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 562718 496226
rect 562098 496102 562718 496170
rect 562098 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 562718 496102
rect 562098 495978 562718 496046
rect 562098 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 562718 495978
rect 562098 478350 562718 495922
rect 562098 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 562718 478350
rect 562098 478226 562718 478294
rect 562098 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 562718 478226
rect 562098 478102 562718 478170
rect 562098 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 562718 478102
rect 562098 477978 562718 478046
rect 562098 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 562718 477978
rect 562098 460350 562718 477922
rect 562098 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 562718 460350
rect 562098 460226 562718 460294
rect 562098 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 562718 460226
rect 562098 460102 562718 460170
rect 562098 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 562718 460102
rect 562098 459978 562718 460046
rect 562098 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 562718 459978
rect 562098 442350 562718 459922
rect 562098 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 562718 442350
rect 562098 442226 562718 442294
rect 562098 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 562718 442226
rect 562098 442102 562718 442170
rect 562098 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 562718 442102
rect 562098 441978 562718 442046
rect 562098 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 562718 441978
rect 562098 424350 562718 441922
rect 562098 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 562718 424350
rect 562098 424226 562718 424294
rect 562098 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 562718 424226
rect 562098 424102 562718 424170
rect 562098 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 562718 424102
rect 562098 423978 562718 424046
rect 562098 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 562718 423978
rect 562098 406350 562718 423922
rect 562098 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 562718 406350
rect 562098 406226 562718 406294
rect 562098 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 562718 406226
rect 562098 406102 562718 406170
rect 562098 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 562718 406102
rect 562098 405978 562718 406046
rect 562098 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 562718 405978
rect 558378 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 558998 400350
rect 558378 400226 558998 400294
rect 558378 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 558998 400226
rect 558378 400102 558998 400170
rect 558378 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 558998 400102
rect 558378 399978 558998 400046
rect 558378 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 558998 399978
rect 551068 399112 551124 399122
rect 549500 398932 549556 398942
rect 532476 397018 532532 397028
rect 532476 396788 532532 396962
rect 532476 396722 532532 396732
rect 556668 396838 556724 396848
rect 556668 396676 556724 396782
rect 550620 396658 550676 396668
rect 556668 396610 556724 396620
rect 550620 396564 550676 396602
rect 550620 396498 550676 396508
rect 538524 394884 538580 394894
rect 538524 394790 538580 394802
rect 558378 394038 558998 399922
rect 559468 398278 559524 398288
rect 471996 392354 472052 392364
rect 362124 392308 362180 392318
rect 441756 392272 441812 392282
rect 362124 391798 362180 392252
rect 362124 391732 362180 391742
rect 379808 388350 380128 388384
rect 379808 388294 379878 388350
rect 379934 388294 380002 388350
rect 380058 388294 380128 388350
rect 379808 388226 380128 388294
rect 379808 388170 379878 388226
rect 379934 388170 380002 388226
rect 380058 388170 380128 388226
rect 379808 388102 380128 388170
rect 379808 388046 379878 388102
rect 379934 388046 380002 388102
rect 380058 388046 380128 388102
rect 379808 387978 380128 388046
rect 379808 387922 379878 387978
rect 379934 387922 380002 387978
rect 380058 387922 380128 387978
rect 379808 387888 380128 387922
rect 410528 388350 410848 388384
rect 410528 388294 410598 388350
rect 410654 388294 410722 388350
rect 410778 388294 410848 388350
rect 410528 388226 410848 388294
rect 410528 388170 410598 388226
rect 410654 388170 410722 388226
rect 410778 388170 410848 388226
rect 410528 388102 410848 388170
rect 410528 388046 410598 388102
rect 410654 388046 410722 388102
rect 410778 388046 410848 388102
rect 410528 387978 410848 388046
rect 410528 387922 410598 387978
rect 410654 387922 410722 387978
rect 410778 387922 410848 387978
rect 410528 387888 410848 387922
rect 441248 388350 441568 388384
rect 441248 388294 441318 388350
rect 441374 388294 441442 388350
rect 441498 388294 441568 388350
rect 441248 388226 441568 388294
rect 441248 388170 441318 388226
rect 441374 388170 441442 388226
rect 441498 388170 441568 388226
rect 441248 388102 441568 388170
rect 441248 388046 441318 388102
rect 441374 388046 441442 388102
rect 441498 388046 441568 388102
rect 441248 387978 441568 388046
rect 441248 387922 441318 387978
rect 441374 387922 441442 387978
rect 441498 387922 441568 387978
rect 441248 387888 441568 387922
rect 471968 388350 472288 388384
rect 471968 388294 472038 388350
rect 472094 388294 472162 388350
rect 472218 388294 472288 388350
rect 471968 388226 472288 388294
rect 471968 388170 472038 388226
rect 472094 388170 472162 388226
rect 472218 388170 472288 388226
rect 471968 388102 472288 388170
rect 471968 388046 472038 388102
rect 472094 388046 472162 388102
rect 472218 388046 472288 388102
rect 471968 387978 472288 388046
rect 471968 387922 472038 387978
rect 472094 387922 472162 387978
rect 472218 387922 472288 387978
rect 471968 387888 472288 387922
rect 502688 388350 503008 388384
rect 502688 388294 502758 388350
rect 502814 388294 502882 388350
rect 502938 388294 503008 388350
rect 502688 388226 503008 388294
rect 502688 388170 502758 388226
rect 502814 388170 502882 388226
rect 502938 388170 503008 388226
rect 502688 388102 503008 388170
rect 502688 388046 502758 388102
rect 502814 388046 502882 388102
rect 502938 388046 503008 388102
rect 502688 387978 503008 388046
rect 502688 387922 502758 387978
rect 502814 387922 502882 387978
rect 502938 387922 503008 387978
rect 502688 387888 503008 387922
rect 533408 388350 533728 388384
rect 533408 388294 533478 388350
rect 533534 388294 533602 388350
rect 533658 388294 533728 388350
rect 533408 388226 533728 388294
rect 533408 388170 533478 388226
rect 533534 388170 533602 388226
rect 533658 388170 533728 388226
rect 533408 388102 533728 388170
rect 533408 388046 533478 388102
rect 533534 388046 533602 388102
rect 533658 388046 533728 388102
rect 533408 387978 533728 388046
rect 533408 387922 533478 387978
rect 533534 387922 533602 387978
rect 533658 387922 533728 387978
rect 533408 387888 533728 387922
rect 362012 384692 362180 384748
rect 362124 383158 362180 384692
rect 362124 383092 362180 383102
rect 364448 382350 364768 382384
rect 364448 382294 364518 382350
rect 364574 382294 364642 382350
rect 364698 382294 364768 382350
rect 364448 382226 364768 382294
rect 364448 382170 364518 382226
rect 364574 382170 364642 382226
rect 364698 382170 364768 382226
rect 364448 382102 364768 382170
rect 364448 382046 364518 382102
rect 364574 382046 364642 382102
rect 364698 382046 364768 382102
rect 364448 381978 364768 382046
rect 364448 381922 364518 381978
rect 364574 381922 364642 381978
rect 364698 381922 364768 381978
rect 364448 381888 364768 381922
rect 395168 382350 395488 382384
rect 395168 382294 395238 382350
rect 395294 382294 395362 382350
rect 395418 382294 395488 382350
rect 395168 382226 395488 382294
rect 395168 382170 395238 382226
rect 395294 382170 395362 382226
rect 395418 382170 395488 382226
rect 395168 382102 395488 382170
rect 395168 382046 395238 382102
rect 395294 382046 395362 382102
rect 395418 382046 395488 382102
rect 395168 381978 395488 382046
rect 395168 381922 395238 381978
rect 395294 381922 395362 381978
rect 395418 381922 395488 381978
rect 395168 381888 395488 381922
rect 425888 382350 426208 382384
rect 425888 382294 425958 382350
rect 426014 382294 426082 382350
rect 426138 382294 426208 382350
rect 425888 382226 426208 382294
rect 425888 382170 425958 382226
rect 426014 382170 426082 382226
rect 426138 382170 426208 382226
rect 425888 382102 426208 382170
rect 425888 382046 425958 382102
rect 426014 382046 426082 382102
rect 426138 382046 426208 382102
rect 425888 381978 426208 382046
rect 425888 381922 425958 381978
rect 426014 381922 426082 381978
rect 426138 381922 426208 381978
rect 425888 381888 426208 381922
rect 456608 382350 456928 382384
rect 456608 382294 456678 382350
rect 456734 382294 456802 382350
rect 456858 382294 456928 382350
rect 456608 382226 456928 382294
rect 456608 382170 456678 382226
rect 456734 382170 456802 382226
rect 456858 382170 456928 382226
rect 456608 382102 456928 382170
rect 456608 382046 456678 382102
rect 456734 382046 456802 382102
rect 456858 382046 456928 382102
rect 456608 381978 456928 382046
rect 456608 381922 456678 381978
rect 456734 381922 456802 381978
rect 456858 381922 456928 381978
rect 456608 381888 456928 381922
rect 487328 382350 487648 382384
rect 487328 382294 487398 382350
rect 487454 382294 487522 382350
rect 487578 382294 487648 382350
rect 487328 382226 487648 382294
rect 487328 382170 487398 382226
rect 487454 382170 487522 382226
rect 487578 382170 487648 382226
rect 487328 382102 487648 382170
rect 487328 382046 487398 382102
rect 487454 382046 487522 382102
rect 487578 382046 487648 382102
rect 487328 381978 487648 382046
rect 487328 381922 487398 381978
rect 487454 381922 487522 381978
rect 487578 381922 487648 381978
rect 487328 381888 487648 381922
rect 518048 382350 518368 382384
rect 518048 382294 518118 382350
rect 518174 382294 518242 382350
rect 518298 382294 518368 382350
rect 518048 382226 518368 382294
rect 518048 382170 518118 382226
rect 518174 382170 518242 382226
rect 518298 382170 518368 382226
rect 518048 382102 518368 382170
rect 518048 382046 518118 382102
rect 518174 382046 518242 382102
rect 518298 382046 518368 382102
rect 518048 381978 518368 382046
rect 518048 381922 518118 381978
rect 518174 381922 518242 381978
rect 518298 381922 518368 381978
rect 518048 381888 518368 381922
rect 548768 382350 549088 382384
rect 548768 382294 548838 382350
rect 548894 382294 548962 382350
rect 549018 382294 549088 382350
rect 548768 382226 549088 382294
rect 548768 382170 548838 382226
rect 548894 382170 548962 382226
rect 549018 382170 549088 382226
rect 548768 382102 549088 382170
rect 548768 382046 548838 382102
rect 548894 382046 548962 382102
rect 549018 382046 549088 382102
rect 548768 381978 549088 382046
rect 548768 381922 548838 381978
rect 548894 381922 548962 381978
rect 549018 381922 549088 381978
rect 548768 381888 549088 381922
rect 379808 370350 380128 370384
rect 379808 370294 379878 370350
rect 379934 370294 380002 370350
rect 380058 370294 380128 370350
rect 379808 370226 380128 370294
rect 379808 370170 379878 370226
rect 379934 370170 380002 370226
rect 380058 370170 380128 370226
rect 379808 370102 380128 370170
rect 379808 370046 379878 370102
rect 379934 370046 380002 370102
rect 380058 370046 380128 370102
rect 379808 369978 380128 370046
rect 379808 369922 379878 369978
rect 379934 369922 380002 369978
rect 380058 369922 380128 369978
rect 379808 369888 380128 369922
rect 410528 370350 410848 370384
rect 410528 370294 410598 370350
rect 410654 370294 410722 370350
rect 410778 370294 410848 370350
rect 410528 370226 410848 370294
rect 410528 370170 410598 370226
rect 410654 370170 410722 370226
rect 410778 370170 410848 370226
rect 410528 370102 410848 370170
rect 410528 370046 410598 370102
rect 410654 370046 410722 370102
rect 410778 370046 410848 370102
rect 410528 369978 410848 370046
rect 410528 369922 410598 369978
rect 410654 369922 410722 369978
rect 410778 369922 410848 369978
rect 410528 369888 410848 369922
rect 441248 370350 441568 370384
rect 441248 370294 441318 370350
rect 441374 370294 441442 370350
rect 441498 370294 441568 370350
rect 441248 370226 441568 370294
rect 441248 370170 441318 370226
rect 441374 370170 441442 370226
rect 441498 370170 441568 370226
rect 441248 370102 441568 370170
rect 441248 370046 441318 370102
rect 441374 370046 441442 370102
rect 441498 370046 441568 370102
rect 441248 369978 441568 370046
rect 441248 369922 441318 369978
rect 441374 369922 441442 369978
rect 441498 369922 441568 369978
rect 441248 369888 441568 369922
rect 471968 370350 472288 370384
rect 471968 370294 472038 370350
rect 472094 370294 472162 370350
rect 472218 370294 472288 370350
rect 471968 370226 472288 370294
rect 471968 370170 472038 370226
rect 472094 370170 472162 370226
rect 472218 370170 472288 370226
rect 471968 370102 472288 370170
rect 471968 370046 472038 370102
rect 472094 370046 472162 370102
rect 472218 370046 472288 370102
rect 471968 369978 472288 370046
rect 471968 369922 472038 369978
rect 472094 369922 472162 369978
rect 472218 369922 472288 369978
rect 471968 369888 472288 369922
rect 502688 370350 503008 370384
rect 502688 370294 502758 370350
rect 502814 370294 502882 370350
rect 502938 370294 503008 370350
rect 502688 370226 503008 370294
rect 502688 370170 502758 370226
rect 502814 370170 502882 370226
rect 502938 370170 503008 370226
rect 502688 370102 503008 370170
rect 502688 370046 502758 370102
rect 502814 370046 502882 370102
rect 502938 370046 503008 370102
rect 502688 369978 503008 370046
rect 502688 369922 502758 369978
rect 502814 369922 502882 369978
rect 502938 369922 503008 369978
rect 502688 369888 503008 369922
rect 533408 370350 533728 370384
rect 533408 370294 533478 370350
rect 533534 370294 533602 370350
rect 533658 370294 533728 370350
rect 533408 370226 533728 370294
rect 533408 370170 533478 370226
rect 533534 370170 533602 370226
rect 533658 370170 533728 370226
rect 533408 370102 533728 370170
rect 533408 370046 533478 370102
rect 533534 370046 533602 370102
rect 533658 370046 533728 370102
rect 533408 369978 533728 370046
rect 533408 369922 533478 369978
rect 533534 369922 533602 369978
rect 533658 369922 533728 369978
rect 533408 369888 533728 369922
rect 364448 364350 364768 364384
rect 364448 364294 364518 364350
rect 364574 364294 364642 364350
rect 364698 364294 364768 364350
rect 364448 364226 364768 364294
rect 364448 364170 364518 364226
rect 364574 364170 364642 364226
rect 364698 364170 364768 364226
rect 364448 364102 364768 364170
rect 364448 364046 364518 364102
rect 364574 364046 364642 364102
rect 364698 364046 364768 364102
rect 364448 363978 364768 364046
rect 364448 363922 364518 363978
rect 364574 363922 364642 363978
rect 364698 363922 364768 363978
rect 364448 363888 364768 363922
rect 395168 364350 395488 364384
rect 395168 364294 395238 364350
rect 395294 364294 395362 364350
rect 395418 364294 395488 364350
rect 395168 364226 395488 364294
rect 395168 364170 395238 364226
rect 395294 364170 395362 364226
rect 395418 364170 395488 364226
rect 395168 364102 395488 364170
rect 395168 364046 395238 364102
rect 395294 364046 395362 364102
rect 395418 364046 395488 364102
rect 395168 363978 395488 364046
rect 395168 363922 395238 363978
rect 395294 363922 395362 363978
rect 395418 363922 395488 363978
rect 395168 363888 395488 363922
rect 425888 364350 426208 364384
rect 425888 364294 425958 364350
rect 426014 364294 426082 364350
rect 426138 364294 426208 364350
rect 425888 364226 426208 364294
rect 425888 364170 425958 364226
rect 426014 364170 426082 364226
rect 426138 364170 426208 364226
rect 425888 364102 426208 364170
rect 425888 364046 425958 364102
rect 426014 364046 426082 364102
rect 426138 364046 426208 364102
rect 425888 363978 426208 364046
rect 425888 363922 425958 363978
rect 426014 363922 426082 363978
rect 426138 363922 426208 363978
rect 425888 363888 426208 363922
rect 456608 364350 456928 364384
rect 456608 364294 456678 364350
rect 456734 364294 456802 364350
rect 456858 364294 456928 364350
rect 456608 364226 456928 364294
rect 456608 364170 456678 364226
rect 456734 364170 456802 364226
rect 456858 364170 456928 364226
rect 456608 364102 456928 364170
rect 456608 364046 456678 364102
rect 456734 364046 456802 364102
rect 456858 364046 456928 364102
rect 456608 363978 456928 364046
rect 456608 363922 456678 363978
rect 456734 363922 456802 363978
rect 456858 363922 456928 363978
rect 456608 363888 456928 363922
rect 487328 364350 487648 364384
rect 487328 364294 487398 364350
rect 487454 364294 487522 364350
rect 487578 364294 487648 364350
rect 487328 364226 487648 364294
rect 487328 364170 487398 364226
rect 487454 364170 487522 364226
rect 487578 364170 487648 364226
rect 487328 364102 487648 364170
rect 487328 364046 487398 364102
rect 487454 364046 487522 364102
rect 487578 364046 487648 364102
rect 487328 363978 487648 364046
rect 487328 363922 487398 363978
rect 487454 363922 487522 363978
rect 487578 363922 487648 363978
rect 487328 363888 487648 363922
rect 518048 364350 518368 364384
rect 518048 364294 518118 364350
rect 518174 364294 518242 364350
rect 518298 364294 518368 364350
rect 518048 364226 518368 364294
rect 518048 364170 518118 364226
rect 518174 364170 518242 364226
rect 518298 364170 518368 364226
rect 518048 364102 518368 364170
rect 518048 364046 518118 364102
rect 518174 364046 518242 364102
rect 518298 364046 518368 364102
rect 518048 363978 518368 364046
rect 518048 363922 518118 363978
rect 518174 363922 518242 363978
rect 518298 363922 518368 363978
rect 518048 363888 518368 363922
rect 548768 364350 549088 364384
rect 548768 364294 548838 364350
rect 548894 364294 548962 364350
rect 549018 364294 549088 364350
rect 548768 364226 549088 364294
rect 548768 364170 548838 364226
rect 548894 364170 548962 364226
rect 549018 364170 549088 364226
rect 548768 364102 549088 364170
rect 548768 364046 548838 364102
rect 548894 364046 548962 364102
rect 549018 364046 549088 364102
rect 548768 363978 549088 364046
rect 548768 363922 548838 363978
rect 548894 363922 548962 363978
rect 549018 363922 549088 363978
rect 548768 363888 549088 363922
rect 379808 352350 380128 352384
rect 379808 352294 379878 352350
rect 379934 352294 380002 352350
rect 380058 352294 380128 352350
rect 379808 352226 380128 352294
rect 379808 352170 379878 352226
rect 379934 352170 380002 352226
rect 380058 352170 380128 352226
rect 379808 352102 380128 352170
rect 379808 352046 379878 352102
rect 379934 352046 380002 352102
rect 380058 352046 380128 352102
rect 379808 351978 380128 352046
rect 379808 351922 379878 351978
rect 379934 351922 380002 351978
rect 380058 351922 380128 351978
rect 379808 351888 380128 351922
rect 410528 352350 410848 352384
rect 410528 352294 410598 352350
rect 410654 352294 410722 352350
rect 410778 352294 410848 352350
rect 410528 352226 410848 352294
rect 410528 352170 410598 352226
rect 410654 352170 410722 352226
rect 410778 352170 410848 352226
rect 410528 352102 410848 352170
rect 410528 352046 410598 352102
rect 410654 352046 410722 352102
rect 410778 352046 410848 352102
rect 410528 351978 410848 352046
rect 410528 351922 410598 351978
rect 410654 351922 410722 351978
rect 410778 351922 410848 351978
rect 410528 351888 410848 351922
rect 441248 352350 441568 352384
rect 441248 352294 441318 352350
rect 441374 352294 441442 352350
rect 441498 352294 441568 352350
rect 441248 352226 441568 352294
rect 441248 352170 441318 352226
rect 441374 352170 441442 352226
rect 441498 352170 441568 352226
rect 441248 352102 441568 352170
rect 441248 352046 441318 352102
rect 441374 352046 441442 352102
rect 441498 352046 441568 352102
rect 441248 351978 441568 352046
rect 441248 351922 441318 351978
rect 441374 351922 441442 351978
rect 441498 351922 441568 351978
rect 441248 351888 441568 351922
rect 471968 352350 472288 352384
rect 471968 352294 472038 352350
rect 472094 352294 472162 352350
rect 472218 352294 472288 352350
rect 471968 352226 472288 352294
rect 471968 352170 472038 352226
rect 472094 352170 472162 352226
rect 472218 352170 472288 352226
rect 471968 352102 472288 352170
rect 471968 352046 472038 352102
rect 472094 352046 472162 352102
rect 472218 352046 472288 352102
rect 471968 351978 472288 352046
rect 471968 351922 472038 351978
rect 472094 351922 472162 351978
rect 472218 351922 472288 351978
rect 471968 351888 472288 351922
rect 502688 352350 503008 352384
rect 502688 352294 502758 352350
rect 502814 352294 502882 352350
rect 502938 352294 503008 352350
rect 502688 352226 503008 352294
rect 502688 352170 502758 352226
rect 502814 352170 502882 352226
rect 502938 352170 503008 352226
rect 502688 352102 503008 352170
rect 502688 352046 502758 352102
rect 502814 352046 502882 352102
rect 502938 352046 503008 352102
rect 502688 351978 503008 352046
rect 502688 351922 502758 351978
rect 502814 351922 502882 351978
rect 502938 351922 503008 351978
rect 502688 351888 503008 351922
rect 533408 352350 533728 352384
rect 533408 352294 533478 352350
rect 533534 352294 533602 352350
rect 533658 352294 533728 352350
rect 533408 352226 533728 352294
rect 533408 352170 533478 352226
rect 533534 352170 533602 352226
rect 533658 352170 533728 352226
rect 533408 352102 533728 352170
rect 533408 352046 533478 352102
rect 533534 352046 533602 352102
rect 533658 352046 533728 352102
rect 533408 351978 533728 352046
rect 533408 351922 533478 351978
rect 533534 351922 533602 351978
rect 533658 351922 533728 351978
rect 533408 351888 533728 351922
rect 364448 346350 364768 346384
rect 364448 346294 364518 346350
rect 364574 346294 364642 346350
rect 364698 346294 364768 346350
rect 364448 346226 364768 346294
rect 364448 346170 364518 346226
rect 364574 346170 364642 346226
rect 364698 346170 364768 346226
rect 364448 346102 364768 346170
rect 364448 346046 364518 346102
rect 364574 346046 364642 346102
rect 364698 346046 364768 346102
rect 364448 345978 364768 346046
rect 364448 345922 364518 345978
rect 364574 345922 364642 345978
rect 364698 345922 364768 345978
rect 364448 345888 364768 345922
rect 395168 346350 395488 346384
rect 395168 346294 395238 346350
rect 395294 346294 395362 346350
rect 395418 346294 395488 346350
rect 395168 346226 395488 346294
rect 395168 346170 395238 346226
rect 395294 346170 395362 346226
rect 395418 346170 395488 346226
rect 395168 346102 395488 346170
rect 395168 346046 395238 346102
rect 395294 346046 395362 346102
rect 395418 346046 395488 346102
rect 395168 345978 395488 346046
rect 395168 345922 395238 345978
rect 395294 345922 395362 345978
rect 395418 345922 395488 345978
rect 395168 345888 395488 345922
rect 425888 346350 426208 346384
rect 425888 346294 425958 346350
rect 426014 346294 426082 346350
rect 426138 346294 426208 346350
rect 425888 346226 426208 346294
rect 425888 346170 425958 346226
rect 426014 346170 426082 346226
rect 426138 346170 426208 346226
rect 425888 346102 426208 346170
rect 425888 346046 425958 346102
rect 426014 346046 426082 346102
rect 426138 346046 426208 346102
rect 425888 345978 426208 346046
rect 425888 345922 425958 345978
rect 426014 345922 426082 345978
rect 426138 345922 426208 345978
rect 425888 345888 426208 345922
rect 456608 346350 456928 346384
rect 456608 346294 456678 346350
rect 456734 346294 456802 346350
rect 456858 346294 456928 346350
rect 456608 346226 456928 346294
rect 456608 346170 456678 346226
rect 456734 346170 456802 346226
rect 456858 346170 456928 346226
rect 456608 346102 456928 346170
rect 456608 346046 456678 346102
rect 456734 346046 456802 346102
rect 456858 346046 456928 346102
rect 456608 345978 456928 346046
rect 456608 345922 456678 345978
rect 456734 345922 456802 345978
rect 456858 345922 456928 345978
rect 456608 345888 456928 345922
rect 487328 346350 487648 346384
rect 487328 346294 487398 346350
rect 487454 346294 487522 346350
rect 487578 346294 487648 346350
rect 487328 346226 487648 346294
rect 487328 346170 487398 346226
rect 487454 346170 487522 346226
rect 487578 346170 487648 346226
rect 487328 346102 487648 346170
rect 487328 346046 487398 346102
rect 487454 346046 487522 346102
rect 487578 346046 487648 346102
rect 487328 345978 487648 346046
rect 487328 345922 487398 345978
rect 487454 345922 487522 345978
rect 487578 345922 487648 345978
rect 487328 345888 487648 345922
rect 518048 346350 518368 346384
rect 518048 346294 518118 346350
rect 518174 346294 518242 346350
rect 518298 346294 518368 346350
rect 518048 346226 518368 346294
rect 518048 346170 518118 346226
rect 518174 346170 518242 346226
rect 518298 346170 518368 346226
rect 518048 346102 518368 346170
rect 518048 346046 518118 346102
rect 518174 346046 518242 346102
rect 518298 346046 518368 346102
rect 518048 345978 518368 346046
rect 518048 345922 518118 345978
rect 518174 345922 518242 345978
rect 518298 345922 518368 345978
rect 518048 345888 518368 345922
rect 548768 346350 549088 346384
rect 548768 346294 548838 346350
rect 548894 346294 548962 346350
rect 549018 346294 549088 346350
rect 548768 346226 549088 346294
rect 548768 346170 548838 346226
rect 548894 346170 548962 346226
rect 549018 346170 549088 346226
rect 548768 346102 549088 346170
rect 548768 346046 548838 346102
rect 548894 346046 548962 346102
rect 549018 346046 549088 346102
rect 548768 345978 549088 346046
rect 548768 345922 548838 345978
rect 548894 345922 548962 345978
rect 549018 345922 549088 345978
rect 548768 345888 549088 345922
rect 379808 334350 380128 334384
rect 379808 334294 379878 334350
rect 379934 334294 380002 334350
rect 380058 334294 380128 334350
rect 379808 334226 380128 334294
rect 379808 334170 379878 334226
rect 379934 334170 380002 334226
rect 380058 334170 380128 334226
rect 379808 334102 380128 334170
rect 379808 334046 379878 334102
rect 379934 334046 380002 334102
rect 380058 334046 380128 334102
rect 379808 333978 380128 334046
rect 379808 333922 379878 333978
rect 379934 333922 380002 333978
rect 380058 333922 380128 333978
rect 379808 333888 380128 333922
rect 410528 334350 410848 334384
rect 410528 334294 410598 334350
rect 410654 334294 410722 334350
rect 410778 334294 410848 334350
rect 410528 334226 410848 334294
rect 410528 334170 410598 334226
rect 410654 334170 410722 334226
rect 410778 334170 410848 334226
rect 410528 334102 410848 334170
rect 410528 334046 410598 334102
rect 410654 334046 410722 334102
rect 410778 334046 410848 334102
rect 410528 333978 410848 334046
rect 410528 333922 410598 333978
rect 410654 333922 410722 333978
rect 410778 333922 410848 333978
rect 410528 333888 410848 333922
rect 441248 334350 441568 334384
rect 441248 334294 441318 334350
rect 441374 334294 441442 334350
rect 441498 334294 441568 334350
rect 441248 334226 441568 334294
rect 441248 334170 441318 334226
rect 441374 334170 441442 334226
rect 441498 334170 441568 334226
rect 441248 334102 441568 334170
rect 441248 334046 441318 334102
rect 441374 334046 441442 334102
rect 441498 334046 441568 334102
rect 441248 333978 441568 334046
rect 441248 333922 441318 333978
rect 441374 333922 441442 333978
rect 441498 333922 441568 333978
rect 441248 333888 441568 333922
rect 471968 334350 472288 334384
rect 471968 334294 472038 334350
rect 472094 334294 472162 334350
rect 472218 334294 472288 334350
rect 471968 334226 472288 334294
rect 471968 334170 472038 334226
rect 472094 334170 472162 334226
rect 472218 334170 472288 334226
rect 471968 334102 472288 334170
rect 471968 334046 472038 334102
rect 472094 334046 472162 334102
rect 472218 334046 472288 334102
rect 471968 333978 472288 334046
rect 471968 333922 472038 333978
rect 472094 333922 472162 333978
rect 472218 333922 472288 333978
rect 471968 333888 472288 333922
rect 502688 334350 503008 334384
rect 502688 334294 502758 334350
rect 502814 334294 502882 334350
rect 502938 334294 503008 334350
rect 502688 334226 503008 334294
rect 502688 334170 502758 334226
rect 502814 334170 502882 334226
rect 502938 334170 503008 334226
rect 502688 334102 503008 334170
rect 502688 334046 502758 334102
rect 502814 334046 502882 334102
rect 502938 334046 503008 334102
rect 502688 333978 503008 334046
rect 502688 333922 502758 333978
rect 502814 333922 502882 333978
rect 502938 333922 503008 333978
rect 502688 333888 503008 333922
rect 533408 334350 533728 334384
rect 533408 334294 533478 334350
rect 533534 334294 533602 334350
rect 533658 334294 533728 334350
rect 533408 334226 533728 334294
rect 533408 334170 533478 334226
rect 533534 334170 533602 334226
rect 533658 334170 533728 334226
rect 533408 334102 533728 334170
rect 533408 334046 533478 334102
rect 533534 334046 533602 334102
rect 533658 334046 533728 334102
rect 533408 333978 533728 334046
rect 533408 333922 533478 333978
rect 533534 333922 533602 333978
rect 533658 333922 533728 333978
rect 533408 333888 533728 333922
rect 364448 328350 364768 328384
rect 364448 328294 364518 328350
rect 364574 328294 364642 328350
rect 364698 328294 364768 328350
rect 364448 328226 364768 328294
rect 364448 328170 364518 328226
rect 364574 328170 364642 328226
rect 364698 328170 364768 328226
rect 364448 328102 364768 328170
rect 364448 328046 364518 328102
rect 364574 328046 364642 328102
rect 364698 328046 364768 328102
rect 364448 327978 364768 328046
rect 364448 327922 364518 327978
rect 364574 327922 364642 327978
rect 364698 327922 364768 327978
rect 364448 327888 364768 327922
rect 395168 328350 395488 328384
rect 395168 328294 395238 328350
rect 395294 328294 395362 328350
rect 395418 328294 395488 328350
rect 395168 328226 395488 328294
rect 395168 328170 395238 328226
rect 395294 328170 395362 328226
rect 395418 328170 395488 328226
rect 395168 328102 395488 328170
rect 395168 328046 395238 328102
rect 395294 328046 395362 328102
rect 395418 328046 395488 328102
rect 395168 327978 395488 328046
rect 395168 327922 395238 327978
rect 395294 327922 395362 327978
rect 395418 327922 395488 327978
rect 395168 327888 395488 327922
rect 425888 328350 426208 328384
rect 425888 328294 425958 328350
rect 426014 328294 426082 328350
rect 426138 328294 426208 328350
rect 425888 328226 426208 328294
rect 425888 328170 425958 328226
rect 426014 328170 426082 328226
rect 426138 328170 426208 328226
rect 425888 328102 426208 328170
rect 425888 328046 425958 328102
rect 426014 328046 426082 328102
rect 426138 328046 426208 328102
rect 425888 327978 426208 328046
rect 425888 327922 425958 327978
rect 426014 327922 426082 327978
rect 426138 327922 426208 327978
rect 425888 327888 426208 327922
rect 456608 328350 456928 328384
rect 456608 328294 456678 328350
rect 456734 328294 456802 328350
rect 456858 328294 456928 328350
rect 456608 328226 456928 328294
rect 456608 328170 456678 328226
rect 456734 328170 456802 328226
rect 456858 328170 456928 328226
rect 456608 328102 456928 328170
rect 456608 328046 456678 328102
rect 456734 328046 456802 328102
rect 456858 328046 456928 328102
rect 456608 327978 456928 328046
rect 456608 327922 456678 327978
rect 456734 327922 456802 327978
rect 456858 327922 456928 327978
rect 456608 327888 456928 327922
rect 487328 328350 487648 328384
rect 487328 328294 487398 328350
rect 487454 328294 487522 328350
rect 487578 328294 487648 328350
rect 487328 328226 487648 328294
rect 487328 328170 487398 328226
rect 487454 328170 487522 328226
rect 487578 328170 487648 328226
rect 487328 328102 487648 328170
rect 487328 328046 487398 328102
rect 487454 328046 487522 328102
rect 487578 328046 487648 328102
rect 487328 327978 487648 328046
rect 487328 327922 487398 327978
rect 487454 327922 487522 327978
rect 487578 327922 487648 327978
rect 487328 327888 487648 327922
rect 518048 328350 518368 328384
rect 518048 328294 518118 328350
rect 518174 328294 518242 328350
rect 518298 328294 518368 328350
rect 518048 328226 518368 328294
rect 518048 328170 518118 328226
rect 518174 328170 518242 328226
rect 518298 328170 518368 328226
rect 518048 328102 518368 328170
rect 518048 328046 518118 328102
rect 518174 328046 518242 328102
rect 518298 328046 518368 328102
rect 518048 327978 518368 328046
rect 518048 327922 518118 327978
rect 518174 327922 518242 327978
rect 518298 327922 518368 327978
rect 518048 327888 518368 327922
rect 548768 328350 549088 328384
rect 548768 328294 548838 328350
rect 548894 328294 548962 328350
rect 549018 328294 549088 328350
rect 548768 328226 549088 328294
rect 548768 328170 548838 328226
rect 548894 328170 548962 328226
rect 549018 328170 549088 328226
rect 548768 328102 549088 328170
rect 548768 328046 548838 328102
rect 548894 328046 548962 328102
rect 549018 328046 549088 328102
rect 548768 327978 549088 328046
rect 548768 327922 548838 327978
rect 548894 327922 548962 327978
rect 549018 327922 549088 327978
rect 548768 327888 549088 327922
rect 360108 319788 360164 319798
rect 359884 317604 359940 317614
rect 360108 317548 360164 319732
rect 359884 308638 359940 317548
rect 359996 317492 360164 317548
rect 359996 308998 360052 317492
rect 379808 316350 380128 316384
rect 379808 316294 379878 316350
rect 379934 316294 380002 316350
rect 380058 316294 380128 316350
rect 379808 316226 380128 316294
rect 379808 316170 379878 316226
rect 379934 316170 380002 316226
rect 380058 316170 380128 316226
rect 379808 316102 380128 316170
rect 379808 316046 379878 316102
rect 379934 316046 380002 316102
rect 380058 316046 380128 316102
rect 379808 315978 380128 316046
rect 379808 315922 379878 315978
rect 379934 315922 380002 315978
rect 380058 315922 380128 315978
rect 379808 315888 380128 315922
rect 410528 316350 410848 316384
rect 410528 316294 410598 316350
rect 410654 316294 410722 316350
rect 410778 316294 410848 316350
rect 410528 316226 410848 316294
rect 410528 316170 410598 316226
rect 410654 316170 410722 316226
rect 410778 316170 410848 316226
rect 410528 316102 410848 316170
rect 410528 316046 410598 316102
rect 410654 316046 410722 316102
rect 410778 316046 410848 316102
rect 410528 315978 410848 316046
rect 410528 315922 410598 315978
rect 410654 315922 410722 315978
rect 410778 315922 410848 315978
rect 410528 315888 410848 315922
rect 441248 316350 441568 316384
rect 441248 316294 441318 316350
rect 441374 316294 441442 316350
rect 441498 316294 441568 316350
rect 441248 316226 441568 316294
rect 441248 316170 441318 316226
rect 441374 316170 441442 316226
rect 441498 316170 441568 316226
rect 441248 316102 441568 316170
rect 441248 316046 441318 316102
rect 441374 316046 441442 316102
rect 441498 316046 441568 316102
rect 441248 315978 441568 316046
rect 441248 315922 441318 315978
rect 441374 315922 441442 315978
rect 441498 315922 441568 315978
rect 441248 315888 441568 315922
rect 471968 316350 472288 316384
rect 471968 316294 472038 316350
rect 472094 316294 472162 316350
rect 472218 316294 472288 316350
rect 471968 316226 472288 316294
rect 471968 316170 472038 316226
rect 472094 316170 472162 316226
rect 472218 316170 472288 316226
rect 471968 316102 472288 316170
rect 471968 316046 472038 316102
rect 472094 316046 472162 316102
rect 472218 316046 472288 316102
rect 471968 315978 472288 316046
rect 471968 315922 472038 315978
rect 472094 315922 472162 315978
rect 472218 315922 472288 315978
rect 471968 315888 472288 315922
rect 502688 316350 503008 316384
rect 502688 316294 502758 316350
rect 502814 316294 502882 316350
rect 502938 316294 503008 316350
rect 502688 316226 503008 316294
rect 502688 316170 502758 316226
rect 502814 316170 502882 316226
rect 502938 316170 503008 316226
rect 502688 316102 503008 316170
rect 502688 316046 502758 316102
rect 502814 316046 502882 316102
rect 502938 316046 503008 316102
rect 502688 315978 503008 316046
rect 502688 315922 502758 315978
rect 502814 315922 502882 315978
rect 502938 315922 503008 315978
rect 502688 315888 503008 315922
rect 533408 316350 533728 316384
rect 533408 316294 533478 316350
rect 533534 316294 533602 316350
rect 533658 316294 533728 316350
rect 533408 316226 533728 316294
rect 533408 316170 533478 316226
rect 533534 316170 533602 316226
rect 533658 316170 533728 316226
rect 533408 316102 533728 316170
rect 533408 316046 533478 316102
rect 533534 316046 533602 316102
rect 533658 316046 533728 316102
rect 533408 315978 533728 316046
rect 533408 315922 533478 315978
rect 533534 315922 533602 315978
rect 533658 315922 533728 315978
rect 533408 315888 533728 315922
rect 364448 310350 364768 310384
rect 364448 310294 364518 310350
rect 364574 310294 364642 310350
rect 364698 310294 364768 310350
rect 364448 310226 364768 310294
rect 364448 310170 364518 310226
rect 364574 310170 364642 310226
rect 364698 310170 364768 310226
rect 364448 310102 364768 310170
rect 364448 310046 364518 310102
rect 364574 310046 364642 310102
rect 364698 310046 364768 310102
rect 364448 309978 364768 310046
rect 364448 309922 364518 309978
rect 364574 309922 364642 309978
rect 364698 309922 364768 309978
rect 364448 309888 364768 309922
rect 395168 310350 395488 310384
rect 395168 310294 395238 310350
rect 395294 310294 395362 310350
rect 395418 310294 395488 310350
rect 395168 310226 395488 310294
rect 395168 310170 395238 310226
rect 395294 310170 395362 310226
rect 395418 310170 395488 310226
rect 395168 310102 395488 310170
rect 395168 310046 395238 310102
rect 395294 310046 395362 310102
rect 395418 310046 395488 310102
rect 395168 309978 395488 310046
rect 395168 309922 395238 309978
rect 395294 309922 395362 309978
rect 395418 309922 395488 309978
rect 395168 309888 395488 309922
rect 425888 310350 426208 310384
rect 425888 310294 425958 310350
rect 426014 310294 426082 310350
rect 426138 310294 426208 310350
rect 425888 310226 426208 310294
rect 425888 310170 425958 310226
rect 426014 310170 426082 310226
rect 426138 310170 426208 310226
rect 425888 310102 426208 310170
rect 425888 310046 425958 310102
rect 426014 310046 426082 310102
rect 426138 310046 426208 310102
rect 425888 309978 426208 310046
rect 425888 309922 425958 309978
rect 426014 309922 426082 309978
rect 426138 309922 426208 309978
rect 425888 309888 426208 309922
rect 456608 310350 456928 310384
rect 456608 310294 456678 310350
rect 456734 310294 456802 310350
rect 456858 310294 456928 310350
rect 456608 310226 456928 310294
rect 456608 310170 456678 310226
rect 456734 310170 456802 310226
rect 456858 310170 456928 310226
rect 456608 310102 456928 310170
rect 456608 310046 456678 310102
rect 456734 310046 456802 310102
rect 456858 310046 456928 310102
rect 456608 309978 456928 310046
rect 456608 309922 456678 309978
rect 456734 309922 456802 309978
rect 456858 309922 456928 309978
rect 456608 309888 456928 309922
rect 487328 310350 487648 310384
rect 487328 310294 487398 310350
rect 487454 310294 487522 310350
rect 487578 310294 487648 310350
rect 487328 310226 487648 310294
rect 487328 310170 487398 310226
rect 487454 310170 487522 310226
rect 487578 310170 487648 310226
rect 487328 310102 487648 310170
rect 487328 310046 487398 310102
rect 487454 310046 487522 310102
rect 487578 310046 487648 310102
rect 487328 309978 487648 310046
rect 487328 309922 487398 309978
rect 487454 309922 487522 309978
rect 487578 309922 487648 309978
rect 487328 309888 487648 309922
rect 518048 310350 518368 310384
rect 518048 310294 518118 310350
rect 518174 310294 518242 310350
rect 518298 310294 518368 310350
rect 518048 310226 518368 310294
rect 518048 310170 518118 310226
rect 518174 310170 518242 310226
rect 518298 310170 518368 310226
rect 518048 310102 518368 310170
rect 518048 310046 518118 310102
rect 518174 310046 518242 310102
rect 518298 310046 518368 310102
rect 518048 309978 518368 310046
rect 518048 309922 518118 309978
rect 518174 309922 518242 309978
rect 518298 309922 518368 309978
rect 518048 309888 518368 309922
rect 548768 310350 549088 310384
rect 548768 310294 548838 310350
rect 548894 310294 548962 310350
rect 549018 310294 549088 310350
rect 548768 310226 549088 310294
rect 548768 310170 548838 310226
rect 548894 310170 548962 310226
rect 549018 310170 549088 310226
rect 548768 310102 549088 310170
rect 548768 310046 548838 310102
rect 548894 310046 548962 310102
rect 549018 310046 549088 310102
rect 548768 309978 549088 310046
rect 548768 309922 548838 309978
rect 548894 309922 548962 309978
rect 549018 309922 549088 309978
rect 548768 309888 549088 309922
rect 359996 308942 360164 308998
rect 359884 308572 359940 308582
rect 360108 308638 360164 308942
rect 360108 308572 360164 308582
rect 360108 308458 360164 308468
rect 360108 305788 360164 308402
rect 360332 308278 360388 308288
rect 360108 305732 360276 305788
rect 360220 298918 360276 305732
rect 360108 298862 360276 298918
rect 359772 240146 359828 240156
rect 359884 296100 359940 296110
rect 359660 235956 359716 235966
rect 359660 235852 359716 235862
rect 359660 216132 359716 216142
rect 359660 165508 359716 216076
rect 359884 215038 359940 296044
rect 359996 287398 360052 287408
rect 359996 235918 360052 287342
rect 359996 235852 360052 235862
rect 359884 214982 360052 215038
rect 359996 211708 360052 214982
rect 359884 211652 360052 211708
rect 359884 209300 359940 211652
rect 359884 209234 359940 209244
rect 359884 206052 359940 206062
rect 360108 206038 360164 298862
rect 359940 205996 360164 206038
rect 359884 205982 360164 205996
rect 359884 205828 359940 205838
rect 359772 196196 359828 196206
rect 359772 191818 359828 196140
rect 359772 191752 359828 191762
rect 359772 191660 359828 191670
rect 359772 186058 359828 191604
rect 359884 186228 359940 205772
rect 359884 186162 359940 186172
rect 359772 185992 359828 186002
rect 359884 186004 359940 186014
rect 359772 185698 359828 185708
rect 359772 181412 359828 185642
rect 359772 181346 359828 181356
rect 359660 165442 359716 165452
rect 359772 178052 359828 178062
rect 359548 116946 359604 116956
rect 358652 52658 358708 52668
rect 355292 48066 355348 48076
rect 353612 45154 353668 45164
rect 359772 45108 359828 177996
rect 359884 115858 359940 185948
rect 359996 185878 360052 185888
rect 359996 118804 360052 185822
rect 360108 157078 360164 205982
rect 360220 296758 360276 296768
rect 360220 185698 360276 296702
rect 360220 185632 360276 185642
rect 360332 172228 360388 308222
rect 379808 298350 380128 298384
rect 379808 298294 379878 298350
rect 379934 298294 380002 298350
rect 380058 298294 380128 298350
rect 379808 298226 380128 298294
rect 379808 298170 379878 298226
rect 379934 298170 380002 298226
rect 380058 298170 380128 298226
rect 379808 298102 380128 298170
rect 379808 298046 379878 298102
rect 379934 298046 380002 298102
rect 380058 298046 380128 298102
rect 379808 297978 380128 298046
rect 379808 297922 379878 297978
rect 379934 297922 380002 297978
rect 380058 297922 380128 297978
rect 379808 297888 380128 297922
rect 410528 298350 410848 298384
rect 410528 298294 410598 298350
rect 410654 298294 410722 298350
rect 410778 298294 410848 298350
rect 410528 298226 410848 298294
rect 410528 298170 410598 298226
rect 410654 298170 410722 298226
rect 410778 298170 410848 298226
rect 410528 298102 410848 298170
rect 410528 298046 410598 298102
rect 410654 298046 410722 298102
rect 410778 298046 410848 298102
rect 410528 297978 410848 298046
rect 410528 297922 410598 297978
rect 410654 297922 410722 297978
rect 410778 297922 410848 297978
rect 410528 297888 410848 297922
rect 441248 298350 441568 298384
rect 441248 298294 441318 298350
rect 441374 298294 441442 298350
rect 441498 298294 441568 298350
rect 441248 298226 441568 298294
rect 441248 298170 441318 298226
rect 441374 298170 441442 298226
rect 441498 298170 441568 298226
rect 441248 298102 441568 298170
rect 441248 298046 441318 298102
rect 441374 298046 441442 298102
rect 441498 298046 441568 298102
rect 441248 297978 441568 298046
rect 441248 297922 441318 297978
rect 441374 297922 441442 297978
rect 441498 297922 441568 297978
rect 441248 297888 441568 297922
rect 471968 298350 472288 298384
rect 471968 298294 472038 298350
rect 472094 298294 472162 298350
rect 472218 298294 472288 298350
rect 471968 298226 472288 298294
rect 471968 298170 472038 298226
rect 472094 298170 472162 298226
rect 472218 298170 472288 298226
rect 471968 298102 472288 298170
rect 471968 298046 472038 298102
rect 472094 298046 472162 298102
rect 472218 298046 472288 298102
rect 471968 297978 472288 298046
rect 471968 297922 472038 297978
rect 472094 297922 472162 297978
rect 472218 297922 472288 297978
rect 471968 297888 472288 297922
rect 502688 298350 503008 298384
rect 502688 298294 502758 298350
rect 502814 298294 502882 298350
rect 502938 298294 503008 298350
rect 502688 298226 503008 298294
rect 502688 298170 502758 298226
rect 502814 298170 502882 298226
rect 502938 298170 503008 298226
rect 502688 298102 503008 298170
rect 502688 298046 502758 298102
rect 502814 298046 502882 298102
rect 502938 298046 503008 298102
rect 502688 297978 503008 298046
rect 502688 297922 502758 297978
rect 502814 297922 502882 297978
rect 502938 297922 503008 297978
rect 502688 297888 503008 297922
rect 533408 298350 533728 298384
rect 533408 298294 533478 298350
rect 533534 298294 533602 298350
rect 533658 298294 533728 298350
rect 533408 298226 533728 298294
rect 533408 298170 533478 298226
rect 533534 298170 533602 298226
rect 533658 298170 533728 298226
rect 533408 298102 533728 298170
rect 533408 298046 533478 298102
rect 533534 298046 533602 298102
rect 533658 298046 533728 298102
rect 533408 297978 533728 298046
rect 533408 297922 533478 297978
rect 533534 297922 533602 297978
rect 533658 297922 533728 297978
rect 533408 297888 533728 297922
rect 362012 292618 362068 292628
rect 360332 172162 360388 172172
rect 360444 255718 360500 255728
rect 360108 157012 360164 157022
rect 359996 118738 360052 118748
rect 360444 117124 360500 255662
rect 361788 235918 361844 235928
rect 360556 191818 360612 191828
rect 360556 172116 360612 191762
rect 361228 184618 361284 184628
rect 361116 184562 361228 184618
rect 361116 182098 361172 184562
rect 361228 184552 361284 184562
rect 361788 183876 361844 235862
rect 361900 193978 361956 193988
rect 361900 184618 361956 193922
rect 361900 184552 361956 184562
rect 361340 183820 361844 183876
rect 361340 182638 361396 183820
rect 361340 182582 361844 182638
rect 361116 182042 361732 182098
rect 361564 181018 361620 181028
rect 361452 176338 361508 176348
rect 361452 175364 361508 176282
rect 361452 175298 361508 175308
rect 360556 172050 360612 172060
rect 361564 168028 361620 180962
rect 361676 174580 361732 182042
rect 361676 174514 361732 174524
rect 361564 167972 361732 168028
rect 361676 162596 361732 167972
rect 361676 162530 361732 162540
rect 361788 118580 361844 182582
rect 362012 118692 362068 292562
rect 364448 292350 364768 292384
rect 364448 292294 364518 292350
rect 364574 292294 364642 292350
rect 364698 292294 364768 292350
rect 364448 292226 364768 292294
rect 364448 292170 364518 292226
rect 364574 292170 364642 292226
rect 364698 292170 364768 292226
rect 364448 292102 364768 292170
rect 364448 292046 364518 292102
rect 364574 292046 364642 292102
rect 364698 292046 364768 292102
rect 364448 291978 364768 292046
rect 364448 291922 364518 291978
rect 364574 291922 364642 291978
rect 364698 291922 364768 291978
rect 364448 291888 364768 291922
rect 395168 292350 395488 292384
rect 395168 292294 395238 292350
rect 395294 292294 395362 292350
rect 395418 292294 395488 292350
rect 395168 292226 395488 292294
rect 395168 292170 395238 292226
rect 395294 292170 395362 292226
rect 395418 292170 395488 292226
rect 395168 292102 395488 292170
rect 395168 292046 395238 292102
rect 395294 292046 395362 292102
rect 395418 292046 395488 292102
rect 395168 291978 395488 292046
rect 395168 291922 395238 291978
rect 395294 291922 395362 291978
rect 395418 291922 395488 291978
rect 395168 291888 395488 291922
rect 425888 292350 426208 292384
rect 425888 292294 425958 292350
rect 426014 292294 426082 292350
rect 426138 292294 426208 292350
rect 425888 292226 426208 292294
rect 425888 292170 425958 292226
rect 426014 292170 426082 292226
rect 426138 292170 426208 292226
rect 425888 292102 426208 292170
rect 425888 292046 425958 292102
rect 426014 292046 426082 292102
rect 426138 292046 426208 292102
rect 425888 291978 426208 292046
rect 425888 291922 425958 291978
rect 426014 291922 426082 291978
rect 426138 291922 426208 291978
rect 425888 291888 426208 291922
rect 456608 292350 456928 292384
rect 456608 292294 456678 292350
rect 456734 292294 456802 292350
rect 456858 292294 456928 292350
rect 456608 292226 456928 292294
rect 456608 292170 456678 292226
rect 456734 292170 456802 292226
rect 456858 292170 456928 292226
rect 456608 292102 456928 292170
rect 456608 292046 456678 292102
rect 456734 292046 456802 292102
rect 456858 292046 456928 292102
rect 456608 291978 456928 292046
rect 456608 291922 456678 291978
rect 456734 291922 456802 291978
rect 456858 291922 456928 291978
rect 456608 291888 456928 291922
rect 487328 292350 487648 292384
rect 487328 292294 487398 292350
rect 487454 292294 487522 292350
rect 487578 292294 487648 292350
rect 487328 292226 487648 292294
rect 487328 292170 487398 292226
rect 487454 292170 487522 292226
rect 487578 292170 487648 292226
rect 487328 292102 487648 292170
rect 487328 292046 487398 292102
rect 487454 292046 487522 292102
rect 487578 292046 487648 292102
rect 487328 291978 487648 292046
rect 487328 291922 487398 291978
rect 487454 291922 487522 291978
rect 487578 291922 487648 291978
rect 487328 291888 487648 291922
rect 518048 292350 518368 292384
rect 518048 292294 518118 292350
rect 518174 292294 518242 292350
rect 518298 292294 518368 292350
rect 518048 292226 518368 292294
rect 518048 292170 518118 292226
rect 518174 292170 518242 292226
rect 518298 292170 518368 292226
rect 518048 292102 518368 292170
rect 518048 292046 518118 292102
rect 518174 292046 518242 292102
rect 518298 292046 518368 292102
rect 518048 291978 518368 292046
rect 518048 291922 518118 291978
rect 518174 291922 518242 291978
rect 518298 291922 518368 291978
rect 518048 291888 518368 291922
rect 548768 292350 549088 292384
rect 548768 292294 548838 292350
rect 548894 292294 548962 292350
rect 549018 292294 549088 292350
rect 548768 292226 549088 292294
rect 548768 292170 548838 292226
rect 548894 292170 548962 292226
rect 549018 292170 549088 292226
rect 548768 292102 549088 292170
rect 548768 292046 548838 292102
rect 548894 292046 548962 292102
rect 549018 292046 549088 292102
rect 548768 291978 549088 292046
rect 548768 291922 548838 291978
rect 548894 291922 548962 291978
rect 549018 291922 549088 291978
rect 548768 291888 549088 291922
rect 379808 280350 380128 280384
rect 379808 280294 379878 280350
rect 379934 280294 380002 280350
rect 380058 280294 380128 280350
rect 379808 280226 380128 280294
rect 379808 280170 379878 280226
rect 379934 280170 380002 280226
rect 380058 280170 380128 280226
rect 379808 280102 380128 280170
rect 379808 280046 379878 280102
rect 379934 280046 380002 280102
rect 380058 280046 380128 280102
rect 379808 279978 380128 280046
rect 379808 279922 379878 279978
rect 379934 279922 380002 279978
rect 380058 279922 380128 279978
rect 379808 279888 380128 279922
rect 410528 280350 410848 280384
rect 410528 280294 410598 280350
rect 410654 280294 410722 280350
rect 410778 280294 410848 280350
rect 410528 280226 410848 280294
rect 410528 280170 410598 280226
rect 410654 280170 410722 280226
rect 410778 280170 410848 280226
rect 410528 280102 410848 280170
rect 410528 280046 410598 280102
rect 410654 280046 410722 280102
rect 410778 280046 410848 280102
rect 410528 279978 410848 280046
rect 410528 279922 410598 279978
rect 410654 279922 410722 279978
rect 410778 279922 410848 279978
rect 410528 279888 410848 279922
rect 441248 280350 441568 280384
rect 441248 280294 441318 280350
rect 441374 280294 441442 280350
rect 441498 280294 441568 280350
rect 441248 280226 441568 280294
rect 441248 280170 441318 280226
rect 441374 280170 441442 280226
rect 441498 280170 441568 280226
rect 441248 280102 441568 280170
rect 441248 280046 441318 280102
rect 441374 280046 441442 280102
rect 441498 280046 441568 280102
rect 441248 279978 441568 280046
rect 441248 279922 441318 279978
rect 441374 279922 441442 279978
rect 441498 279922 441568 279978
rect 441248 279888 441568 279922
rect 471968 280350 472288 280384
rect 471968 280294 472038 280350
rect 472094 280294 472162 280350
rect 472218 280294 472288 280350
rect 471968 280226 472288 280294
rect 471968 280170 472038 280226
rect 472094 280170 472162 280226
rect 472218 280170 472288 280226
rect 471968 280102 472288 280170
rect 471968 280046 472038 280102
rect 472094 280046 472162 280102
rect 472218 280046 472288 280102
rect 471968 279978 472288 280046
rect 471968 279922 472038 279978
rect 472094 279922 472162 279978
rect 472218 279922 472288 279978
rect 471968 279888 472288 279922
rect 502688 280350 503008 280384
rect 502688 280294 502758 280350
rect 502814 280294 502882 280350
rect 502938 280294 503008 280350
rect 502688 280226 503008 280294
rect 502688 280170 502758 280226
rect 502814 280170 502882 280226
rect 502938 280170 503008 280226
rect 502688 280102 503008 280170
rect 502688 280046 502758 280102
rect 502814 280046 502882 280102
rect 502938 280046 503008 280102
rect 502688 279978 503008 280046
rect 502688 279922 502758 279978
rect 502814 279922 502882 279978
rect 502938 279922 503008 279978
rect 502688 279888 503008 279922
rect 533408 280350 533728 280384
rect 533408 280294 533478 280350
rect 533534 280294 533602 280350
rect 533658 280294 533728 280350
rect 533408 280226 533728 280294
rect 533408 280170 533478 280226
rect 533534 280170 533602 280226
rect 533658 280170 533728 280226
rect 533408 280102 533728 280170
rect 533408 280046 533478 280102
rect 533534 280046 533602 280102
rect 533658 280046 533728 280102
rect 533408 279978 533728 280046
rect 533408 279922 533478 279978
rect 533534 279922 533602 279978
rect 533658 279922 533728 279978
rect 533408 279888 533728 279922
rect 364448 274350 364768 274384
rect 364448 274294 364518 274350
rect 364574 274294 364642 274350
rect 364698 274294 364768 274350
rect 364448 274226 364768 274294
rect 364448 274170 364518 274226
rect 364574 274170 364642 274226
rect 364698 274170 364768 274226
rect 364448 274102 364768 274170
rect 364448 274046 364518 274102
rect 364574 274046 364642 274102
rect 364698 274046 364768 274102
rect 364448 273978 364768 274046
rect 364448 273922 364518 273978
rect 364574 273922 364642 273978
rect 364698 273922 364768 273978
rect 364448 273888 364768 273922
rect 395168 274350 395488 274384
rect 395168 274294 395238 274350
rect 395294 274294 395362 274350
rect 395418 274294 395488 274350
rect 395168 274226 395488 274294
rect 395168 274170 395238 274226
rect 395294 274170 395362 274226
rect 395418 274170 395488 274226
rect 395168 274102 395488 274170
rect 395168 274046 395238 274102
rect 395294 274046 395362 274102
rect 395418 274046 395488 274102
rect 395168 273978 395488 274046
rect 395168 273922 395238 273978
rect 395294 273922 395362 273978
rect 395418 273922 395488 273978
rect 395168 273888 395488 273922
rect 425888 274350 426208 274384
rect 425888 274294 425958 274350
rect 426014 274294 426082 274350
rect 426138 274294 426208 274350
rect 425888 274226 426208 274294
rect 425888 274170 425958 274226
rect 426014 274170 426082 274226
rect 426138 274170 426208 274226
rect 425888 274102 426208 274170
rect 425888 274046 425958 274102
rect 426014 274046 426082 274102
rect 426138 274046 426208 274102
rect 425888 273978 426208 274046
rect 425888 273922 425958 273978
rect 426014 273922 426082 273978
rect 426138 273922 426208 273978
rect 425888 273888 426208 273922
rect 456608 274350 456928 274384
rect 456608 274294 456678 274350
rect 456734 274294 456802 274350
rect 456858 274294 456928 274350
rect 456608 274226 456928 274294
rect 456608 274170 456678 274226
rect 456734 274170 456802 274226
rect 456858 274170 456928 274226
rect 456608 274102 456928 274170
rect 456608 274046 456678 274102
rect 456734 274046 456802 274102
rect 456858 274046 456928 274102
rect 456608 273978 456928 274046
rect 456608 273922 456678 273978
rect 456734 273922 456802 273978
rect 456858 273922 456928 273978
rect 456608 273888 456928 273922
rect 487328 274350 487648 274384
rect 487328 274294 487398 274350
rect 487454 274294 487522 274350
rect 487578 274294 487648 274350
rect 487328 274226 487648 274294
rect 487328 274170 487398 274226
rect 487454 274170 487522 274226
rect 487578 274170 487648 274226
rect 487328 274102 487648 274170
rect 487328 274046 487398 274102
rect 487454 274046 487522 274102
rect 487578 274046 487648 274102
rect 487328 273978 487648 274046
rect 487328 273922 487398 273978
rect 487454 273922 487522 273978
rect 487578 273922 487648 273978
rect 487328 273888 487648 273922
rect 518048 274350 518368 274384
rect 518048 274294 518118 274350
rect 518174 274294 518242 274350
rect 518298 274294 518368 274350
rect 518048 274226 518368 274294
rect 518048 274170 518118 274226
rect 518174 274170 518242 274226
rect 518298 274170 518368 274226
rect 518048 274102 518368 274170
rect 518048 274046 518118 274102
rect 518174 274046 518242 274102
rect 518298 274046 518368 274102
rect 518048 273978 518368 274046
rect 518048 273922 518118 273978
rect 518174 273922 518242 273978
rect 518298 273922 518368 273978
rect 518048 273888 518368 273922
rect 548768 274350 549088 274384
rect 548768 274294 548838 274350
rect 548894 274294 548962 274350
rect 549018 274294 549088 274350
rect 548768 274226 549088 274294
rect 548768 274170 548838 274226
rect 548894 274170 548962 274226
rect 549018 274170 549088 274226
rect 548768 274102 549088 274170
rect 548768 274046 548838 274102
rect 548894 274046 548962 274102
rect 549018 274046 549088 274102
rect 548768 273978 549088 274046
rect 548768 273922 548838 273978
rect 548894 273922 548962 273978
rect 549018 273922 549088 273978
rect 548768 273888 549088 273922
rect 379808 262350 380128 262384
rect 379808 262294 379878 262350
rect 379934 262294 380002 262350
rect 380058 262294 380128 262350
rect 379808 262226 380128 262294
rect 379808 262170 379878 262226
rect 379934 262170 380002 262226
rect 380058 262170 380128 262226
rect 379808 262102 380128 262170
rect 379808 262046 379878 262102
rect 379934 262046 380002 262102
rect 380058 262046 380128 262102
rect 379808 261978 380128 262046
rect 379808 261922 379878 261978
rect 379934 261922 380002 261978
rect 380058 261922 380128 261978
rect 379808 261888 380128 261922
rect 410528 262350 410848 262384
rect 410528 262294 410598 262350
rect 410654 262294 410722 262350
rect 410778 262294 410848 262350
rect 410528 262226 410848 262294
rect 410528 262170 410598 262226
rect 410654 262170 410722 262226
rect 410778 262170 410848 262226
rect 410528 262102 410848 262170
rect 410528 262046 410598 262102
rect 410654 262046 410722 262102
rect 410778 262046 410848 262102
rect 410528 261978 410848 262046
rect 410528 261922 410598 261978
rect 410654 261922 410722 261978
rect 410778 261922 410848 261978
rect 410528 261888 410848 261922
rect 441248 262350 441568 262384
rect 441248 262294 441318 262350
rect 441374 262294 441442 262350
rect 441498 262294 441568 262350
rect 441248 262226 441568 262294
rect 441248 262170 441318 262226
rect 441374 262170 441442 262226
rect 441498 262170 441568 262226
rect 441248 262102 441568 262170
rect 441248 262046 441318 262102
rect 441374 262046 441442 262102
rect 441498 262046 441568 262102
rect 441248 261978 441568 262046
rect 441248 261922 441318 261978
rect 441374 261922 441442 261978
rect 441498 261922 441568 261978
rect 441248 261888 441568 261922
rect 471968 262350 472288 262384
rect 471968 262294 472038 262350
rect 472094 262294 472162 262350
rect 472218 262294 472288 262350
rect 471968 262226 472288 262294
rect 471968 262170 472038 262226
rect 472094 262170 472162 262226
rect 472218 262170 472288 262226
rect 471968 262102 472288 262170
rect 471968 262046 472038 262102
rect 472094 262046 472162 262102
rect 472218 262046 472288 262102
rect 471968 261978 472288 262046
rect 471968 261922 472038 261978
rect 472094 261922 472162 261978
rect 472218 261922 472288 261978
rect 471968 261888 472288 261922
rect 502688 262350 503008 262384
rect 502688 262294 502758 262350
rect 502814 262294 502882 262350
rect 502938 262294 503008 262350
rect 502688 262226 503008 262294
rect 502688 262170 502758 262226
rect 502814 262170 502882 262226
rect 502938 262170 503008 262226
rect 502688 262102 503008 262170
rect 502688 262046 502758 262102
rect 502814 262046 502882 262102
rect 502938 262046 503008 262102
rect 502688 261978 503008 262046
rect 502688 261922 502758 261978
rect 502814 261922 502882 261978
rect 502938 261922 503008 261978
rect 502688 261888 503008 261922
rect 533408 262350 533728 262384
rect 533408 262294 533478 262350
rect 533534 262294 533602 262350
rect 533658 262294 533728 262350
rect 533408 262226 533728 262294
rect 533408 262170 533478 262226
rect 533534 262170 533602 262226
rect 533658 262170 533728 262226
rect 533408 262102 533728 262170
rect 533408 262046 533478 262102
rect 533534 262046 533602 262102
rect 533658 262046 533728 262102
rect 533408 261978 533728 262046
rect 533408 261922 533478 261978
rect 533534 261922 533602 261978
rect 533658 261922 533728 261978
rect 533408 261888 533728 261922
rect 364448 256350 364768 256384
rect 364448 256294 364518 256350
rect 364574 256294 364642 256350
rect 364698 256294 364768 256350
rect 364448 256226 364768 256294
rect 364448 256170 364518 256226
rect 364574 256170 364642 256226
rect 364698 256170 364768 256226
rect 364448 256102 364768 256170
rect 364448 256046 364518 256102
rect 364574 256046 364642 256102
rect 364698 256046 364768 256102
rect 364448 255978 364768 256046
rect 364448 255922 364518 255978
rect 364574 255922 364642 255978
rect 364698 255922 364768 255978
rect 364448 255888 364768 255922
rect 395168 256350 395488 256384
rect 395168 256294 395238 256350
rect 395294 256294 395362 256350
rect 395418 256294 395488 256350
rect 395168 256226 395488 256294
rect 395168 256170 395238 256226
rect 395294 256170 395362 256226
rect 395418 256170 395488 256226
rect 395168 256102 395488 256170
rect 395168 256046 395238 256102
rect 395294 256046 395362 256102
rect 395418 256046 395488 256102
rect 395168 255978 395488 256046
rect 395168 255922 395238 255978
rect 395294 255922 395362 255978
rect 395418 255922 395488 255978
rect 395168 255888 395488 255922
rect 425888 256350 426208 256384
rect 425888 256294 425958 256350
rect 426014 256294 426082 256350
rect 426138 256294 426208 256350
rect 425888 256226 426208 256294
rect 425888 256170 425958 256226
rect 426014 256170 426082 256226
rect 426138 256170 426208 256226
rect 425888 256102 426208 256170
rect 425888 256046 425958 256102
rect 426014 256046 426082 256102
rect 426138 256046 426208 256102
rect 425888 255978 426208 256046
rect 425888 255922 425958 255978
rect 426014 255922 426082 255978
rect 426138 255922 426208 255978
rect 425888 255888 426208 255922
rect 456608 256350 456928 256384
rect 456608 256294 456678 256350
rect 456734 256294 456802 256350
rect 456858 256294 456928 256350
rect 456608 256226 456928 256294
rect 456608 256170 456678 256226
rect 456734 256170 456802 256226
rect 456858 256170 456928 256226
rect 456608 256102 456928 256170
rect 456608 256046 456678 256102
rect 456734 256046 456802 256102
rect 456858 256046 456928 256102
rect 456608 255978 456928 256046
rect 456608 255922 456678 255978
rect 456734 255922 456802 255978
rect 456858 255922 456928 255978
rect 456608 255888 456928 255922
rect 487328 256350 487648 256384
rect 487328 256294 487398 256350
rect 487454 256294 487522 256350
rect 487578 256294 487648 256350
rect 487328 256226 487648 256294
rect 487328 256170 487398 256226
rect 487454 256170 487522 256226
rect 487578 256170 487648 256226
rect 487328 256102 487648 256170
rect 487328 256046 487398 256102
rect 487454 256046 487522 256102
rect 487578 256046 487648 256102
rect 487328 255978 487648 256046
rect 487328 255922 487398 255978
rect 487454 255922 487522 255978
rect 487578 255922 487648 255978
rect 487328 255888 487648 255922
rect 518048 256350 518368 256384
rect 518048 256294 518118 256350
rect 518174 256294 518242 256350
rect 518298 256294 518368 256350
rect 518048 256226 518368 256294
rect 518048 256170 518118 256226
rect 518174 256170 518242 256226
rect 518298 256170 518368 256226
rect 518048 256102 518368 256170
rect 518048 256046 518118 256102
rect 518174 256046 518242 256102
rect 518298 256046 518368 256102
rect 518048 255978 518368 256046
rect 518048 255922 518118 255978
rect 518174 255922 518242 255978
rect 518298 255922 518368 255978
rect 518048 255888 518368 255922
rect 548768 256350 549088 256384
rect 548768 256294 548838 256350
rect 548894 256294 548962 256350
rect 549018 256294 549088 256350
rect 548768 256226 549088 256294
rect 548768 256170 548838 256226
rect 548894 256170 548962 256226
rect 549018 256170 549088 256226
rect 548768 256102 549088 256170
rect 548768 256046 548838 256102
rect 548894 256046 548962 256102
rect 549018 256046 549088 256102
rect 548768 255978 549088 256046
rect 548768 255922 548838 255978
rect 548894 255922 548962 255978
rect 549018 255922 549088 255978
rect 548768 255888 549088 255922
rect 379808 244350 380128 244384
rect 379808 244294 379878 244350
rect 379934 244294 380002 244350
rect 380058 244294 380128 244350
rect 379808 244226 380128 244294
rect 379808 244170 379878 244226
rect 379934 244170 380002 244226
rect 380058 244170 380128 244226
rect 379808 244102 380128 244170
rect 379808 244046 379878 244102
rect 379934 244046 380002 244102
rect 380058 244046 380128 244102
rect 379808 243978 380128 244046
rect 379808 243922 379878 243978
rect 379934 243922 380002 243978
rect 380058 243922 380128 243978
rect 379808 243888 380128 243922
rect 410528 244350 410848 244384
rect 410528 244294 410598 244350
rect 410654 244294 410722 244350
rect 410778 244294 410848 244350
rect 410528 244226 410848 244294
rect 410528 244170 410598 244226
rect 410654 244170 410722 244226
rect 410778 244170 410848 244226
rect 410528 244102 410848 244170
rect 410528 244046 410598 244102
rect 410654 244046 410722 244102
rect 410778 244046 410848 244102
rect 410528 243978 410848 244046
rect 410528 243922 410598 243978
rect 410654 243922 410722 243978
rect 410778 243922 410848 243978
rect 410528 243888 410848 243922
rect 441248 244350 441568 244384
rect 441248 244294 441318 244350
rect 441374 244294 441442 244350
rect 441498 244294 441568 244350
rect 441248 244226 441568 244294
rect 441248 244170 441318 244226
rect 441374 244170 441442 244226
rect 441498 244170 441568 244226
rect 441248 244102 441568 244170
rect 441248 244046 441318 244102
rect 441374 244046 441442 244102
rect 441498 244046 441568 244102
rect 441248 243978 441568 244046
rect 441248 243922 441318 243978
rect 441374 243922 441442 243978
rect 441498 243922 441568 243978
rect 441248 243888 441568 243922
rect 471968 244350 472288 244384
rect 471968 244294 472038 244350
rect 472094 244294 472162 244350
rect 472218 244294 472288 244350
rect 471968 244226 472288 244294
rect 471968 244170 472038 244226
rect 472094 244170 472162 244226
rect 472218 244170 472288 244226
rect 471968 244102 472288 244170
rect 471968 244046 472038 244102
rect 472094 244046 472162 244102
rect 472218 244046 472288 244102
rect 471968 243978 472288 244046
rect 471968 243922 472038 243978
rect 472094 243922 472162 243978
rect 472218 243922 472288 243978
rect 471968 243888 472288 243922
rect 502688 244350 503008 244384
rect 502688 244294 502758 244350
rect 502814 244294 502882 244350
rect 502938 244294 503008 244350
rect 502688 244226 503008 244294
rect 502688 244170 502758 244226
rect 502814 244170 502882 244226
rect 502938 244170 503008 244226
rect 502688 244102 503008 244170
rect 502688 244046 502758 244102
rect 502814 244046 502882 244102
rect 502938 244046 503008 244102
rect 502688 243978 503008 244046
rect 502688 243922 502758 243978
rect 502814 243922 502882 243978
rect 502938 243922 503008 243978
rect 502688 243888 503008 243922
rect 533408 244350 533728 244384
rect 533408 244294 533478 244350
rect 533534 244294 533602 244350
rect 533658 244294 533728 244350
rect 533408 244226 533728 244294
rect 533408 244170 533478 244226
rect 533534 244170 533602 244226
rect 533658 244170 533728 244226
rect 533408 244102 533728 244170
rect 533408 244046 533478 244102
rect 533534 244046 533602 244102
rect 533658 244046 533728 244102
rect 533408 243978 533728 244046
rect 533408 243922 533478 243978
rect 533534 243922 533602 243978
rect 533658 243922 533728 243978
rect 533408 243888 533728 243922
rect 364448 238350 364768 238384
rect 364448 238294 364518 238350
rect 364574 238294 364642 238350
rect 364698 238294 364768 238350
rect 364448 238226 364768 238294
rect 364448 238170 364518 238226
rect 364574 238170 364642 238226
rect 364698 238170 364768 238226
rect 364448 238102 364768 238170
rect 364448 238046 364518 238102
rect 364574 238046 364642 238102
rect 364698 238046 364768 238102
rect 364448 237978 364768 238046
rect 364448 237922 364518 237978
rect 364574 237922 364642 237978
rect 364698 237922 364768 237978
rect 364448 237888 364768 237922
rect 395168 238350 395488 238384
rect 395168 238294 395238 238350
rect 395294 238294 395362 238350
rect 395418 238294 395488 238350
rect 395168 238226 395488 238294
rect 395168 238170 395238 238226
rect 395294 238170 395362 238226
rect 395418 238170 395488 238226
rect 395168 238102 395488 238170
rect 395168 238046 395238 238102
rect 395294 238046 395362 238102
rect 395418 238046 395488 238102
rect 395168 237978 395488 238046
rect 395168 237922 395238 237978
rect 395294 237922 395362 237978
rect 395418 237922 395488 237978
rect 395168 237888 395488 237922
rect 425888 238350 426208 238384
rect 425888 238294 425958 238350
rect 426014 238294 426082 238350
rect 426138 238294 426208 238350
rect 425888 238226 426208 238294
rect 425888 238170 425958 238226
rect 426014 238170 426082 238226
rect 426138 238170 426208 238226
rect 425888 238102 426208 238170
rect 425888 238046 425958 238102
rect 426014 238046 426082 238102
rect 426138 238046 426208 238102
rect 425888 237978 426208 238046
rect 425888 237922 425958 237978
rect 426014 237922 426082 237978
rect 426138 237922 426208 237978
rect 425888 237888 426208 237922
rect 456608 238350 456928 238384
rect 456608 238294 456678 238350
rect 456734 238294 456802 238350
rect 456858 238294 456928 238350
rect 456608 238226 456928 238294
rect 456608 238170 456678 238226
rect 456734 238170 456802 238226
rect 456858 238170 456928 238226
rect 456608 238102 456928 238170
rect 456608 238046 456678 238102
rect 456734 238046 456802 238102
rect 456858 238046 456928 238102
rect 456608 237978 456928 238046
rect 456608 237922 456678 237978
rect 456734 237922 456802 237978
rect 456858 237922 456928 237978
rect 456608 237888 456928 237922
rect 487328 238350 487648 238384
rect 487328 238294 487398 238350
rect 487454 238294 487522 238350
rect 487578 238294 487648 238350
rect 487328 238226 487648 238294
rect 487328 238170 487398 238226
rect 487454 238170 487522 238226
rect 487578 238170 487648 238226
rect 487328 238102 487648 238170
rect 487328 238046 487398 238102
rect 487454 238046 487522 238102
rect 487578 238046 487648 238102
rect 487328 237978 487648 238046
rect 487328 237922 487398 237978
rect 487454 237922 487522 237978
rect 487578 237922 487648 237978
rect 487328 237888 487648 237922
rect 518048 238350 518368 238384
rect 518048 238294 518118 238350
rect 518174 238294 518242 238350
rect 518298 238294 518368 238350
rect 518048 238226 518368 238294
rect 518048 238170 518118 238226
rect 518174 238170 518242 238226
rect 518298 238170 518368 238226
rect 518048 238102 518368 238170
rect 518048 238046 518118 238102
rect 518174 238046 518242 238102
rect 518298 238046 518368 238102
rect 518048 237978 518368 238046
rect 518048 237922 518118 237978
rect 518174 237922 518242 237978
rect 518298 237922 518368 237978
rect 518048 237888 518368 237922
rect 548768 238350 549088 238384
rect 548768 238294 548838 238350
rect 548894 238294 548962 238350
rect 549018 238294 549088 238350
rect 548768 238226 549088 238294
rect 548768 238170 548838 238226
rect 548894 238170 548962 238226
rect 549018 238170 549088 238226
rect 548768 238102 549088 238170
rect 548768 238046 548838 238102
rect 548894 238046 548962 238102
rect 549018 238046 549088 238102
rect 548768 237978 549088 238046
rect 548768 237922 548838 237978
rect 548894 237922 548962 237978
rect 549018 237922 549088 237978
rect 548768 237888 549088 237922
rect 379808 226350 380128 226384
rect 379808 226294 379878 226350
rect 379934 226294 380002 226350
rect 380058 226294 380128 226350
rect 379808 226226 380128 226294
rect 379808 226170 379878 226226
rect 379934 226170 380002 226226
rect 380058 226170 380128 226226
rect 379808 226102 380128 226170
rect 379808 226046 379878 226102
rect 379934 226046 380002 226102
rect 380058 226046 380128 226102
rect 379808 225978 380128 226046
rect 379808 225922 379878 225978
rect 379934 225922 380002 225978
rect 380058 225922 380128 225978
rect 379808 225888 380128 225922
rect 410528 226350 410848 226384
rect 410528 226294 410598 226350
rect 410654 226294 410722 226350
rect 410778 226294 410848 226350
rect 410528 226226 410848 226294
rect 410528 226170 410598 226226
rect 410654 226170 410722 226226
rect 410778 226170 410848 226226
rect 410528 226102 410848 226170
rect 410528 226046 410598 226102
rect 410654 226046 410722 226102
rect 410778 226046 410848 226102
rect 410528 225978 410848 226046
rect 410528 225922 410598 225978
rect 410654 225922 410722 225978
rect 410778 225922 410848 225978
rect 410528 225888 410848 225922
rect 441248 226350 441568 226384
rect 441248 226294 441318 226350
rect 441374 226294 441442 226350
rect 441498 226294 441568 226350
rect 441248 226226 441568 226294
rect 441248 226170 441318 226226
rect 441374 226170 441442 226226
rect 441498 226170 441568 226226
rect 441248 226102 441568 226170
rect 441248 226046 441318 226102
rect 441374 226046 441442 226102
rect 441498 226046 441568 226102
rect 441248 225978 441568 226046
rect 441248 225922 441318 225978
rect 441374 225922 441442 225978
rect 441498 225922 441568 225978
rect 441248 225888 441568 225922
rect 471968 226350 472288 226384
rect 471968 226294 472038 226350
rect 472094 226294 472162 226350
rect 472218 226294 472288 226350
rect 471968 226226 472288 226294
rect 471968 226170 472038 226226
rect 472094 226170 472162 226226
rect 472218 226170 472288 226226
rect 471968 226102 472288 226170
rect 471968 226046 472038 226102
rect 472094 226046 472162 226102
rect 472218 226046 472288 226102
rect 471968 225978 472288 226046
rect 471968 225922 472038 225978
rect 472094 225922 472162 225978
rect 472218 225922 472288 225978
rect 471968 225888 472288 225922
rect 502688 226350 503008 226384
rect 502688 226294 502758 226350
rect 502814 226294 502882 226350
rect 502938 226294 503008 226350
rect 502688 226226 503008 226294
rect 502688 226170 502758 226226
rect 502814 226170 502882 226226
rect 502938 226170 503008 226226
rect 502688 226102 503008 226170
rect 502688 226046 502758 226102
rect 502814 226046 502882 226102
rect 502938 226046 503008 226102
rect 502688 225978 503008 226046
rect 502688 225922 502758 225978
rect 502814 225922 502882 225978
rect 502938 225922 503008 225978
rect 502688 225888 503008 225922
rect 533408 226350 533728 226384
rect 533408 226294 533478 226350
rect 533534 226294 533602 226350
rect 533658 226294 533728 226350
rect 533408 226226 533728 226294
rect 533408 226170 533478 226226
rect 533534 226170 533602 226226
rect 533658 226170 533728 226226
rect 533408 226102 533728 226170
rect 533408 226046 533478 226102
rect 533534 226046 533602 226102
rect 533658 226046 533728 226102
rect 533408 225978 533728 226046
rect 533408 225922 533478 225978
rect 533534 225922 533602 225978
rect 533658 225922 533728 225978
rect 533408 225888 533728 225922
rect 364448 220350 364768 220384
rect 364448 220294 364518 220350
rect 364574 220294 364642 220350
rect 364698 220294 364768 220350
rect 364448 220226 364768 220294
rect 364448 220170 364518 220226
rect 364574 220170 364642 220226
rect 364698 220170 364768 220226
rect 364448 220102 364768 220170
rect 364448 220046 364518 220102
rect 364574 220046 364642 220102
rect 364698 220046 364768 220102
rect 364448 219978 364768 220046
rect 364448 219922 364518 219978
rect 364574 219922 364642 219978
rect 364698 219922 364768 219978
rect 364448 219888 364768 219922
rect 395168 220350 395488 220384
rect 395168 220294 395238 220350
rect 395294 220294 395362 220350
rect 395418 220294 395488 220350
rect 395168 220226 395488 220294
rect 395168 220170 395238 220226
rect 395294 220170 395362 220226
rect 395418 220170 395488 220226
rect 395168 220102 395488 220170
rect 395168 220046 395238 220102
rect 395294 220046 395362 220102
rect 395418 220046 395488 220102
rect 395168 219978 395488 220046
rect 395168 219922 395238 219978
rect 395294 219922 395362 219978
rect 395418 219922 395488 219978
rect 395168 219888 395488 219922
rect 425888 220350 426208 220384
rect 425888 220294 425958 220350
rect 426014 220294 426082 220350
rect 426138 220294 426208 220350
rect 425888 220226 426208 220294
rect 425888 220170 425958 220226
rect 426014 220170 426082 220226
rect 426138 220170 426208 220226
rect 425888 220102 426208 220170
rect 425888 220046 425958 220102
rect 426014 220046 426082 220102
rect 426138 220046 426208 220102
rect 425888 219978 426208 220046
rect 425888 219922 425958 219978
rect 426014 219922 426082 219978
rect 426138 219922 426208 219978
rect 425888 219888 426208 219922
rect 456608 220350 456928 220384
rect 456608 220294 456678 220350
rect 456734 220294 456802 220350
rect 456858 220294 456928 220350
rect 456608 220226 456928 220294
rect 456608 220170 456678 220226
rect 456734 220170 456802 220226
rect 456858 220170 456928 220226
rect 456608 220102 456928 220170
rect 456608 220046 456678 220102
rect 456734 220046 456802 220102
rect 456858 220046 456928 220102
rect 456608 219978 456928 220046
rect 456608 219922 456678 219978
rect 456734 219922 456802 219978
rect 456858 219922 456928 219978
rect 456608 219888 456928 219922
rect 487328 220350 487648 220384
rect 487328 220294 487398 220350
rect 487454 220294 487522 220350
rect 487578 220294 487648 220350
rect 487328 220226 487648 220294
rect 487328 220170 487398 220226
rect 487454 220170 487522 220226
rect 487578 220170 487648 220226
rect 487328 220102 487648 220170
rect 487328 220046 487398 220102
rect 487454 220046 487522 220102
rect 487578 220046 487648 220102
rect 487328 219978 487648 220046
rect 487328 219922 487398 219978
rect 487454 219922 487522 219978
rect 487578 219922 487648 219978
rect 487328 219888 487648 219922
rect 518048 220350 518368 220384
rect 518048 220294 518118 220350
rect 518174 220294 518242 220350
rect 518298 220294 518368 220350
rect 518048 220226 518368 220294
rect 518048 220170 518118 220226
rect 518174 220170 518242 220226
rect 518298 220170 518368 220226
rect 518048 220102 518368 220170
rect 518048 220046 518118 220102
rect 518174 220046 518242 220102
rect 518298 220046 518368 220102
rect 518048 219978 518368 220046
rect 518048 219922 518118 219978
rect 518174 219922 518242 219978
rect 518298 219922 518368 219978
rect 518048 219888 518368 219922
rect 548768 220350 549088 220384
rect 548768 220294 548838 220350
rect 548894 220294 548962 220350
rect 549018 220294 549088 220350
rect 548768 220226 549088 220294
rect 548768 220170 548838 220226
rect 548894 220170 548962 220226
rect 549018 220170 549088 220226
rect 548768 220102 549088 220170
rect 548768 220046 548838 220102
rect 548894 220046 548962 220102
rect 549018 220046 549088 220102
rect 548768 219978 549088 220046
rect 548768 219922 548838 219978
rect 548894 219922 548962 219978
rect 549018 219922 549088 219978
rect 548768 219888 549088 219922
rect 379808 208350 380128 208384
rect 379808 208294 379878 208350
rect 379934 208294 380002 208350
rect 380058 208294 380128 208350
rect 379808 208226 380128 208294
rect 379808 208170 379878 208226
rect 379934 208170 380002 208226
rect 380058 208170 380128 208226
rect 379808 208102 380128 208170
rect 379808 208046 379878 208102
rect 379934 208046 380002 208102
rect 380058 208046 380128 208102
rect 379808 207978 380128 208046
rect 379808 207922 379878 207978
rect 379934 207922 380002 207978
rect 380058 207922 380128 207978
rect 379808 207888 380128 207922
rect 410528 208350 410848 208384
rect 410528 208294 410598 208350
rect 410654 208294 410722 208350
rect 410778 208294 410848 208350
rect 410528 208226 410848 208294
rect 410528 208170 410598 208226
rect 410654 208170 410722 208226
rect 410778 208170 410848 208226
rect 410528 208102 410848 208170
rect 410528 208046 410598 208102
rect 410654 208046 410722 208102
rect 410778 208046 410848 208102
rect 410528 207978 410848 208046
rect 410528 207922 410598 207978
rect 410654 207922 410722 207978
rect 410778 207922 410848 207978
rect 410528 207888 410848 207922
rect 441248 208350 441568 208384
rect 441248 208294 441318 208350
rect 441374 208294 441442 208350
rect 441498 208294 441568 208350
rect 441248 208226 441568 208294
rect 441248 208170 441318 208226
rect 441374 208170 441442 208226
rect 441498 208170 441568 208226
rect 441248 208102 441568 208170
rect 441248 208046 441318 208102
rect 441374 208046 441442 208102
rect 441498 208046 441568 208102
rect 441248 207978 441568 208046
rect 441248 207922 441318 207978
rect 441374 207922 441442 207978
rect 441498 207922 441568 207978
rect 441248 207888 441568 207922
rect 471968 208350 472288 208384
rect 471968 208294 472038 208350
rect 472094 208294 472162 208350
rect 472218 208294 472288 208350
rect 471968 208226 472288 208294
rect 471968 208170 472038 208226
rect 472094 208170 472162 208226
rect 472218 208170 472288 208226
rect 471968 208102 472288 208170
rect 471968 208046 472038 208102
rect 472094 208046 472162 208102
rect 472218 208046 472288 208102
rect 471968 207978 472288 208046
rect 471968 207922 472038 207978
rect 472094 207922 472162 207978
rect 472218 207922 472288 207978
rect 471968 207888 472288 207922
rect 502688 208350 503008 208384
rect 502688 208294 502758 208350
rect 502814 208294 502882 208350
rect 502938 208294 503008 208350
rect 502688 208226 503008 208294
rect 502688 208170 502758 208226
rect 502814 208170 502882 208226
rect 502938 208170 503008 208226
rect 502688 208102 503008 208170
rect 502688 208046 502758 208102
rect 502814 208046 502882 208102
rect 502938 208046 503008 208102
rect 502688 207978 503008 208046
rect 502688 207922 502758 207978
rect 502814 207922 502882 207978
rect 502938 207922 503008 207978
rect 502688 207888 503008 207922
rect 533408 208350 533728 208384
rect 533408 208294 533478 208350
rect 533534 208294 533602 208350
rect 533658 208294 533728 208350
rect 533408 208226 533728 208294
rect 533408 208170 533478 208226
rect 533534 208170 533602 208226
rect 533658 208170 533728 208226
rect 533408 208102 533728 208170
rect 533408 208046 533478 208102
rect 533534 208046 533602 208102
rect 533658 208046 533728 208102
rect 533408 207978 533728 208046
rect 533408 207922 533478 207978
rect 533534 207922 533602 207978
rect 533658 207922 533728 207978
rect 533408 207888 533728 207922
rect 364448 202350 364768 202384
rect 364448 202294 364518 202350
rect 364574 202294 364642 202350
rect 364698 202294 364768 202350
rect 364448 202226 364768 202294
rect 364448 202170 364518 202226
rect 364574 202170 364642 202226
rect 364698 202170 364768 202226
rect 364448 202102 364768 202170
rect 364448 202046 364518 202102
rect 364574 202046 364642 202102
rect 364698 202046 364768 202102
rect 364448 201978 364768 202046
rect 364448 201922 364518 201978
rect 364574 201922 364642 201978
rect 364698 201922 364768 201978
rect 364448 201888 364768 201922
rect 395168 202350 395488 202384
rect 395168 202294 395238 202350
rect 395294 202294 395362 202350
rect 395418 202294 395488 202350
rect 395168 202226 395488 202294
rect 395168 202170 395238 202226
rect 395294 202170 395362 202226
rect 395418 202170 395488 202226
rect 395168 202102 395488 202170
rect 395168 202046 395238 202102
rect 395294 202046 395362 202102
rect 395418 202046 395488 202102
rect 395168 201978 395488 202046
rect 395168 201922 395238 201978
rect 395294 201922 395362 201978
rect 395418 201922 395488 201978
rect 395168 201888 395488 201922
rect 425888 202350 426208 202384
rect 425888 202294 425958 202350
rect 426014 202294 426082 202350
rect 426138 202294 426208 202350
rect 425888 202226 426208 202294
rect 425888 202170 425958 202226
rect 426014 202170 426082 202226
rect 426138 202170 426208 202226
rect 425888 202102 426208 202170
rect 425888 202046 425958 202102
rect 426014 202046 426082 202102
rect 426138 202046 426208 202102
rect 425888 201978 426208 202046
rect 425888 201922 425958 201978
rect 426014 201922 426082 201978
rect 426138 201922 426208 201978
rect 425888 201888 426208 201922
rect 456608 202350 456928 202384
rect 456608 202294 456678 202350
rect 456734 202294 456802 202350
rect 456858 202294 456928 202350
rect 456608 202226 456928 202294
rect 456608 202170 456678 202226
rect 456734 202170 456802 202226
rect 456858 202170 456928 202226
rect 456608 202102 456928 202170
rect 456608 202046 456678 202102
rect 456734 202046 456802 202102
rect 456858 202046 456928 202102
rect 456608 201978 456928 202046
rect 456608 201922 456678 201978
rect 456734 201922 456802 201978
rect 456858 201922 456928 201978
rect 456608 201888 456928 201922
rect 487328 202350 487648 202384
rect 487328 202294 487398 202350
rect 487454 202294 487522 202350
rect 487578 202294 487648 202350
rect 487328 202226 487648 202294
rect 487328 202170 487398 202226
rect 487454 202170 487522 202226
rect 487578 202170 487648 202226
rect 487328 202102 487648 202170
rect 487328 202046 487398 202102
rect 487454 202046 487522 202102
rect 487578 202046 487648 202102
rect 487328 201978 487648 202046
rect 487328 201922 487398 201978
rect 487454 201922 487522 201978
rect 487578 201922 487648 201978
rect 487328 201888 487648 201922
rect 518048 202350 518368 202384
rect 518048 202294 518118 202350
rect 518174 202294 518242 202350
rect 518298 202294 518368 202350
rect 518048 202226 518368 202294
rect 518048 202170 518118 202226
rect 518174 202170 518242 202226
rect 518298 202170 518368 202226
rect 518048 202102 518368 202170
rect 518048 202046 518118 202102
rect 518174 202046 518242 202102
rect 518298 202046 518368 202102
rect 518048 201978 518368 202046
rect 518048 201922 518118 201978
rect 518174 201922 518242 201978
rect 518298 201922 518368 201978
rect 518048 201888 518368 201922
rect 548768 202350 549088 202384
rect 548768 202294 548838 202350
rect 548894 202294 548962 202350
rect 549018 202294 549088 202350
rect 548768 202226 549088 202294
rect 548768 202170 548838 202226
rect 548894 202170 548962 202226
rect 549018 202170 549088 202226
rect 548768 202102 549088 202170
rect 548768 202046 548838 202102
rect 548894 202046 548962 202102
rect 549018 202046 549088 202102
rect 548768 201978 549088 202046
rect 548768 201922 548838 201978
rect 548894 201922 548962 201978
rect 549018 201922 549088 201978
rect 548768 201888 549088 201922
rect 362124 195778 362180 195788
rect 362124 174468 362180 195722
rect 379808 190350 380128 190384
rect 379808 190294 379878 190350
rect 379934 190294 380002 190350
rect 380058 190294 380128 190350
rect 379808 190226 380128 190294
rect 379808 190170 379878 190226
rect 379934 190170 380002 190226
rect 380058 190170 380128 190226
rect 379808 190102 380128 190170
rect 379808 190046 379878 190102
rect 379934 190046 380002 190102
rect 380058 190046 380128 190102
rect 379808 189978 380128 190046
rect 379808 189922 379878 189978
rect 379934 189922 380002 189978
rect 380058 189922 380128 189978
rect 379808 189888 380128 189922
rect 410528 190350 410848 190384
rect 410528 190294 410598 190350
rect 410654 190294 410722 190350
rect 410778 190294 410848 190350
rect 410528 190226 410848 190294
rect 410528 190170 410598 190226
rect 410654 190170 410722 190226
rect 410778 190170 410848 190226
rect 410528 190102 410848 190170
rect 410528 190046 410598 190102
rect 410654 190046 410722 190102
rect 410778 190046 410848 190102
rect 410528 189978 410848 190046
rect 410528 189922 410598 189978
rect 410654 189922 410722 189978
rect 410778 189922 410848 189978
rect 410528 189888 410848 189922
rect 441248 190350 441568 190384
rect 441248 190294 441318 190350
rect 441374 190294 441442 190350
rect 441498 190294 441568 190350
rect 441248 190226 441568 190294
rect 441248 190170 441318 190226
rect 441374 190170 441442 190226
rect 441498 190170 441568 190226
rect 441248 190102 441568 190170
rect 441248 190046 441318 190102
rect 441374 190046 441442 190102
rect 441498 190046 441568 190102
rect 441248 189978 441568 190046
rect 441248 189922 441318 189978
rect 441374 189922 441442 189978
rect 441498 189922 441568 189978
rect 441248 189888 441568 189922
rect 471968 190350 472288 190384
rect 471968 190294 472038 190350
rect 472094 190294 472162 190350
rect 472218 190294 472288 190350
rect 471968 190226 472288 190294
rect 471968 190170 472038 190226
rect 472094 190170 472162 190226
rect 472218 190170 472288 190226
rect 471968 190102 472288 190170
rect 471968 190046 472038 190102
rect 472094 190046 472162 190102
rect 472218 190046 472288 190102
rect 471968 189978 472288 190046
rect 471968 189922 472038 189978
rect 472094 189922 472162 189978
rect 472218 189922 472288 189978
rect 471968 189888 472288 189922
rect 502688 190350 503008 190384
rect 502688 190294 502758 190350
rect 502814 190294 502882 190350
rect 502938 190294 503008 190350
rect 502688 190226 503008 190294
rect 502688 190170 502758 190226
rect 502814 190170 502882 190226
rect 502938 190170 503008 190226
rect 502688 190102 503008 190170
rect 502688 190046 502758 190102
rect 502814 190046 502882 190102
rect 502938 190046 503008 190102
rect 502688 189978 503008 190046
rect 502688 189922 502758 189978
rect 502814 189922 502882 189978
rect 502938 189922 503008 189978
rect 502688 189888 503008 189922
rect 533408 190350 533728 190384
rect 533408 190294 533478 190350
rect 533534 190294 533602 190350
rect 533658 190294 533728 190350
rect 533408 190226 533728 190294
rect 533408 190170 533478 190226
rect 533534 190170 533602 190226
rect 533658 190170 533728 190226
rect 533408 190102 533728 190170
rect 533408 190046 533478 190102
rect 533534 190046 533602 190102
rect 533658 190046 533728 190102
rect 533408 189978 533728 190046
rect 533408 189922 533478 189978
rect 533534 189922 533602 189978
rect 533658 189922 533728 189978
rect 533408 189888 533728 189922
rect 364448 184350 364768 184384
rect 364448 184294 364518 184350
rect 364574 184294 364642 184350
rect 364698 184294 364768 184350
rect 364448 184226 364768 184294
rect 364448 184170 364518 184226
rect 364574 184170 364642 184226
rect 364698 184170 364768 184226
rect 364448 184102 364768 184170
rect 364448 184046 364518 184102
rect 364574 184046 364642 184102
rect 364698 184046 364768 184102
rect 364448 183978 364768 184046
rect 364448 183922 364518 183978
rect 364574 183922 364642 183978
rect 364698 183922 364768 183978
rect 364448 183888 364768 183922
rect 395168 184350 395488 184384
rect 395168 184294 395238 184350
rect 395294 184294 395362 184350
rect 395418 184294 395488 184350
rect 395168 184226 395488 184294
rect 395168 184170 395238 184226
rect 395294 184170 395362 184226
rect 395418 184170 395488 184226
rect 395168 184102 395488 184170
rect 395168 184046 395238 184102
rect 395294 184046 395362 184102
rect 395418 184046 395488 184102
rect 395168 183978 395488 184046
rect 395168 183922 395238 183978
rect 395294 183922 395362 183978
rect 395418 183922 395488 183978
rect 395168 183888 395488 183922
rect 425888 184350 426208 184384
rect 425888 184294 425958 184350
rect 426014 184294 426082 184350
rect 426138 184294 426208 184350
rect 425888 184226 426208 184294
rect 425888 184170 425958 184226
rect 426014 184170 426082 184226
rect 426138 184170 426208 184226
rect 425888 184102 426208 184170
rect 425888 184046 425958 184102
rect 426014 184046 426082 184102
rect 426138 184046 426208 184102
rect 425888 183978 426208 184046
rect 425888 183922 425958 183978
rect 426014 183922 426082 183978
rect 426138 183922 426208 183978
rect 425888 183888 426208 183922
rect 456608 184350 456928 184384
rect 456608 184294 456678 184350
rect 456734 184294 456802 184350
rect 456858 184294 456928 184350
rect 456608 184226 456928 184294
rect 456608 184170 456678 184226
rect 456734 184170 456802 184226
rect 456858 184170 456928 184226
rect 456608 184102 456928 184170
rect 456608 184046 456678 184102
rect 456734 184046 456802 184102
rect 456858 184046 456928 184102
rect 456608 183978 456928 184046
rect 456608 183922 456678 183978
rect 456734 183922 456802 183978
rect 456858 183922 456928 183978
rect 456608 183888 456928 183922
rect 487328 184350 487648 184384
rect 487328 184294 487398 184350
rect 487454 184294 487522 184350
rect 487578 184294 487648 184350
rect 487328 184226 487648 184294
rect 487328 184170 487398 184226
rect 487454 184170 487522 184226
rect 487578 184170 487648 184226
rect 487328 184102 487648 184170
rect 487328 184046 487398 184102
rect 487454 184046 487522 184102
rect 487578 184046 487648 184102
rect 487328 183978 487648 184046
rect 487328 183922 487398 183978
rect 487454 183922 487522 183978
rect 487578 183922 487648 183978
rect 487328 183888 487648 183922
rect 518048 184350 518368 184384
rect 518048 184294 518118 184350
rect 518174 184294 518242 184350
rect 518298 184294 518368 184350
rect 518048 184226 518368 184294
rect 518048 184170 518118 184226
rect 518174 184170 518242 184226
rect 518298 184170 518368 184226
rect 518048 184102 518368 184170
rect 518048 184046 518118 184102
rect 518174 184046 518242 184102
rect 518298 184046 518368 184102
rect 518048 183978 518368 184046
rect 518048 183922 518118 183978
rect 518174 183922 518242 183978
rect 518298 183922 518368 183978
rect 518048 183888 518368 183922
rect 548768 184350 549088 184384
rect 548768 184294 548838 184350
rect 548894 184294 548962 184350
rect 549018 184294 549088 184350
rect 548768 184226 549088 184294
rect 548768 184170 548838 184226
rect 548894 184170 548962 184226
rect 549018 184170 549088 184226
rect 548768 184102 549088 184170
rect 548768 184046 548838 184102
rect 548894 184046 548962 184102
rect 549018 184046 549088 184102
rect 548768 183978 549088 184046
rect 548768 183922 548838 183978
rect 548894 183922 548962 183978
rect 549018 183922 549088 183978
rect 548768 183888 549088 183922
rect 375228 175258 375284 175290
rect 375228 175186 375284 175196
rect 362124 174402 362180 174412
rect 417564 174692 417620 174702
rect 417564 173998 417620 174636
rect 417564 173932 417620 173942
rect 362012 118626 362068 118636
rect 374058 166350 374678 173466
rect 374058 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 374678 166350
rect 374058 166226 374678 166294
rect 374058 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 374678 166226
rect 374058 166102 374678 166170
rect 374058 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 374678 166102
rect 374058 165978 374678 166046
rect 374058 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 374678 165978
rect 374058 148350 374678 165922
rect 374058 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 374678 148350
rect 374058 148226 374678 148294
rect 374058 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 374678 148226
rect 374058 148102 374678 148170
rect 374058 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 374678 148102
rect 374058 147978 374678 148046
rect 374058 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 374678 147978
rect 374058 130350 374678 147922
rect 374058 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 374678 130350
rect 374058 130226 374678 130294
rect 374058 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 374678 130226
rect 374058 130102 374678 130170
rect 374058 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 374678 130102
rect 374058 129978 374678 130046
rect 374058 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 374678 129978
rect 361788 118514 361844 118524
rect 360444 117058 360500 117068
rect 359884 115792 359940 115802
rect 374058 115262 374678 129922
rect 377778 172350 378398 173466
rect 377778 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 378398 172350
rect 377778 172226 378398 172294
rect 377778 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 378398 172226
rect 377778 172102 378398 172170
rect 377778 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 378398 172102
rect 377778 171978 378398 172046
rect 377778 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 378398 171978
rect 377778 154350 378398 171922
rect 377778 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 378398 154350
rect 377778 154226 378398 154294
rect 377778 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 378398 154226
rect 377778 154102 378398 154170
rect 377778 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 378398 154102
rect 377778 153978 378398 154046
rect 377778 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 378398 153978
rect 377778 136350 378398 153922
rect 377778 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 378398 136350
rect 377778 136226 378398 136294
rect 377778 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 378398 136226
rect 377778 136102 378398 136170
rect 377778 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 378398 136102
rect 377778 135978 378398 136046
rect 377778 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 378398 135978
rect 377778 118350 378398 135922
rect 404778 166350 405398 173466
rect 404778 166294 404874 166350
rect 404930 166294 404998 166350
rect 405054 166294 405122 166350
rect 405178 166294 405246 166350
rect 405302 166294 405398 166350
rect 404778 166226 405398 166294
rect 404778 166170 404874 166226
rect 404930 166170 404998 166226
rect 405054 166170 405122 166226
rect 405178 166170 405246 166226
rect 405302 166170 405398 166226
rect 404778 166102 405398 166170
rect 404778 166046 404874 166102
rect 404930 166046 404998 166102
rect 405054 166046 405122 166102
rect 405178 166046 405246 166102
rect 405302 166046 405398 166102
rect 404778 165978 405398 166046
rect 404778 165922 404874 165978
rect 404930 165922 404998 165978
rect 405054 165922 405122 165978
rect 405178 165922 405246 165978
rect 405302 165922 405398 165978
rect 404778 148350 405398 165922
rect 404778 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 405398 148350
rect 404778 148226 405398 148294
rect 404778 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 405398 148226
rect 404778 148102 405398 148170
rect 404778 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 405398 148102
rect 404778 147978 405398 148046
rect 404778 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 405398 147978
rect 404778 130350 405398 147922
rect 404778 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 405398 130350
rect 404778 130226 405398 130294
rect 404778 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 405398 130226
rect 404778 130102 405398 130170
rect 404778 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 405398 130102
rect 404778 129978 405398 130046
rect 404778 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 405398 129978
rect 394940 124318 394996 124328
rect 388892 124138 388948 124148
rect 386876 123778 386932 123788
rect 384860 123598 384916 123608
rect 384860 122724 384916 123542
rect 384860 122658 384916 122668
rect 386876 122724 386932 123722
rect 386876 122658 386932 122668
rect 388892 122724 388948 124082
rect 388892 122658 388948 122668
rect 390908 123958 390964 123968
rect 390908 122724 390964 123902
rect 390908 122658 390964 122668
rect 394940 122724 394996 124262
rect 394940 122658 394996 122668
rect 377778 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 378398 118350
rect 377778 118226 378398 118294
rect 377778 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 378398 118226
rect 377778 118102 378398 118170
rect 377778 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 378398 118102
rect 377778 117978 378398 118046
rect 377778 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 378398 117978
rect 377778 115262 378398 117922
rect 404778 115262 405398 129922
rect 408498 172350 409118 173466
rect 408498 172294 408594 172350
rect 408650 172294 408718 172350
rect 408774 172294 408842 172350
rect 408898 172294 408966 172350
rect 409022 172294 409118 172350
rect 408498 172226 409118 172294
rect 408498 172170 408594 172226
rect 408650 172170 408718 172226
rect 408774 172170 408842 172226
rect 408898 172170 408966 172226
rect 409022 172170 409118 172226
rect 408498 172102 409118 172170
rect 408498 172046 408594 172102
rect 408650 172046 408718 172102
rect 408774 172046 408842 172102
rect 408898 172046 408966 172102
rect 409022 172046 409118 172102
rect 408498 171978 409118 172046
rect 408498 171922 408594 171978
rect 408650 171922 408718 171978
rect 408774 171922 408842 171978
rect 408898 171922 408966 171978
rect 409022 171922 409118 171978
rect 408498 154350 409118 171922
rect 408498 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 409118 154350
rect 408498 154226 409118 154294
rect 408498 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 409118 154226
rect 408498 154102 409118 154170
rect 408498 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 409118 154102
rect 408498 153978 409118 154046
rect 408498 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 409118 153978
rect 408498 136350 409118 153922
rect 435498 166350 436118 173466
rect 435498 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 436118 166350
rect 435498 166226 436118 166294
rect 435498 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 436118 166226
rect 435498 166102 436118 166170
rect 435498 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 436118 166102
rect 435498 165978 436118 166046
rect 435498 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 436118 165978
rect 435498 148350 436118 165922
rect 435498 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 436118 148350
rect 435498 148226 436118 148294
rect 435498 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 436118 148226
rect 435498 148102 436118 148170
rect 435498 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 436118 148102
rect 435498 147978 436118 148046
rect 435498 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 436118 147978
rect 408498 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 409118 136350
rect 408498 136226 409118 136294
rect 408498 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 409118 136226
rect 408498 136102 409118 136170
rect 408498 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 409118 136102
rect 408498 135978 409118 136046
rect 408498 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 409118 135978
rect 408498 118350 409118 135922
rect 414988 136918 415044 136928
rect 411628 133498 411684 133508
rect 411628 122724 411684 133442
rect 411628 122658 411684 122668
rect 414988 122724 415044 136862
rect 414988 122658 415044 122668
rect 435498 130350 436118 147922
rect 435498 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 436118 130350
rect 435498 130226 436118 130294
rect 435498 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 436118 130226
rect 435498 130102 436118 130170
rect 435498 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 436118 130102
rect 435498 129978 436118 130046
rect 435498 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 436118 129978
rect 408498 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 409118 118350
rect 408498 118226 409118 118294
rect 408498 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 409118 118226
rect 408498 118102 409118 118170
rect 408498 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 409118 118102
rect 408498 117978 409118 118046
rect 408498 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 409118 117978
rect 408498 115262 409118 117922
rect 421708 120484 421764 120494
rect 421708 116116 421764 120428
rect 421708 116050 421764 116060
rect 421820 118804 421876 118814
rect 364448 112350 364768 112384
rect 364448 112294 364518 112350
rect 364574 112294 364642 112350
rect 364698 112294 364768 112350
rect 364448 112226 364768 112294
rect 364448 112170 364518 112226
rect 364574 112170 364642 112226
rect 364698 112170 364768 112226
rect 364448 112102 364768 112170
rect 364448 112046 364518 112102
rect 364574 112046 364642 112102
rect 364698 112046 364768 112102
rect 364448 111978 364768 112046
rect 364448 111922 364518 111978
rect 364574 111922 364642 111978
rect 364698 111922 364768 111978
rect 364448 111888 364768 111922
rect 395168 112350 395488 112384
rect 395168 112294 395238 112350
rect 395294 112294 395362 112350
rect 395418 112294 395488 112350
rect 395168 112226 395488 112294
rect 395168 112170 395238 112226
rect 395294 112170 395362 112226
rect 395418 112170 395488 112226
rect 395168 112102 395488 112170
rect 395168 112046 395238 112102
rect 395294 112046 395362 112102
rect 395418 112046 395488 112102
rect 395168 111978 395488 112046
rect 395168 111922 395238 111978
rect 395294 111922 395362 111978
rect 395418 111922 395488 111978
rect 395168 111888 395488 111922
rect 421820 109172 421876 118748
rect 425852 116116 425908 116126
rect 421820 109106 421876 109116
rect 424172 109172 424228 109182
rect 379808 100350 380128 100384
rect 379808 100294 379878 100350
rect 379934 100294 380002 100350
rect 380058 100294 380128 100350
rect 379808 100226 380128 100294
rect 379808 100170 379878 100226
rect 379934 100170 380002 100226
rect 380058 100170 380128 100226
rect 379808 100102 380128 100170
rect 379808 100046 379878 100102
rect 379934 100046 380002 100102
rect 380058 100046 380128 100102
rect 379808 99978 380128 100046
rect 379808 99922 379878 99978
rect 379934 99922 380002 99978
rect 380058 99922 380128 99978
rect 379808 99888 380128 99922
rect 410528 100350 410848 100384
rect 410528 100294 410598 100350
rect 410654 100294 410722 100350
rect 410778 100294 410848 100350
rect 410528 100226 410848 100294
rect 410528 100170 410598 100226
rect 410654 100170 410722 100226
rect 410778 100170 410848 100226
rect 410528 100102 410848 100170
rect 410528 100046 410598 100102
rect 410654 100046 410722 100102
rect 410778 100046 410848 100102
rect 410528 99978 410848 100046
rect 410528 99922 410598 99978
rect 410654 99922 410722 99978
rect 410778 99922 410848 99978
rect 410528 99888 410848 99922
rect 364448 94350 364768 94384
rect 364448 94294 364518 94350
rect 364574 94294 364642 94350
rect 364698 94294 364768 94350
rect 364448 94226 364768 94294
rect 364448 94170 364518 94226
rect 364574 94170 364642 94226
rect 364698 94170 364768 94226
rect 364448 94102 364768 94170
rect 364448 94046 364518 94102
rect 364574 94046 364642 94102
rect 364698 94046 364768 94102
rect 364448 93978 364768 94046
rect 364448 93922 364518 93978
rect 364574 93922 364642 93978
rect 364698 93922 364768 93978
rect 364448 93888 364768 93922
rect 395168 94350 395488 94384
rect 395168 94294 395238 94350
rect 395294 94294 395362 94350
rect 395418 94294 395488 94350
rect 395168 94226 395488 94294
rect 395168 94170 395238 94226
rect 395294 94170 395362 94226
rect 395418 94170 395488 94226
rect 395168 94102 395488 94170
rect 395168 94046 395238 94102
rect 395294 94046 395362 94102
rect 395418 94046 395488 94102
rect 395168 93978 395488 94046
rect 395168 93922 395238 93978
rect 395294 93922 395362 93978
rect 395418 93922 395488 93978
rect 395168 93888 395488 93922
rect 379808 82350 380128 82384
rect 379808 82294 379878 82350
rect 379934 82294 380002 82350
rect 380058 82294 380128 82350
rect 379808 82226 380128 82294
rect 379808 82170 379878 82226
rect 379934 82170 380002 82226
rect 380058 82170 380128 82226
rect 379808 82102 380128 82170
rect 379808 82046 379878 82102
rect 379934 82046 380002 82102
rect 380058 82046 380128 82102
rect 379808 81978 380128 82046
rect 379808 81922 379878 81978
rect 379934 81922 380002 81978
rect 380058 81922 380128 81978
rect 379808 81888 380128 81922
rect 410528 82350 410848 82384
rect 410528 82294 410598 82350
rect 410654 82294 410722 82350
rect 410778 82294 410848 82350
rect 410528 82226 410848 82294
rect 410528 82170 410598 82226
rect 410654 82170 410722 82226
rect 410778 82170 410848 82226
rect 410528 82102 410848 82170
rect 410528 82046 410598 82102
rect 410654 82046 410722 82102
rect 410778 82046 410848 82102
rect 410528 81978 410848 82046
rect 410528 81922 410598 81978
rect 410654 81922 410722 81978
rect 410778 81922 410848 81978
rect 410528 81888 410848 81922
rect 364448 76350 364768 76384
rect 364448 76294 364518 76350
rect 364574 76294 364642 76350
rect 364698 76294 364768 76350
rect 364448 76226 364768 76294
rect 364448 76170 364518 76226
rect 364574 76170 364642 76226
rect 364698 76170 364768 76226
rect 364448 76102 364768 76170
rect 364448 76046 364518 76102
rect 364574 76046 364642 76102
rect 364698 76046 364768 76102
rect 364448 75978 364768 76046
rect 364448 75922 364518 75978
rect 364574 75922 364642 75978
rect 364698 75922 364768 75978
rect 364448 75888 364768 75922
rect 395168 76350 395488 76384
rect 395168 76294 395238 76350
rect 395294 76294 395362 76350
rect 395418 76294 395488 76350
rect 395168 76226 395488 76294
rect 395168 76170 395238 76226
rect 395294 76170 395362 76226
rect 395418 76170 395488 76226
rect 395168 76102 395488 76170
rect 395168 76046 395238 76102
rect 395294 76046 395362 76102
rect 395418 76046 395488 76102
rect 395168 75978 395488 76046
rect 395168 75922 395238 75978
rect 395294 75922 395362 75978
rect 395418 75922 395488 75978
rect 395168 75888 395488 75922
rect 424172 66388 424228 109116
rect 424172 66322 424228 66332
rect 379808 64350 380128 64384
rect 379808 64294 379878 64350
rect 379934 64294 380002 64350
rect 380058 64294 380128 64350
rect 379808 64226 380128 64294
rect 379808 64170 379878 64226
rect 379934 64170 380002 64226
rect 380058 64170 380128 64226
rect 379808 64102 380128 64170
rect 379808 64046 379878 64102
rect 379934 64046 380002 64102
rect 380058 64046 380128 64102
rect 379808 63978 380128 64046
rect 379808 63922 379878 63978
rect 379934 63922 380002 63978
rect 380058 63922 380128 63978
rect 379808 63888 380128 63922
rect 410528 64350 410848 64384
rect 410528 64294 410598 64350
rect 410654 64294 410722 64350
rect 410778 64294 410848 64350
rect 410528 64226 410848 64294
rect 410528 64170 410598 64226
rect 410654 64170 410722 64226
rect 410778 64170 410848 64226
rect 410528 64102 410848 64170
rect 410528 64046 410598 64102
rect 410654 64046 410722 64102
rect 410778 64046 410848 64102
rect 410528 63978 410848 64046
rect 410528 63922 410598 63978
rect 410654 63922 410722 63978
rect 410778 63922 410848 63978
rect 410528 63888 410848 63922
rect 425852 60676 425908 116060
rect 425852 60610 425908 60620
rect 435498 112350 436118 129922
rect 435498 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 436118 112350
rect 435498 112226 436118 112294
rect 435498 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 436118 112226
rect 435498 112102 436118 112170
rect 435498 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 436118 112102
rect 435498 111978 436118 112046
rect 435498 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 436118 111978
rect 435498 94350 436118 111922
rect 435498 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 436118 94350
rect 435498 94226 436118 94294
rect 435498 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 436118 94226
rect 435498 94102 436118 94170
rect 435498 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 436118 94102
rect 435498 93978 436118 94046
rect 435498 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 436118 93978
rect 435498 76350 436118 93922
rect 435498 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 436118 76350
rect 435498 76226 436118 76294
rect 435498 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 436118 76226
rect 435498 76102 436118 76170
rect 435498 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 436118 76102
rect 435498 75978 436118 76046
rect 435498 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 436118 75978
rect 364448 58350 364768 58384
rect 364448 58294 364518 58350
rect 364574 58294 364642 58350
rect 364698 58294 364768 58350
rect 364448 58226 364768 58294
rect 364448 58170 364518 58226
rect 364574 58170 364642 58226
rect 364698 58170 364768 58226
rect 364448 58102 364768 58170
rect 364448 58046 364518 58102
rect 364574 58046 364642 58102
rect 364698 58046 364768 58102
rect 364448 57978 364768 58046
rect 364448 57922 364518 57978
rect 364574 57922 364642 57978
rect 364698 57922 364768 57978
rect 364448 57888 364768 57922
rect 395168 58350 395488 58384
rect 395168 58294 395238 58350
rect 395294 58294 395362 58350
rect 395418 58294 395488 58350
rect 395168 58226 395488 58294
rect 395168 58170 395238 58226
rect 395294 58170 395362 58226
rect 395418 58170 395488 58226
rect 395168 58102 395488 58170
rect 395168 58046 395238 58102
rect 395294 58046 395362 58102
rect 395418 58046 395488 58102
rect 395168 57978 395488 58046
rect 395168 57922 395238 57978
rect 395294 57922 395362 57978
rect 395418 57922 395488 57978
rect 395168 57888 395488 57922
rect 435498 58350 436118 75922
rect 435498 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 436118 58350
rect 435498 58226 436118 58294
rect 435498 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 436118 58226
rect 435498 58102 436118 58170
rect 435498 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 436118 58102
rect 435498 57978 436118 58046
rect 435498 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 436118 57978
rect 359772 45042 359828 45052
rect 347058 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 347678 28350
rect 347058 28226 347678 28294
rect 347058 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 347678 28226
rect 347058 28102 347678 28170
rect 347058 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 347678 28102
rect 347058 27978 347678 28046
rect 347058 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 347678 27978
rect 347058 10350 347678 27922
rect 347058 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 347678 10350
rect 347058 10226 347678 10294
rect 347058 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 347678 10226
rect 347058 10102 347678 10170
rect 347058 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 347678 10102
rect 347058 9978 347678 10046
rect 347058 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 347678 9978
rect 347058 -1120 347678 9922
rect 347058 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 347678 -1120
rect 347058 -1244 347678 -1176
rect 347058 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 347678 -1244
rect 347058 -1368 347678 -1300
rect 347058 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 347678 -1368
rect 347058 -1492 347678 -1424
rect 347058 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 347678 -1492
rect 347058 -1644 347678 -1548
rect 374058 40350 374678 53730
rect 374058 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 374678 40350
rect 374058 40226 374678 40294
rect 374058 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 374678 40226
rect 374058 40102 374678 40170
rect 374058 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 374678 40102
rect 374058 39978 374678 40046
rect 374058 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 374678 39978
rect 374058 22350 374678 39922
rect 374058 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 374678 22350
rect 374058 22226 374678 22294
rect 374058 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 374678 22226
rect 374058 22102 374678 22170
rect 374058 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 374678 22102
rect 374058 21978 374678 22046
rect 374058 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 374678 21978
rect 374058 4350 374678 21922
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 374058 4102 374678 4170
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 374058 -160 374678 3922
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 377778 46350 378398 53730
rect 377778 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 378398 46350
rect 377778 46226 378398 46294
rect 377778 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 378398 46226
rect 377778 46102 378398 46170
rect 377778 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 378398 46102
rect 377778 45978 378398 46046
rect 377778 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 378398 45978
rect 377778 28350 378398 45922
rect 377778 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 378398 28350
rect 377778 28226 378398 28294
rect 377778 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 378398 28226
rect 377778 28102 378398 28170
rect 377778 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 378398 28102
rect 377778 27978 378398 28046
rect 377778 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 378398 27978
rect 377778 10350 378398 27922
rect 377778 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 378398 10350
rect 377778 10226 378398 10294
rect 377778 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 378398 10226
rect 377778 10102 378398 10170
rect 377778 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 378398 10102
rect 377778 9978 378398 10046
rect 377778 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 378398 9978
rect 377778 -1120 378398 9922
rect 377778 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 378398 -1120
rect 377778 -1244 378398 -1176
rect 377778 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 378398 -1244
rect 377778 -1368 378398 -1300
rect 377778 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 378398 -1368
rect 377778 -1492 378398 -1424
rect 377778 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 378398 -1492
rect 377778 -1644 378398 -1548
rect 404778 40350 405398 53730
rect 404778 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 405398 40350
rect 404778 40226 405398 40294
rect 404778 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 405398 40226
rect 404778 40102 405398 40170
rect 404778 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 405398 40102
rect 404778 39978 405398 40046
rect 404778 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 405398 39978
rect 404778 22350 405398 39922
rect 404778 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 405398 22350
rect 404778 22226 405398 22294
rect 404778 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 405398 22226
rect 404778 22102 405398 22170
rect 404778 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 405398 22102
rect 404778 21978 405398 22046
rect 404778 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 405398 21978
rect 404778 4350 405398 21922
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 404778 4102 405398 4170
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 404778 -160 405398 3922
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 408498 46350 409118 53730
rect 408498 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 409118 46350
rect 408498 46226 409118 46294
rect 408498 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 409118 46226
rect 408498 46102 409118 46170
rect 408498 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 409118 46102
rect 408498 45978 409118 46046
rect 408498 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 409118 45978
rect 408498 28350 409118 45922
rect 408498 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 409118 28350
rect 408498 28226 409118 28294
rect 408498 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 409118 28226
rect 408498 28102 409118 28170
rect 408498 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 409118 28102
rect 408498 27978 409118 28046
rect 408498 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 409118 27978
rect 408498 10350 409118 27922
rect 408498 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 409118 10350
rect 408498 10226 409118 10294
rect 408498 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 409118 10226
rect 408498 10102 409118 10170
rect 408498 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 409118 10102
rect 408498 9978 409118 10046
rect 408498 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 409118 9978
rect 408498 -1120 409118 9922
rect 408498 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 409118 -1120
rect 408498 -1244 409118 -1176
rect 408498 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 409118 -1244
rect 408498 -1368 409118 -1300
rect 408498 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 409118 -1368
rect 408498 -1492 409118 -1424
rect 408498 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 409118 -1492
rect 408498 -1644 409118 -1548
rect 435498 40350 436118 57922
rect 435498 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 436118 40350
rect 435498 40226 436118 40294
rect 435498 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 436118 40226
rect 435498 40102 436118 40170
rect 435498 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 436118 40102
rect 435498 39978 436118 40046
rect 435498 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 436118 39978
rect 435498 22350 436118 39922
rect 435498 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 436118 22350
rect 435498 22226 436118 22294
rect 435498 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 436118 22226
rect 435498 22102 436118 22170
rect 435498 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 436118 22102
rect 435498 21978 436118 22046
rect 435498 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 436118 21978
rect 435498 4350 436118 21922
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 435498 4102 436118 4170
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 435498 -160 436118 3922
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 439218 172350 439838 173466
rect 439218 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 439838 172350
rect 439218 172226 439838 172294
rect 439218 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 439838 172226
rect 439218 172102 439838 172170
rect 439218 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 439838 172102
rect 439218 171978 439838 172046
rect 439218 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 439838 171978
rect 439218 154350 439838 171922
rect 469938 172350 470558 173466
rect 469938 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 470558 172350
rect 469938 172226 470558 172294
rect 469938 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 470558 172226
rect 469938 172102 470558 172170
rect 469938 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 470558 172102
rect 469938 171978 470558 172046
rect 469938 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 470558 171978
rect 439218 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 439838 154350
rect 439218 154226 439838 154294
rect 439218 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 439838 154226
rect 439218 154102 439838 154170
rect 439218 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 439838 154102
rect 439218 153978 439838 154046
rect 439218 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 439838 153978
rect 439218 136350 439838 153922
rect 439218 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 439838 136350
rect 439218 136226 439838 136294
rect 439218 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 439838 136226
rect 439218 136102 439838 136170
rect 439218 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 439838 136102
rect 439218 135978 439838 136046
rect 439218 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 439838 135978
rect 439218 118350 439838 135922
rect 457772 170772 457828 170782
rect 457660 131908 457716 131918
rect 457660 130564 457716 131852
rect 457660 130498 457716 130508
rect 457660 121940 457716 121950
rect 457660 118916 457716 121884
rect 457660 118850 457716 118860
rect 457660 118580 457716 118590
rect 439218 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 439838 118350
rect 439218 118226 439838 118294
rect 439218 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 439838 118226
rect 439218 118102 439838 118170
rect 439218 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 439838 118102
rect 439218 117978 439838 118046
rect 439218 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 439838 117978
rect 439218 100350 439838 117922
rect 457548 118468 457604 118478
rect 457548 114268 457604 118412
rect 457660 116900 457716 118524
rect 457660 116834 457716 116844
rect 457660 115892 457716 115902
rect 457660 115792 457716 115802
rect 457548 114212 457716 114268
rect 439218 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 439838 100350
rect 439218 100226 439838 100294
rect 439218 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 439838 100226
rect 439218 100102 439838 100170
rect 439218 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 439838 100102
rect 439218 99978 439838 100046
rect 439218 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 439838 99978
rect 439218 82350 439838 99922
rect 457660 95620 457716 114212
rect 457660 95554 457716 95564
rect 439218 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 439838 82350
rect 439218 82226 439838 82294
rect 439218 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 439838 82226
rect 439218 82102 439838 82170
rect 439218 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 439838 82102
rect 439218 81978 439838 82046
rect 439218 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 439838 81978
rect 439218 64350 439838 81922
rect 457772 81060 457828 170716
rect 457884 169316 457940 169326
rect 457884 83972 457940 169260
rect 457996 162484 458052 162494
rect 457996 148596 458052 162428
rect 469938 154350 470558 171922
rect 490588 173098 490644 173108
rect 469938 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 470558 154350
rect 469938 154226 470558 154294
rect 469938 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 470558 154226
rect 469938 154102 470558 154170
rect 469938 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 470558 154102
rect 469938 153978 470558 154046
rect 488908 168778 488964 168788
rect 488908 154084 488964 168722
rect 490588 154308 490644 173042
rect 500658 172350 501278 173466
rect 500658 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 501278 172350
rect 500658 172226 501278 172294
rect 500658 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 501278 172226
rect 500658 172102 501278 172170
rect 500658 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 501278 172102
rect 500658 171978 501278 172046
rect 500658 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 501278 171978
rect 490588 154242 490644 154252
rect 493164 157078 493220 157088
rect 488908 154018 488964 154028
rect 469938 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 470558 153978
rect 469938 149870 470558 153922
rect 493164 153300 493220 157022
rect 493164 153234 493220 153244
rect 500658 154350 501278 171922
rect 500658 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 501278 154350
rect 500658 154226 501278 154294
rect 500658 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 501278 154226
rect 500658 154102 501278 154170
rect 500658 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 501278 154102
rect 500658 153978 501278 154046
rect 500658 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 501278 153978
rect 482076 150598 482132 150608
rect 463372 149828 463428 149838
rect 457996 148530 458052 148540
rect 462028 149044 462084 149054
rect 462028 146098 462084 148988
rect 463372 147718 463428 149772
rect 482076 149716 482132 150542
rect 500658 149870 501278 153922
rect 531378 172350 531998 173466
rect 559468 173012 559524 398222
rect 559468 172946 559524 172956
rect 559580 395398 559636 395408
rect 559580 172676 559636 395342
rect 562098 388350 562718 405922
rect 565292 535780 565348 535790
rect 565292 404398 565348 535724
rect 568652 522564 568708 522574
rect 566972 482916 567028 482926
rect 566972 408178 567028 482860
rect 568652 411058 568708 522508
rect 568652 410992 568708 411002
rect 570332 456484 570388 456494
rect 566972 408112 567028 408122
rect 565292 404332 565348 404342
rect 570332 404218 570388 456428
rect 584668 409438 584724 590156
rect 589098 580350 589718 596784
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 589098 562350 589718 579922
rect 590492 588644 590548 588654
rect 590492 575540 590548 588588
rect 590492 575474 590548 575484
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 584668 409372 584724 409382
rect 585452 562212 585508 562222
rect 585452 409078 585508 562156
rect 585452 409012 585508 409022
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 589098 544350 589718 561922
rect 590492 567924 590548 567934
rect 590492 549220 590548 567868
rect 590492 549154 590548 549164
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 589098 526350 589718 543922
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 589098 508350 589718 525922
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 589098 472350 589718 489922
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 589098 454350 589718 471922
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 589098 436350 589718 453922
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 589098 418350 589718 435922
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 570332 404152 570388 404162
rect 572012 402058 572068 402068
rect 562098 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 562718 388350
rect 562098 388226 562718 388294
rect 562098 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 562718 388226
rect 562098 388102 562718 388170
rect 562098 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 562718 388102
rect 562098 387978 562718 388046
rect 562098 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 562718 387978
rect 562098 370350 562718 387922
rect 562098 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 562718 370350
rect 562098 370226 562718 370294
rect 562098 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 562718 370226
rect 562098 370102 562718 370170
rect 562098 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 562718 370102
rect 562098 369978 562718 370046
rect 562098 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 562718 369978
rect 562098 352350 562718 369922
rect 562098 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 562718 352350
rect 562098 352226 562718 352294
rect 562098 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 562718 352226
rect 562098 352102 562718 352170
rect 562098 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 562718 352102
rect 562098 351978 562718 352046
rect 562098 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 562718 351978
rect 562098 334350 562718 351922
rect 562098 334294 562194 334350
rect 562250 334294 562318 334350
rect 562374 334294 562442 334350
rect 562498 334294 562566 334350
rect 562622 334294 562718 334350
rect 562098 334226 562718 334294
rect 562098 334170 562194 334226
rect 562250 334170 562318 334226
rect 562374 334170 562442 334226
rect 562498 334170 562566 334226
rect 562622 334170 562718 334226
rect 562098 334102 562718 334170
rect 562098 334046 562194 334102
rect 562250 334046 562318 334102
rect 562374 334046 562442 334102
rect 562498 334046 562566 334102
rect 562622 334046 562718 334102
rect 562098 333978 562718 334046
rect 562098 333922 562194 333978
rect 562250 333922 562318 333978
rect 562374 333922 562442 333978
rect 562498 333922 562566 333978
rect 562622 333922 562718 333978
rect 562098 316350 562718 333922
rect 562098 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 562718 316350
rect 562098 316226 562718 316294
rect 562098 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 562718 316226
rect 562098 316102 562718 316170
rect 562098 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 562718 316102
rect 562098 315978 562718 316046
rect 562098 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 562718 315978
rect 562098 298350 562718 315922
rect 562098 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 562718 298350
rect 562098 298226 562718 298294
rect 562098 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 562718 298226
rect 562098 298102 562718 298170
rect 562098 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 562718 298102
rect 562098 297978 562718 298046
rect 562098 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 562718 297978
rect 562098 280350 562718 297922
rect 562098 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 562718 280350
rect 562098 280226 562718 280294
rect 562098 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 562718 280226
rect 562098 280102 562718 280170
rect 562098 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 562718 280102
rect 562098 279978 562718 280046
rect 562098 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 562718 279978
rect 562098 262350 562718 279922
rect 562098 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 562718 262350
rect 562098 262226 562718 262294
rect 562098 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 562718 262226
rect 562098 262102 562718 262170
rect 562098 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 562718 262102
rect 562098 261978 562718 262046
rect 562098 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 562718 261978
rect 562098 244350 562718 261922
rect 562098 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 562718 244350
rect 562098 244226 562718 244294
rect 562098 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 562718 244226
rect 562098 244102 562718 244170
rect 562098 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 562718 244102
rect 562098 243978 562718 244046
rect 562098 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 562718 243978
rect 562098 226350 562718 243922
rect 562098 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 562718 226350
rect 562098 226226 562718 226294
rect 562098 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 562718 226226
rect 562098 226102 562718 226170
rect 562098 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 562718 226102
rect 562098 225978 562718 226046
rect 562098 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 562718 225978
rect 562098 208350 562718 225922
rect 562098 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 562718 208350
rect 562098 208226 562718 208294
rect 562098 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 562718 208226
rect 562098 208102 562718 208170
rect 562098 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 562718 208102
rect 562098 207978 562718 208046
rect 562098 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 562718 207978
rect 562098 190350 562718 207922
rect 562098 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 562718 190350
rect 562098 190226 562718 190294
rect 562098 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 562718 190226
rect 562098 190102 562718 190170
rect 562098 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 562718 190102
rect 562098 189978 562718 190046
rect 562098 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 562718 189978
rect 559580 172610 559636 172620
rect 561148 173818 561204 173828
rect 531378 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 531998 172350
rect 531378 172226 531998 172294
rect 531378 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 531998 172226
rect 531378 172102 531998 172170
rect 531378 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 531998 172102
rect 531378 171978 531998 172046
rect 531378 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 531998 171978
rect 531378 154350 531998 171922
rect 531378 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 531998 154350
rect 531378 154226 531998 154294
rect 531378 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 531998 154226
rect 531378 154102 531998 154170
rect 531378 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 531998 154102
rect 531378 153978 531998 154046
rect 531378 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 531998 153978
rect 502572 153658 502628 153668
rect 502572 152964 502628 153602
rect 502572 152898 502628 152908
rect 503132 153478 503188 153488
rect 503132 152964 503188 153422
rect 503132 152898 503188 152908
rect 506828 150276 506884 150286
rect 482076 149650 482132 149660
rect 501004 149158 501060 149166
rect 501452 149158 501508 149166
rect 501004 149156 501508 149158
rect 501060 149102 501452 149156
rect 501004 149090 501060 149100
rect 501452 149090 501508 149100
rect 506828 149156 506884 150220
rect 531378 149870 531998 153922
rect 559468 172228 559524 172238
rect 506828 149090 506884 149100
rect 463372 147652 463428 147662
rect 462028 146032 462084 146042
rect 479808 136350 480128 136384
rect 479808 136294 479878 136350
rect 479934 136294 480002 136350
rect 480058 136294 480128 136350
rect 479808 136226 480128 136294
rect 479808 136170 479878 136226
rect 479934 136170 480002 136226
rect 480058 136170 480128 136226
rect 479808 136102 480128 136170
rect 479808 136046 479878 136102
rect 479934 136046 480002 136102
rect 480058 136046 480128 136102
rect 479808 135978 480128 136046
rect 479808 135922 479878 135978
rect 479934 135922 480002 135978
rect 480058 135922 480128 135978
rect 479808 135888 480128 135922
rect 510528 136350 510848 136384
rect 510528 136294 510598 136350
rect 510654 136294 510722 136350
rect 510778 136294 510848 136350
rect 510528 136226 510848 136294
rect 510528 136170 510598 136226
rect 510654 136170 510722 136226
rect 510778 136170 510848 136226
rect 510528 136102 510848 136170
rect 510528 136046 510598 136102
rect 510654 136046 510722 136102
rect 510778 136046 510848 136102
rect 510528 135978 510848 136046
rect 510528 135922 510598 135978
rect 510654 135922 510722 135978
rect 510778 135922 510848 135978
rect 510528 135888 510848 135922
rect 541248 136350 541568 136384
rect 541248 136294 541318 136350
rect 541374 136294 541442 136350
rect 541498 136294 541568 136350
rect 541248 136226 541568 136294
rect 541248 136170 541318 136226
rect 541374 136170 541442 136226
rect 541498 136170 541568 136226
rect 541248 136102 541568 136170
rect 541248 136046 541318 136102
rect 541374 136046 541442 136102
rect 541498 136046 541568 136102
rect 541248 135978 541568 136046
rect 541248 135922 541318 135978
rect 541374 135922 541442 135978
rect 541498 135922 541568 135978
rect 541248 135888 541568 135922
rect 464448 130350 464768 130384
rect 464448 130294 464518 130350
rect 464574 130294 464642 130350
rect 464698 130294 464768 130350
rect 464448 130226 464768 130294
rect 464448 130170 464518 130226
rect 464574 130170 464642 130226
rect 464698 130170 464768 130226
rect 464448 130102 464768 130170
rect 464448 130046 464518 130102
rect 464574 130046 464642 130102
rect 464698 130046 464768 130102
rect 464448 129978 464768 130046
rect 464448 129922 464518 129978
rect 464574 129922 464642 129978
rect 464698 129922 464768 129978
rect 464448 129888 464768 129922
rect 495168 130350 495488 130384
rect 495168 130294 495238 130350
rect 495294 130294 495362 130350
rect 495418 130294 495488 130350
rect 495168 130226 495488 130294
rect 495168 130170 495238 130226
rect 495294 130170 495362 130226
rect 495418 130170 495488 130226
rect 495168 130102 495488 130170
rect 495168 130046 495238 130102
rect 495294 130046 495362 130102
rect 495418 130046 495488 130102
rect 495168 129978 495488 130046
rect 495168 129922 495238 129978
rect 495294 129922 495362 129978
rect 495418 129922 495488 129978
rect 495168 129888 495488 129922
rect 525888 130350 526208 130384
rect 525888 130294 525958 130350
rect 526014 130294 526082 130350
rect 526138 130294 526208 130350
rect 525888 130226 526208 130294
rect 525888 130170 525958 130226
rect 526014 130170 526082 130226
rect 526138 130170 526208 130226
rect 525888 130102 526208 130170
rect 525888 130046 525958 130102
rect 526014 130046 526082 130102
rect 526138 130046 526208 130102
rect 525888 129978 526208 130046
rect 525888 129922 525958 129978
rect 526014 129922 526082 129978
rect 526138 129922 526208 129978
rect 525888 129888 526208 129922
rect 556608 130350 556928 130384
rect 556608 130294 556678 130350
rect 556734 130294 556802 130350
rect 556858 130294 556928 130350
rect 556608 130226 556928 130294
rect 556608 130170 556678 130226
rect 556734 130170 556802 130226
rect 556858 130170 556928 130226
rect 556608 130102 556928 130170
rect 556608 130046 556678 130102
rect 556734 130046 556802 130102
rect 556858 130046 556928 130102
rect 556608 129978 556928 130046
rect 556608 129922 556678 129978
rect 556734 129922 556802 129978
rect 556858 129922 556928 129978
rect 556608 129888 556928 129922
rect 458108 128548 458164 128558
rect 457884 83906 457940 83916
rect 457996 126868 458052 126878
rect 457772 80994 457828 81004
rect 457996 72212 458052 126812
rect 458108 75236 458164 128492
rect 458220 126980 458276 126990
rect 458220 78148 458276 126924
rect 458332 120148 458388 120158
rect 458332 117298 458388 120092
rect 458556 118692 458612 118702
rect 458556 117572 458612 118636
rect 479808 118350 480128 118384
rect 479808 118294 479878 118350
rect 479934 118294 480002 118350
rect 480058 118294 480128 118350
rect 479808 118226 480128 118294
rect 479808 118170 479878 118226
rect 479934 118170 480002 118226
rect 480058 118170 480128 118226
rect 479808 118102 480128 118170
rect 479808 118046 479878 118102
rect 479934 118046 480002 118102
rect 480058 118046 480128 118102
rect 479808 117978 480128 118046
rect 479808 117922 479878 117978
rect 479934 117922 480002 117978
rect 480058 117922 480128 117978
rect 479808 117888 480128 117922
rect 510528 118350 510848 118384
rect 510528 118294 510598 118350
rect 510654 118294 510722 118350
rect 510778 118294 510848 118350
rect 510528 118226 510848 118294
rect 510528 118170 510598 118226
rect 510654 118170 510722 118226
rect 510778 118170 510848 118226
rect 510528 118102 510848 118170
rect 510528 118046 510598 118102
rect 510654 118046 510722 118102
rect 510778 118046 510848 118102
rect 510528 117978 510848 118046
rect 510528 117922 510598 117978
rect 510654 117922 510722 117978
rect 510778 117922 510848 117978
rect 510528 117888 510848 117922
rect 541248 118350 541568 118384
rect 541248 118294 541318 118350
rect 541374 118294 541442 118350
rect 541498 118294 541568 118350
rect 541248 118226 541568 118294
rect 541248 118170 541318 118226
rect 541374 118170 541442 118226
rect 541498 118170 541568 118226
rect 541248 118102 541568 118170
rect 541248 118046 541318 118102
rect 541374 118046 541442 118102
rect 541498 118046 541568 118102
rect 541248 117978 541568 118046
rect 541248 117922 541318 117978
rect 541374 117922 541442 117978
rect 541498 117922 541568 117978
rect 541248 117888 541568 117922
rect 458556 117506 458612 117516
rect 458332 117242 458612 117298
rect 458332 117124 458388 117134
rect 458332 86884 458388 117068
rect 458444 116900 458500 116910
rect 458444 89796 458500 116844
rect 458556 98532 458612 117242
rect 464448 112350 464768 112384
rect 464448 112294 464518 112350
rect 464574 112294 464642 112350
rect 464698 112294 464768 112350
rect 464448 112226 464768 112294
rect 464448 112170 464518 112226
rect 464574 112170 464642 112226
rect 464698 112170 464768 112226
rect 464448 112102 464768 112170
rect 464448 112046 464518 112102
rect 464574 112046 464642 112102
rect 464698 112046 464768 112102
rect 464448 111978 464768 112046
rect 464448 111922 464518 111978
rect 464574 111922 464642 111978
rect 464698 111922 464768 111978
rect 464448 111888 464768 111922
rect 495168 112350 495488 112384
rect 495168 112294 495238 112350
rect 495294 112294 495362 112350
rect 495418 112294 495488 112350
rect 495168 112226 495488 112294
rect 495168 112170 495238 112226
rect 495294 112170 495362 112226
rect 495418 112170 495488 112226
rect 495168 112102 495488 112170
rect 495168 112046 495238 112102
rect 495294 112046 495362 112102
rect 495418 112046 495488 112102
rect 495168 111978 495488 112046
rect 495168 111922 495238 111978
rect 495294 111922 495362 111978
rect 495418 111922 495488 111978
rect 495168 111888 495488 111922
rect 525888 112350 526208 112384
rect 525888 112294 525958 112350
rect 526014 112294 526082 112350
rect 526138 112294 526208 112350
rect 525888 112226 526208 112294
rect 525888 112170 525958 112226
rect 526014 112170 526082 112226
rect 526138 112170 526208 112226
rect 525888 112102 526208 112170
rect 525888 112046 525958 112102
rect 526014 112046 526082 112102
rect 526138 112046 526208 112102
rect 525888 111978 526208 112046
rect 525888 111922 525958 111978
rect 526014 111922 526082 111978
rect 526138 111922 526208 111978
rect 525888 111888 526208 111922
rect 556608 112350 556928 112384
rect 556608 112294 556678 112350
rect 556734 112294 556802 112350
rect 556858 112294 556928 112350
rect 556608 112226 556928 112294
rect 556608 112170 556678 112226
rect 556734 112170 556802 112226
rect 556858 112170 556928 112226
rect 556608 112102 556928 112170
rect 556608 112046 556678 112102
rect 556734 112046 556802 112102
rect 556858 112046 556928 112102
rect 556608 111978 556928 112046
rect 556608 111922 556678 111978
rect 556734 111922 556802 111978
rect 556858 111922 556928 111978
rect 556608 111888 556928 111922
rect 479808 100350 480128 100384
rect 479808 100294 479878 100350
rect 479934 100294 480002 100350
rect 480058 100294 480128 100350
rect 479808 100226 480128 100294
rect 479808 100170 479878 100226
rect 479934 100170 480002 100226
rect 480058 100170 480128 100226
rect 479808 100102 480128 100170
rect 479808 100046 479878 100102
rect 479934 100046 480002 100102
rect 480058 100046 480128 100102
rect 479808 99978 480128 100046
rect 479808 99922 479878 99978
rect 479934 99922 480002 99978
rect 480058 99922 480128 99978
rect 479808 99888 480128 99922
rect 510528 100350 510848 100384
rect 510528 100294 510598 100350
rect 510654 100294 510722 100350
rect 510778 100294 510848 100350
rect 510528 100226 510848 100294
rect 510528 100170 510598 100226
rect 510654 100170 510722 100226
rect 510778 100170 510848 100226
rect 510528 100102 510848 100170
rect 510528 100046 510598 100102
rect 510654 100046 510722 100102
rect 510778 100046 510848 100102
rect 510528 99978 510848 100046
rect 510528 99922 510598 99978
rect 510654 99922 510722 99978
rect 510778 99922 510848 99978
rect 510528 99888 510848 99922
rect 541248 100350 541568 100384
rect 541248 100294 541318 100350
rect 541374 100294 541442 100350
rect 541498 100294 541568 100350
rect 541248 100226 541568 100294
rect 541248 100170 541318 100226
rect 541374 100170 541442 100226
rect 541498 100170 541568 100226
rect 541248 100102 541568 100170
rect 541248 100046 541318 100102
rect 541374 100046 541442 100102
rect 541498 100046 541568 100102
rect 541248 99978 541568 100046
rect 541248 99922 541318 99978
rect 541374 99922 541442 99978
rect 541498 99922 541568 99978
rect 541248 99888 541568 99922
rect 458556 98466 458612 98476
rect 464448 94350 464768 94384
rect 464448 94294 464518 94350
rect 464574 94294 464642 94350
rect 464698 94294 464768 94350
rect 464448 94226 464768 94294
rect 464448 94170 464518 94226
rect 464574 94170 464642 94226
rect 464698 94170 464768 94226
rect 464448 94102 464768 94170
rect 464448 94046 464518 94102
rect 464574 94046 464642 94102
rect 464698 94046 464768 94102
rect 464448 93978 464768 94046
rect 464448 93922 464518 93978
rect 464574 93922 464642 93978
rect 464698 93922 464768 93978
rect 464448 93888 464768 93922
rect 495168 94350 495488 94384
rect 495168 94294 495238 94350
rect 495294 94294 495362 94350
rect 495418 94294 495488 94350
rect 495168 94226 495488 94294
rect 495168 94170 495238 94226
rect 495294 94170 495362 94226
rect 495418 94170 495488 94226
rect 495168 94102 495488 94170
rect 495168 94046 495238 94102
rect 495294 94046 495362 94102
rect 495418 94046 495488 94102
rect 495168 93978 495488 94046
rect 495168 93922 495238 93978
rect 495294 93922 495362 93978
rect 495418 93922 495488 93978
rect 495168 93888 495488 93922
rect 525888 94350 526208 94384
rect 525888 94294 525958 94350
rect 526014 94294 526082 94350
rect 526138 94294 526208 94350
rect 525888 94226 526208 94294
rect 525888 94170 525958 94226
rect 526014 94170 526082 94226
rect 526138 94170 526208 94226
rect 525888 94102 526208 94170
rect 525888 94046 525958 94102
rect 526014 94046 526082 94102
rect 526138 94046 526208 94102
rect 525888 93978 526208 94046
rect 525888 93922 525958 93978
rect 526014 93922 526082 93978
rect 526138 93922 526208 93978
rect 525888 93888 526208 93922
rect 556608 94350 556928 94384
rect 556608 94294 556678 94350
rect 556734 94294 556802 94350
rect 556858 94294 556928 94350
rect 556608 94226 556928 94294
rect 556608 94170 556678 94226
rect 556734 94170 556802 94226
rect 556858 94170 556928 94226
rect 556608 94102 556928 94170
rect 556608 94046 556678 94102
rect 556734 94046 556802 94102
rect 556858 94046 556928 94102
rect 556608 93978 556928 94046
rect 556608 93922 556678 93978
rect 556734 93922 556802 93978
rect 556858 93922 556928 93978
rect 556608 93888 556928 93922
rect 458444 89730 458500 89740
rect 458332 86818 458388 86828
rect 479808 82350 480128 82384
rect 479808 82294 479878 82350
rect 479934 82294 480002 82350
rect 480058 82294 480128 82350
rect 479808 82226 480128 82294
rect 479808 82170 479878 82226
rect 479934 82170 480002 82226
rect 480058 82170 480128 82226
rect 479808 82102 480128 82170
rect 479808 82046 479878 82102
rect 479934 82046 480002 82102
rect 480058 82046 480128 82102
rect 479808 81978 480128 82046
rect 479808 81922 479878 81978
rect 479934 81922 480002 81978
rect 480058 81922 480128 81978
rect 479808 81888 480128 81922
rect 510528 82350 510848 82384
rect 510528 82294 510598 82350
rect 510654 82294 510722 82350
rect 510778 82294 510848 82350
rect 510528 82226 510848 82294
rect 510528 82170 510598 82226
rect 510654 82170 510722 82226
rect 510778 82170 510848 82226
rect 510528 82102 510848 82170
rect 510528 82046 510598 82102
rect 510654 82046 510722 82102
rect 510778 82046 510848 82102
rect 510528 81978 510848 82046
rect 510528 81922 510598 81978
rect 510654 81922 510722 81978
rect 510778 81922 510848 81978
rect 510528 81888 510848 81922
rect 541248 82350 541568 82384
rect 541248 82294 541318 82350
rect 541374 82294 541442 82350
rect 541498 82294 541568 82350
rect 541248 82226 541568 82294
rect 541248 82170 541318 82226
rect 541374 82170 541442 82226
rect 541498 82170 541568 82226
rect 541248 82102 541568 82170
rect 541248 82046 541318 82102
rect 541374 82046 541442 82102
rect 541498 82046 541568 82102
rect 541248 81978 541568 82046
rect 541248 81922 541318 81978
rect 541374 81922 541442 81978
rect 541498 81922 541568 81978
rect 541248 81888 541568 81922
rect 458220 78082 458276 78092
rect 464448 76350 464768 76384
rect 464448 76294 464518 76350
rect 464574 76294 464642 76350
rect 464698 76294 464768 76350
rect 464448 76226 464768 76294
rect 464448 76170 464518 76226
rect 464574 76170 464642 76226
rect 464698 76170 464768 76226
rect 464448 76102 464768 76170
rect 464448 76046 464518 76102
rect 464574 76046 464642 76102
rect 464698 76046 464768 76102
rect 464448 75978 464768 76046
rect 464448 75922 464518 75978
rect 464574 75922 464642 75978
rect 464698 75922 464768 75978
rect 464448 75888 464768 75922
rect 495168 76350 495488 76384
rect 495168 76294 495238 76350
rect 495294 76294 495362 76350
rect 495418 76294 495488 76350
rect 495168 76226 495488 76294
rect 495168 76170 495238 76226
rect 495294 76170 495362 76226
rect 495418 76170 495488 76226
rect 495168 76102 495488 76170
rect 495168 76046 495238 76102
rect 495294 76046 495362 76102
rect 495418 76046 495488 76102
rect 495168 75978 495488 76046
rect 495168 75922 495238 75978
rect 495294 75922 495362 75978
rect 495418 75922 495488 75978
rect 495168 75888 495488 75922
rect 525888 76350 526208 76384
rect 525888 76294 525958 76350
rect 526014 76294 526082 76350
rect 526138 76294 526208 76350
rect 525888 76226 526208 76294
rect 525888 76170 525958 76226
rect 526014 76170 526082 76226
rect 526138 76170 526208 76226
rect 525888 76102 526208 76170
rect 525888 76046 525958 76102
rect 526014 76046 526082 76102
rect 526138 76046 526208 76102
rect 525888 75978 526208 76046
rect 525888 75922 525958 75978
rect 526014 75922 526082 75978
rect 526138 75922 526208 75978
rect 525888 75888 526208 75922
rect 556608 76350 556928 76384
rect 556608 76294 556678 76350
rect 556734 76294 556802 76350
rect 556858 76294 556928 76350
rect 556608 76226 556928 76294
rect 556608 76170 556678 76226
rect 556734 76170 556802 76226
rect 556858 76170 556928 76226
rect 556608 76102 556928 76170
rect 556608 76046 556678 76102
rect 556734 76046 556802 76102
rect 556858 76046 556928 76102
rect 556608 75978 556928 76046
rect 556608 75922 556678 75978
rect 556734 75922 556802 75978
rect 556858 75922 556928 75978
rect 556608 75888 556928 75922
rect 559468 75572 559524 172172
rect 559580 170578 559636 170588
rect 559580 78708 559636 170522
rect 559804 168980 559860 168990
rect 559580 78642 559636 78652
rect 559692 163940 559748 163950
rect 559692 77140 559748 163884
rect 559804 89684 559860 168924
rect 559916 167188 559972 167198
rect 559916 95956 559972 167132
rect 561148 105364 561204 173762
rect 562098 172350 562718 189922
rect 570332 393598 570388 393608
rect 570332 178948 570388 393542
rect 570332 178882 570388 178892
rect 562098 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 562718 172350
rect 562098 172226 562718 172294
rect 562098 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 562718 172226
rect 562098 172102 562718 172170
rect 562098 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 562718 172102
rect 562098 171978 562718 172046
rect 562098 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 562718 171978
rect 561260 158878 561316 158888
rect 561260 125748 561316 158822
rect 561260 125682 561316 125692
rect 562098 154350 562718 171922
rect 563164 168868 563220 168878
rect 562098 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 562718 154350
rect 562098 154226 562718 154294
rect 562098 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 562718 154226
rect 562098 154102 562718 154170
rect 562098 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 562718 154102
rect 562098 153978 562718 154046
rect 562098 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 562718 153978
rect 562098 136350 562718 153922
rect 562098 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 562718 136350
rect 562098 136226 562718 136294
rect 562098 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 562718 136226
rect 562098 136102 562718 136170
rect 562098 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 562718 136102
rect 562098 135978 562718 136046
rect 562098 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 562718 135978
rect 561148 105298 561204 105308
rect 562098 118350 562718 135922
rect 562098 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 562718 118350
rect 562098 118226 562718 118294
rect 562098 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 562718 118226
rect 562098 118102 562718 118170
rect 562098 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 562718 118102
rect 562098 117978 562718 118046
rect 562098 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 562718 117978
rect 559916 95890 559972 95900
rect 562098 100350 562718 117922
rect 562098 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 562718 100350
rect 562098 100226 562718 100294
rect 562098 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 562718 100226
rect 562098 100102 562718 100170
rect 562098 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 562718 100102
rect 562098 99978 562718 100046
rect 562098 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 562718 99978
rect 559804 89618 559860 89628
rect 559692 77074 559748 77084
rect 559804 84980 559860 84990
rect 559468 75506 559524 75516
rect 458108 75170 458164 75180
rect 457996 72146 458052 72156
rect 457772 69300 457828 69310
rect 439218 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 439838 64350
rect 439218 64226 439838 64294
rect 439218 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 439838 64226
rect 439218 64102 439838 64170
rect 439218 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 439838 64102
rect 439218 63978 439838 64046
rect 439218 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 439838 63978
rect 439218 46350 439838 63922
rect 457660 66388 457716 66398
rect 457660 57764 457716 66332
rect 457660 57698 457716 57708
rect 457660 54740 457716 54750
rect 457660 52052 457716 54684
rect 457772 52724 457828 69244
rect 457772 52658 457828 52668
rect 457884 66388 457940 66398
rect 457660 51986 457716 51996
rect 457884 51492 457940 66332
rect 479808 64350 480128 64384
rect 479808 64294 479878 64350
rect 479934 64294 480002 64350
rect 480058 64294 480128 64350
rect 479808 64226 480128 64294
rect 479808 64170 479878 64226
rect 479934 64170 480002 64226
rect 480058 64170 480128 64226
rect 479808 64102 480128 64170
rect 479808 64046 479878 64102
rect 479934 64046 480002 64102
rect 480058 64046 480128 64102
rect 479808 63978 480128 64046
rect 479808 63922 479878 63978
rect 479934 63922 480002 63978
rect 480058 63922 480128 63978
rect 479808 63888 480128 63922
rect 510528 64350 510848 64384
rect 510528 64294 510598 64350
rect 510654 64294 510722 64350
rect 510778 64294 510848 64350
rect 510528 64226 510848 64294
rect 510528 64170 510598 64226
rect 510654 64170 510722 64226
rect 510778 64170 510848 64226
rect 510528 64102 510848 64170
rect 510528 64046 510598 64102
rect 510654 64046 510722 64102
rect 510778 64046 510848 64102
rect 510528 63978 510848 64046
rect 510528 63922 510598 63978
rect 510654 63922 510722 63978
rect 510778 63922 510848 63978
rect 510528 63888 510848 63922
rect 541248 64350 541568 64384
rect 541248 64294 541318 64350
rect 541374 64294 541442 64350
rect 541498 64294 541568 64350
rect 541248 64226 541568 64294
rect 541248 64170 541318 64226
rect 541374 64170 541442 64226
rect 541498 64170 541568 64226
rect 541248 64102 541568 64170
rect 541248 64046 541318 64102
rect 541374 64046 541442 64102
rect 541498 64046 541568 64102
rect 541248 63978 541568 64046
rect 541248 63922 541318 63978
rect 541374 63922 541442 63978
rect 541498 63922 541568 63978
rect 541248 63888 541568 63922
rect 457996 63476 458052 63486
rect 457996 52948 458052 63420
rect 464448 58350 464768 58384
rect 464448 58294 464518 58350
rect 464574 58294 464642 58350
rect 464698 58294 464768 58350
rect 464448 58226 464768 58294
rect 464448 58170 464518 58226
rect 464574 58170 464642 58226
rect 464698 58170 464768 58226
rect 464448 58102 464768 58170
rect 464448 58046 464518 58102
rect 464574 58046 464642 58102
rect 464698 58046 464768 58102
rect 464448 57978 464768 58046
rect 464448 57922 464518 57978
rect 464574 57922 464642 57978
rect 464698 57922 464768 57978
rect 464448 57888 464768 57922
rect 495168 58350 495488 58384
rect 495168 58294 495238 58350
rect 495294 58294 495362 58350
rect 495418 58294 495488 58350
rect 495168 58226 495488 58294
rect 495168 58170 495238 58226
rect 495294 58170 495362 58226
rect 495418 58170 495488 58226
rect 495168 58102 495488 58170
rect 495168 58046 495238 58102
rect 495294 58046 495362 58102
rect 495418 58046 495488 58102
rect 495168 57978 495488 58046
rect 495168 57922 495238 57978
rect 495294 57922 495362 57978
rect 495418 57922 495488 57978
rect 495168 57888 495488 57922
rect 525888 58350 526208 58384
rect 525888 58294 525958 58350
rect 526014 58294 526082 58350
rect 526138 58294 526208 58350
rect 525888 58226 526208 58294
rect 525888 58170 525958 58226
rect 526014 58170 526082 58226
rect 526138 58170 526208 58226
rect 525888 58102 526208 58170
rect 525888 58046 525958 58102
rect 526014 58046 526082 58102
rect 526138 58046 526208 58102
rect 525888 57978 526208 58046
rect 525888 57922 525958 57978
rect 526014 57922 526082 57978
rect 526138 57922 526208 57978
rect 525888 57888 526208 57922
rect 556608 58350 556928 58384
rect 556608 58294 556678 58350
rect 556734 58294 556802 58350
rect 556858 58294 556928 58350
rect 556608 58226 556928 58294
rect 556608 58170 556678 58226
rect 556734 58170 556802 58226
rect 556858 58170 556928 58226
rect 556608 58102 556928 58170
rect 556608 58046 556678 58102
rect 556734 58046 556802 58102
rect 556858 58046 556928 58102
rect 556608 57978 556928 58046
rect 556608 57922 556678 57978
rect 556734 57922 556802 57978
rect 556858 57922 556928 57978
rect 556608 57888 556928 57922
rect 457996 52882 458052 52892
rect 559468 56084 559524 56094
rect 457884 51426 457940 51436
rect 559468 50260 559524 56028
rect 559468 50194 559524 50204
rect 439218 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 439838 46350
rect 439218 46226 439838 46294
rect 439218 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 439838 46226
rect 439218 46102 439838 46170
rect 439218 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 439838 46102
rect 439218 45978 439838 46046
rect 439218 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 439838 45978
rect 439218 28350 439838 45922
rect 439218 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 439838 28350
rect 439218 28226 439838 28294
rect 439218 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 439838 28226
rect 439218 28102 439838 28170
rect 439218 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 439838 28102
rect 439218 27978 439838 28046
rect 439218 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 439838 27978
rect 439218 10350 439838 27922
rect 439218 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 439838 10350
rect 439218 10226 439838 10294
rect 439218 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 439838 10226
rect 439218 10102 439838 10170
rect 439218 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 439838 10102
rect 439218 9978 439838 10046
rect 439218 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 439838 9978
rect 439218 -1120 439838 9922
rect 439218 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 439838 -1120
rect 439218 -1244 439838 -1176
rect 439218 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 439838 -1244
rect 439218 -1368 439838 -1300
rect 439218 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 439838 -1368
rect 439218 -1492 439838 -1424
rect 439218 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 439838 -1492
rect 439218 -1644 439838 -1548
rect 466218 40350 466838 48690
rect 466218 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 466838 40350
rect 466218 40226 466838 40294
rect 466218 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 466838 40226
rect 466218 40102 466838 40170
rect 466218 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 466838 40102
rect 466218 39978 466838 40046
rect 466218 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 466838 39978
rect 466218 22350 466838 39922
rect 466218 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 466838 22350
rect 466218 22226 466838 22294
rect 466218 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 466838 22226
rect 466218 22102 466838 22170
rect 466218 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 466838 22102
rect 466218 21978 466838 22046
rect 466218 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 466838 21978
rect 466218 4350 466838 21922
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 466218 -160 466838 3922
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 469938 46350 470558 48690
rect 469938 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 470558 46350
rect 469938 46226 470558 46294
rect 469938 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 470558 46226
rect 469938 46102 470558 46170
rect 469938 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 470558 46102
rect 469938 45978 470558 46046
rect 469938 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 470558 45978
rect 469938 28350 470558 45922
rect 469938 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 470558 28350
rect 469938 28226 470558 28294
rect 469938 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 470558 28226
rect 469938 28102 470558 28170
rect 469938 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 470558 28102
rect 469938 27978 470558 28046
rect 469938 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 470558 27978
rect 469938 10350 470558 27922
rect 469938 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 470558 10350
rect 469938 10226 470558 10294
rect 469938 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 470558 10226
rect 469938 10102 470558 10170
rect 469938 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 470558 10102
rect 469938 9978 470558 10046
rect 469938 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 470558 9978
rect 469938 -1120 470558 9922
rect 469938 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 470558 -1120
rect 469938 -1244 470558 -1176
rect 469938 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 470558 -1244
rect 469938 -1368 470558 -1300
rect 469938 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 470558 -1368
rect 469938 -1492 470558 -1424
rect 469938 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 470558 -1492
rect 469938 -1644 470558 -1548
rect 496938 40350 497558 48690
rect 496938 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 497558 40350
rect 496938 40226 497558 40294
rect 496938 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 497558 40226
rect 496938 40102 497558 40170
rect 496938 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 497558 40102
rect 496938 39978 497558 40046
rect 496938 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 497558 39978
rect 496938 22350 497558 39922
rect 496938 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 497558 22350
rect 496938 22226 497558 22294
rect 496938 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 497558 22226
rect 496938 22102 497558 22170
rect 496938 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 497558 22102
rect 496938 21978 497558 22046
rect 496938 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 497558 21978
rect 496938 4350 497558 21922
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 496938 4102 497558 4170
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 496938 -160 497558 3922
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 500658 46350 501278 48690
rect 500658 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 501278 46350
rect 500658 46226 501278 46294
rect 500658 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 501278 46226
rect 500658 46102 501278 46170
rect 500658 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 501278 46102
rect 500658 45978 501278 46046
rect 500658 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 501278 45978
rect 500658 28350 501278 45922
rect 500658 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 501278 28350
rect 500658 28226 501278 28294
rect 500658 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 501278 28226
rect 500658 28102 501278 28170
rect 500658 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 501278 28102
rect 500658 27978 501278 28046
rect 500658 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 501278 27978
rect 500658 10350 501278 27922
rect 500658 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 501278 10350
rect 500658 10226 501278 10294
rect 500658 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 501278 10226
rect 500658 10102 501278 10170
rect 500658 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 501278 10102
rect 500658 9978 501278 10046
rect 500658 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 501278 9978
rect 500658 -1120 501278 9922
rect 500658 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 501278 -1120
rect 500658 -1244 501278 -1176
rect 500658 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 501278 -1244
rect 500658 -1368 501278 -1300
rect 500658 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 501278 -1368
rect 500658 -1492 501278 -1424
rect 500658 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 501278 -1492
rect 500658 -1644 501278 -1548
rect 527658 40350 528278 48690
rect 527658 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 528278 40350
rect 527658 40226 528278 40294
rect 527658 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 528278 40226
rect 527658 40102 528278 40170
rect 527658 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 528278 40102
rect 527658 39978 528278 40046
rect 527658 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 528278 39978
rect 527658 22350 528278 39922
rect 527658 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 528278 22350
rect 527658 22226 528278 22294
rect 527658 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 528278 22226
rect 527658 22102 528278 22170
rect 527658 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 528278 22102
rect 527658 21978 528278 22046
rect 527658 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 528278 21978
rect 527658 4350 528278 21922
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 527658 4226 528278 4294
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 527658 4102 528278 4170
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 527658 -160 528278 3922
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 531378 46350 531998 48690
rect 531378 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 531998 46350
rect 531378 46226 531998 46294
rect 531378 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 531998 46226
rect 531378 46102 531998 46170
rect 531378 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 531998 46102
rect 531378 45978 531998 46046
rect 531378 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 531998 45978
rect 531378 28350 531998 45922
rect 531378 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 531998 28350
rect 531378 28226 531998 28294
rect 531378 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 531998 28226
rect 531378 28102 531998 28170
rect 531378 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 531998 28102
rect 531378 27978 531998 28046
rect 531378 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 531998 27978
rect 531378 10350 531998 27922
rect 531378 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 531998 10350
rect 531378 10226 531998 10294
rect 531378 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 531998 10226
rect 531378 10102 531998 10170
rect 531378 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 531998 10102
rect 531378 9978 531998 10046
rect 531378 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 531998 9978
rect 531378 -1120 531998 9922
rect 531378 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 531998 -1120
rect 531378 -1244 531998 -1176
rect 531378 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 531998 -1244
rect 531378 -1368 531998 -1300
rect 531378 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 531998 -1368
rect 531378 -1492 531998 -1424
rect 531378 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 531998 -1492
rect 531378 -1644 531998 -1548
rect 558378 40350 558998 48690
rect 559804 45108 559860 84924
rect 559804 45042 559860 45052
rect 562098 82350 562718 99922
rect 562828 167300 562884 167310
rect 562828 92820 562884 167244
rect 563052 165620 563108 165630
rect 562940 163828 562996 163838
rect 562940 97524 562996 163772
rect 563052 100660 563108 165564
rect 563164 106932 563220 168812
rect 563388 164052 563444 164062
rect 563164 106866 563220 106876
rect 563276 162260 563332 162270
rect 563276 102228 563332 162204
rect 563388 103796 563444 163996
rect 566188 160678 566244 160688
rect 564620 160498 564676 160508
rect 564508 158698 564564 158708
rect 563612 152740 563668 152750
rect 563388 103730 563444 103740
rect 563500 150500 563556 150510
rect 563276 102162 563332 102172
rect 563052 100594 563108 100604
rect 562940 97458 562996 97468
rect 562828 92754 562884 92764
rect 563500 91252 563556 150444
rect 563612 94388 563668 152684
rect 563724 152628 563780 152638
rect 563724 99092 563780 152572
rect 564508 110068 564564 158642
rect 564620 113204 564676 160442
rect 564732 155458 564788 155468
rect 564732 116340 564788 155402
rect 566188 121044 566244 160622
rect 566188 120978 566244 120988
rect 564732 116274 564788 116284
rect 564620 113138 564676 113148
rect 564508 110002 564564 110012
rect 563724 99026 563780 99036
rect 563612 94322 563668 94332
rect 563500 91186 563556 91196
rect 562098 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 562718 82350
rect 562098 82226 562718 82294
rect 562098 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 562718 82226
rect 562098 82102 562718 82170
rect 562098 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 562718 82102
rect 562098 81978 562718 82046
rect 562098 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 562718 81978
rect 562098 64350 562718 81922
rect 562098 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 562718 64350
rect 562098 64226 562718 64294
rect 562098 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 562718 64226
rect 562098 64102 562718 64170
rect 562098 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 562718 64102
rect 562098 63978 562718 64046
rect 562098 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 562718 63978
rect 562098 46350 562718 63922
rect 562098 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 562718 46350
rect 562098 46226 562718 46294
rect 562098 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 562718 46226
rect 562098 46102 562718 46170
rect 562098 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 562718 46102
rect 562098 45978 562718 46046
rect 562098 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 562718 45978
rect 558378 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 558998 40350
rect 558378 40226 558998 40294
rect 558378 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 558998 40226
rect 558378 40102 558998 40170
rect 558378 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 558998 40102
rect 558378 39978 558998 40046
rect 558378 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 558998 39978
rect 558378 22350 558998 39922
rect 558378 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 558998 22350
rect 558378 22226 558998 22294
rect 558378 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 558998 22226
rect 558378 22102 558998 22170
rect 558378 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 558998 22102
rect 558378 21978 558998 22046
rect 558378 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 558998 21978
rect 558378 4350 558998 21922
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 558378 -160 558998 3922
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 562098 28350 562718 45922
rect 562828 83412 562884 83422
rect 562828 45220 562884 83356
rect 562940 74004 562996 74014
rect 562940 50036 562996 73948
rect 563052 66164 563108 66174
rect 563052 50148 563108 66108
rect 563052 50082 563108 50092
rect 563164 64596 563220 64606
rect 562940 49970 562996 49980
rect 563164 48132 563220 64540
rect 563164 48066 563220 48076
rect 562828 45154 562884 45164
rect 562098 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 562718 28350
rect 562098 28226 562718 28294
rect 562098 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 562718 28226
rect 562098 28102 562718 28170
rect 562098 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 562718 28102
rect 562098 27978 562718 28046
rect 562098 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 562718 27978
rect 562098 10350 562718 27922
rect 572012 20356 572068 402002
rect 573692 401878 573748 401888
rect 573692 60004 573748 401822
rect 575372 401698 575428 401708
rect 575372 139300 575428 401642
rect 589098 400350 589718 417922
rect 590492 509348 590548 509358
rect 590492 404038 590548 509292
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 590492 403972 590548 403982
rect 590604 469700 590660 469710
rect 590604 402418 590660 469644
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 590604 402352 590660 402362
rect 590716 430164 590772 430174
rect 590716 402388 590772 430108
rect 590716 402322 590772 402332
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 581308 395218 581364 395228
rect 579628 393778 579684 393788
rect 577052 393418 577108 393428
rect 577052 218596 577108 393362
rect 577052 218530 577108 218540
rect 575372 139234 575428 139244
rect 573692 59938 573748 59948
rect 572012 20290 572068 20300
rect 562098 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 562718 10350
rect 562098 10226 562718 10294
rect 562098 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 562718 10226
rect 562098 10102 562718 10170
rect 562098 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 562718 10102
rect 562098 9978 562718 10046
rect 562098 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 562718 9978
rect 562098 -1120 562718 9922
rect 579628 4228 579684 393722
rect 579628 4162 579684 4172
rect 581308 4228 581364 395162
rect 581308 4162 581364 4172
rect 582988 395038 583044 395048
rect 582988 4228 583044 394982
rect 585452 393238 585508 393248
rect 585452 99876 585508 393182
rect 585452 99810 585508 99820
rect 589098 382350 589718 399922
rect 590940 401604 590996 401614
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 589098 364350 589718 381922
rect 590492 392158 590548 392168
rect 590492 377412 590548 392102
rect 590940 390628 590996 401548
rect 590940 390562 590996 390572
rect 590492 377346 590548 377356
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 589098 363978 589718 364046
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 589098 346350 589718 363922
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 589098 328350 589718 345922
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 589098 310350 589718 327922
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 589098 292350 589718 309922
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 589098 274350 589718 291922
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 589098 256350 589718 273922
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 589098 238350 589718 255922
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 589098 220350 589718 237922
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 589098 202350 589718 219922
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 589098 184350 589718 201922
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 589098 166350 589718 183922
rect 590492 311108 590548 311118
rect 590492 175364 590548 311052
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 590492 175298 590548 175308
rect 590604 271460 590660 271470
rect 590604 173572 590660 271404
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 590716 231924 590772 231934
rect 590716 175476 590772 231868
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 590716 175410 590772 175420
rect 590828 192164 590884 192174
rect 590604 173506 590660 173516
rect 590828 167972 590884 192108
rect 590828 167906 590884 167916
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 589098 148350 589718 165922
rect 590604 165508 590660 165518
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 589098 130350 589718 147922
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 589098 112350 589718 129922
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 582988 4162 583044 4172
rect 589098 94350 589718 111922
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 589098 76350 589718 93922
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 589098 58350 589718 75922
rect 590492 150418 590548 150428
rect 590492 73444 590548 150362
rect 590604 113092 590660 165452
rect 590604 113026 590660 113036
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 590492 73378 590548 73388
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 589098 40350 589718 57922
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 589098 22350 589718 39922
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 589098 4350 589718 21922
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 562098 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 562718 -1120
rect 562098 -1244 562718 -1176
rect 562098 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 562718 -1244
rect 562098 -1368 562718 -1300
rect 562098 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 562718 -1368
rect 562098 -1492 562718 -1424
rect 562098 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 562718 -1492
rect 562098 -1644 562718 -1548
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect 4172 376262 4228 376318
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 4172 247022 4228 247078
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect 4172 206522 4228 206578
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect 4172 164582 4228 164638
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 9234 568294 9290 568350
rect 9358 568294 9414 568350
rect 9482 568294 9538 568350
rect 9606 568294 9662 568350
rect 9234 568170 9290 568226
rect 9358 568170 9414 568226
rect 9482 568170 9538 568226
rect 9606 568170 9662 568226
rect 9234 568046 9290 568102
rect 9358 568046 9414 568102
rect 9482 568046 9538 568102
rect 9606 568046 9662 568102
rect 9234 567922 9290 567978
rect 9358 567922 9414 567978
rect 9482 567922 9538 567978
rect 9606 567922 9662 567978
rect 9234 550294 9290 550350
rect 9358 550294 9414 550350
rect 9482 550294 9538 550350
rect 9606 550294 9662 550350
rect 9234 550170 9290 550226
rect 9358 550170 9414 550226
rect 9482 550170 9538 550226
rect 9606 550170 9662 550226
rect 9234 550046 9290 550102
rect 9358 550046 9414 550102
rect 9482 550046 9538 550102
rect 9606 550046 9662 550102
rect 9234 549922 9290 549978
rect 9358 549922 9414 549978
rect 9482 549922 9538 549978
rect 9606 549922 9662 549978
rect 9234 532294 9290 532350
rect 9358 532294 9414 532350
rect 9482 532294 9538 532350
rect 9606 532294 9662 532350
rect 9234 532170 9290 532226
rect 9358 532170 9414 532226
rect 9482 532170 9538 532226
rect 9606 532170 9662 532226
rect 9234 532046 9290 532102
rect 9358 532046 9414 532102
rect 9482 532046 9538 532102
rect 9606 532046 9662 532102
rect 9234 531922 9290 531978
rect 9358 531922 9414 531978
rect 9482 531922 9538 531978
rect 9606 531922 9662 531978
rect 9234 514294 9290 514350
rect 9358 514294 9414 514350
rect 9482 514294 9538 514350
rect 9606 514294 9662 514350
rect 9234 514170 9290 514226
rect 9358 514170 9414 514226
rect 9482 514170 9538 514226
rect 9606 514170 9662 514226
rect 9234 514046 9290 514102
rect 9358 514046 9414 514102
rect 9482 514046 9538 514102
rect 9606 514046 9662 514102
rect 9234 513922 9290 513978
rect 9358 513922 9414 513978
rect 9482 513922 9538 513978
rect 9606 513922 9662 513978
rect 9234 496294 9290 496350
rect 9358 496294 9414 496350
rect 9482 496294 9538 496350
rect 9606 496294 9662 496350
rect 9234 496170 9290 496226
rect 9358 496170 9414 496226
rect 9482 496170 9538 496226
rect 9606 496170 9662 496226
rect 9234 496046 9290 496102
rect 9358 496046 9414 496102
rect 9482 496046 9538 496102
rect 9606 496046 9662 496102
rect 9234 495922 9290 495978
rect 9358 495922 9414 495978
rect 9482 495922 9538 495978
rect 9606 495922 9662 495978
rect 9234 478294 9290 478350
rect 9358 478294 9414 478350
rect 9482 478294 9538 478350
rect 9606 478294 9662 478350
rect 9234 478170 9290 478226
rect 9358 478170 9414 478226
rect 9482 478170 9538 478226
rect 9606 478170 9662 478226
rect 9234 478046 9290 478102
rect 9358 478046 9414 478102
rect 9482 478046 9538 478102
rect 9606 478046 9662 478102
rect 9234 477922 9290 477978
rect 9358 477922 9414 477978
rect 9482 477922 9538 477978
rect 9606 477922 9662 477978
rect 9234 460294 9290 460350
rect 9358 460294 9414 460350
rect 9482 460294 9538 460350
rect 9606 460294 9662 460350
rect 9234 460170 9290 460226
rect 9358 460170 9414 460226
rect 9482 460170 9538 460226
rect 9606 460170 9662 460226
rect 9234 460046 9290 460102
rect 9358 460046 9414 460102
rect 9482 460046 9538 460102
rect 9606 460046 9662 460102
rect 9234 459922 9290 459978
rect 9358 459922 9414 459978
rect 9482 459922 9538 459978
rect 9606 459922 9662 459978
rect 9234 442294 9290 442350
rect 9358 442294 9414 442350
rect 9482 442294 9538 442350
rect 9606 442294 9662 442350
rect 9234 442170 9290 442226
rect 9358 442170 9414 442226
rect 9482 442170 9538 442226
rect 9606 442170 9662 442226
rect 9234 442046 9290 442102
rect 9358 442046 9414 442102
rect 9482 442046 9538 442102
rect 9606 442046 9662 442102
rect 9234 441922 9290 441978
rect 9358 441922 9414 441978
rect 9482 441922 9538 441978
rect 9606 441922 9662 441978
rect 9234 424294 9290 424350
rect 9358 424294 9414 424350
rect 9482 424294 9538 424350
rect 9606 424294 9662 424350
rect 9234 424170 9290 424226
rect 9358 424170 9414 424226
rect 9482 424170 9538 424226
rect 9606 424170 9662 424226
rect 9234 424046 9290 424102
rect 9358 424046 9414 424102
rect 9482 424046 9538 424102
rect 9606 424046 9662 424102
rect 9234 423922 9290 423978
rect 9358 423922 9414 423978
rect 9482 423922 9538 423978
rect 9606 423922 9662 423978
rect 9234 406294 9290 406350
rect 9358 406294 9414 406350
rect 9482 406294 9538 406350
rect 9606 406294 9662 406350
rect 9234 406170 9290 406226
rect 9358 406170 9414 406226
rect 9482 406170 9538 406226
rect 9606 406170 9662 406226
rect 9234 406046 9290 406102
rect 9358 406046 9414 406102
rect 9482 406046 9538 406102
rect 9606 406046 9662 406102
rect 9234 405922 9290 405978
rect 9358 405922 9414 405978
rect 9482 405922 9538 405978
rect 9606 405922 9662 405978
rect 9234 388294 9290 388350
rect 9358 388294 9414 388350
rect 9482 388294 9538 388350
rect 9606 388294 9662 388350
rect 9234 388170 9290 388226
rect 9358 388170 9414 388226
rect 9482 388170 9538 388226
rect 9606 388170 9662 388226
rect 9234 388046 9290 388102
rect 9358 388046 9414 388102
rect 9482 388046 9538 388102
rect 9606 388046 9662 388102
rect 9234 387922 9290 387978
rect 9358 387922 9414 387978
rect 9482 387922 9538 387978
rect 9606 387922 9662 387978
rect 9234 370294 9290 370350
rect 9358 370294 9414 370350
rect 9482 370294 9538 370350
rect 9606 370294 9662 370350
rect 9234 370170 9290 370226
rect 9358 370170 9414 370226
rect 9482 370170 9538 370226
rect 9606 370170 9662 370226
rect 9234 370046 9290 370102
rect 9358 370046 9414 370102
rect 9482 370046 9538 370102
rect 9606 370046 9662 370102
rect 9234 369922 9290 369978
rect 9358 369922 9414 369978
rect 9482 369922 9538 369978
rect 9606 369922 9662 369978
rect 9234 352294 9290 352350
rect 9358 352294 9414 352350
rect 9482 352294 9538 352350
rect 9606 352294 9662 352350
rect 9234 352170 9290 352226
rect 9358 352170 9414 352226
rect 9482 352170 9538 352226
rect 9606 352170 9662 352226
rect 9234 352046 9290 352102
rect 9358 352046 9414 352102
rect 9482 352046 9538 352102
rect 9606 352046 9662 352102
rect 9234 351922 9290 351978
rect 9358 351922 9414 351978
rect 9482 351922 9538 351978
rect 9606 351922 9662 351978
rect 9234 334294 9290 334350
rect 9358 334294 9414 334350
rect 9482 334294 9538 334350
rect 9606 334294 9662 334350
rect 9234 334170 9290 334226
rect 9358 334170 9414 334226
rect 9482 334170 9538 334226
rect 9606 334170 9662 334226
rect 9234 334046 9290 334102
rect 9358 334046 9414 334102
rect 9482 334046 9538 334102
rect 9606 334046 9662 334102
rect 9234 333922 9290 333978
rect 9358 333922 9414 333978
rect 9482 333922 9538 333978
rect 9606 333922 9662 333978
rect 9234 316294 9290 316350
rect 9358 316294 9414 316350
rect 9482 316294 9538 316350
rect 9606 316294 9662 316350
rect 9234 316170 9290 316226
rect 9358 316170 9414 316226
rect 9482 316170 9538 316226
rect 9606 316170 9662 316226
rect 9234 316046 9290 316102
rect 9358 316046 9414 316102
rect 9482 316046 9538 316102
rect 9606 316046 9662 316102
rect 9234 315922 9290 315978
rect 9358 315922 9414 315978
rect 9482 315922 9538 315978
rect 9606 315922 9662 315978
rect 9234 298294 9290 298350
rect 9358 298294 9414 298350
rect 9482 298294 9538 298350
rect 9606 298294 9662 298350
rect 9234 298170 9290 298226
rect 9358 298170 9414 298226
rect 9482 298170 9538 298226
rect 9606 298170 9662 298226
rect 9234 298046 9290 298102
rect 9358 298046 9414 298102
rect 9482 298046 9538 298102
rect 9606 298046 9662 298102
rect 9234 297922 9290 297978
rect 9358 297922 9414 297978
rect 9482 297922 9538 297978
rect 9606 297922 9662 297978
rect 9234 280294 9290 280350
rect 9358 280294 9414 280350
rect 9482 280294 9538 280350
rect 9606 280294 9662 280350
rect 9234 280170 9290 280226
rect 9358 280170 9414 280226
rect 9482 280170 9538 280226
rect 9606 280170 9662 280226
rect 9234 280046 9290 280102
rect 9358 280046 9414 280102
rect 9482 280046 9538 280102
rect 9606 280046 9662 280102
rect 9234 279922 9290 279978
rect 9358 279922 9414 279978
rect 9482 279922 9538 279978
rect 9606 279922 9662 279978
rect 9234 262294 9290 262350
rect 9358 262294 9414 262350
rect 9482 262294 9538 262350
rect 9606 262294 9662 262350
rect 9234 262170 9290 262226
rect 9358 262170 9414 262226
rect 9482 262170 9538 262226
rect 9606 262170 9662 262226
rect 9234 262046 9290 262102
rect 9358 262046 9414 262102
rect 9482 262046 9538 262102
rect 9606 262046 9662 262102
rect 9234 261922 9290 261978
rect 9358 261922 9414 261978
rect 9482 261922 9538 261978
rect 9606 261922 9662 261978
rect 9234 244294 9290 244350
rect 9358 244294 9414 244350
rect 9482 244294 9538 244350
rect 9606 244294 9662 244350
rect 9234 244170 9290 244226
rect 9358 244170 9414 244226
rect 9482 244170 9538 244226
rect 9606 244170 9662 244226
rect 9234 244046 9290 244102
rect 9358 244046 9414 244102
rect 9482 244046 9538 244102
rect 9606 244046 9662 244102
rect 9234 243922 9290 243978
rect 9358 243922 9414 243978
rect 9482 243922 9538 243978
rect 9606 243922 9662 243978
rect 36234 597156 36290 597212
rect 36358 597156 36414 597212
rect 36482 597156 36538 597212
rect 36606 597156 36662 597212
rect 36234 597032 36290 597088
rect 36358 597032 36414 597088
rect 36482 597032 36538 597088
rect 36606 597032 36662 597088
rect 36234 596908 36290 596964
rect 36358 596908 36414 596964
rect 36482 596908 36538 596964
rect 36606 596908 36662 596964
rect 36234 596784 36290 596840
rect 36358 596784 36414 596840
rect 36482 596784 36538 596840
rect 36606 596784 36662 596840
rect 36234 580294 36290 580350
rect 36358 580294 36414 580350
rect 36482 580294 36538 580350
rect 36606 580294 36662 580350
rect 36234 580170 36290 580226
rect 36358 580170 36414 580226
rect 36482 580170 36538 580226
rect 36606 580170 36662 580226
rect 36234 580046 36290 580102
rect 36358 580046 36414 580102
rect 36482 580046 36538 580102
rect 36606 580046 36662 580102
rect 36234 579922 36290 579978
rect 36358 579922 36414 579978
rect 36482 579922 36538 579978
rect 36606 579922 36662 579978
rect 36234 562294 36290 562350
rect 36358 562294 36414 562350
rect 36482 562294 36538 562350
rect 36606 562294 36662 562350
rect 36234 562170 36290 562226
rect 36358 562170 36414 562226
rect 36482 562170 36538 562226
rect 36606 562170 36662 562226
rect 36234 562046 36290 562102
rect 36358 562046 36414 562102
rect 36482 562046 36538 562102
rect 36606 562046 36662 562102
rect 36234 561922 36290 561978
rect 36358 561922 36414 561978
rect 36482 561922 36538 561978
rect 36606 561922 36662 561978
rect 36234 544294 36290 544350
rect 36358 544294 36414 544350
rect 36482 544294 36538 544350
rect 36606 544294 36662 544350
rect 36234 544170 36290 544226
rect 36358 544170 36414 544226
rect 36482 544170 36538 544226
rect 36606 544170 36662 544226
rect 36234 544046 36290 544102
rect 36358 544046 36414 544102
rect 36482 544046 36538 544102
rect 36606 544046 36662 544102
rect 36234 543922 36290 543978
rect 36358 543922 36414 543978
rect 36482 543922 36538 543978
rect 36606 543922 36662 543978
rect 36234 526294 36290 526350
rect 36358 526294 36414 526350
rect 36482 526294 36538 526350
rect 36606 526294 36662 526350
rect 36234 526170 36290 526226
rect 36358 526170 36414 526226
rect 36482 526170 36538 526226
rect 36606 526170 36662 526226
rect 36234 526046 36290 526102
rect 36358 526046 36414 526102
rect 36482 526046 36538 526102
rect 36606 526046 36662 526102
rect 36234 525922 36290 525978
rect 36358 525922 36414 525978
rect 36482 525922 36538 525978
rect 36606 525922 36662 525978
rect 36234 508294 36290 508350
rect 36358 508294 36414 508350
rect 36482 508294 36538 508350
rect 36606 508294 36662 508350
rect 36234 508170 36290 508226
rect 36358 508170 36414 508226
rect 36482 508170 36538 508226
rect 36606 508170 36662 508226
rect 36234 508046 36290 508102
rect 36358 508046 36414 508102
rect 36482 508046 36538 508102
rect 36606 508046 36662 508102
rect 36234 507922 36290 507978
rect 36358 507922 36414 507978
rect 36482 507922 36538 507978
rect 36606 507922 36662 507978
rect 36234 490294 36290 490350
rect 36358 490294 36414 490350
rect 36482 490294 36538 490350
rect 36606 490294 36662 490350
rect 36234 490170 36290 490226
rect 36358 490170 36414 490226
rect 36482 490170 36538 490226
rect 36606 490170 36662 490226
rect 36234 490046 36290 490102
rect 36358 490046 36414 490102
rect 36482 490046 36538 490102
rect 36606 490046 36662 490102
rect 36234 489922 36290 489978
rect 36358 489922 36414 489978
rect 36482 489922 36538 489978
rect 36606 489922 36662 489978
rect 36234 472294 36290 472350
rect 36358 472294 36414 472350
rect 36482 472294 36538 472350
rect 36606 472294 36662 472350
rect 36234 472170 36290 472226
rect 36358 472170 36414 472226
rect 36482 472170 36538 472226
rect 36606 472170 36662 472226
rect 36234 472046 36290 472102
rect 36358 472046 36414 472102
rect 36482 472046 36538 472102
rect 36606 472046 36662 472102
rect 36234 471922 36290 471978
rect 36358 471922 36414 471978
rect 36482 471922 36538 471978
rect 36606 471922 36662 471978
rect 36234 454294 36290 454350
rect 36358 454294 36414 454350
rect 36482 454294 36538 454350
rect 36606 454294 36662 454350
rect 36234 454170 36290 454226
rect 36358 454170 36414 454226
rect 36482 454170 36538 454226
rect 36606 454170 36662 454226
rect 36234 454046 36290 454102
rect 36358 454046 36414 454102
rect 36482 454046 36538 454102
rect 36606 454046 36662 454102
rect 36234 453922 36290 453978
rect 36358 453922 36414 453978
rect 36482 453922 36538 453978
rect 36606 453922 36662 453978
rect 36234 436294 36290 436350
rect 36358 436294 36414 436350
rect 36482 436294 36538 436350
rect 36606 436294 36662 436350
rect 36234 436170 36290 436226
rect 36358 436170 36414 436226
rect 36482 436170 36538 436226
rect 36606 436170 36662 436226
rect 36234 436046 36290 436102
rect 36358 436046 36414 436102
rect 36482 436046 36538 436102
rect 36606 436046 36662 436102
rect 36234 435922 36290 435978
rect 36358 435922 36414 435978
rect 36482 435922 36538 435978
rect 36606 435922 36662 435978
rect 36234 418294 36290 418350
rect 36358 418294 36414 418350
rect 36482 418294 36538 418350
rect 36606 418294 36662 418350
rect 36234 418170 36290 418226
rect 36358 418170 36414 418226
rect 36482 418170 36538 418226
rect 36606 418170 36662 418226
rect 36234 418046 36290 418102
rect 36358 418046 36414 418102
rect 36482 418046 36538 418102
rect 36606 418046 36662 418102
rect 36234 417922 36290 417978
rect 36358 417922 36414 417978
rect 36482 417922 36538 417978
rect 36606 417922 36662 417978
rect 36234 400294 36290 400350
rect 36358 400294 36414 400350
rect 36482 400294 36538 400350
rect 36606 400294 36662 400350
rect 36234 400170 36290 400226
rect 36358 400170 36414 400226
rect 36482 400170 36538 400226
rect 36606 400170 36662 400226
rect 36234 400046 36290 400102
rect 36358 400046 36414 400102
rect 36482 400046 36538 400102
rect 36606 400046 36662 400102
rect 36234 399922 36290 399978
rect 36358 399922 36414 399978
rect 36482 399922 36538 399978
rect 36606 399922 36662 399978
rect 36234 382294 36290 382350
rect 36358 382294 36414 382350
rect 36482 382294 36538 382350
rect 36606 382294 36662 382350
rect 36234 382170 36290 382226
rect 36358 382170 36414 382226
rect 36482 382170 36538 382226
rect 36606 382170 36662 382226
rect 36234 382046 36290 382102
rect 36358 382046 36414 382102
rect 36482 382046 36538 382102
rect 36606 382046 36662 382102
rect 36234 381922 36290 381978
rect 36358 381922 36414 381978
rect 36482 381922 36538 381978
rect 36606 381922 36662 381978
rect 36234 364294 36290 364350
rect 36358 364294 36414 364350
rect 36482 364294 36538 364350
rect 36606 364294 36662 364350
rect 36234 364170 36290 364226
rect 36358 364170 36414 364226
rect 36482 364170 36538 364226
rect 36606 364170 36662 364226
rect 36234 364046 36290 364102
rect 36358 364046 36414 364102
rect 36482 364046 36538 364102
rect 36606 364046 36662 364102
rect 36234 363922 36290 363978
rect 36358 363922 36414 363978
rect 36482 363922 36538 363978
rect 36606 363922 36662 363978
rect 36234 346294 36290 346350
rect 36358 346294 36414 346350
rect 36482 346294 36538 346350
rect 36606 346294 36662 346350
rect 36234 346170 36290 346226
rect 36358 346170 36414 346226
rect 36482 346170 36538 346226
rect 36606 346170 36662 346226
rect 36234 346046 36290 346102
rect 36358 346046 36414 346102
rect 36482 346046 36538 346102
rect 36606 346046 36662 346102
rect 36234 345922 36290 345978
rect 36358 345922 36414 345978
rect 36482 345922 36538 345978
rect 36606 345922 36662 345978
rect 36234 328294 36290 328350
rect 36358 328294 36414 328350
rect 36482 328294 36538 328350
rect 36606 328294 36662 328350
rect 36234 328170 36290 328226
rect 36358 328170 36414 328226
rect 36482 328170 36538 328226
rect 36606 328170 36662 328226
rect 36234 328046 36290 328102
rect 36358 328046 36414 328102
rect 36482 328046 36538 328102
rect 36606 328046 36662 328102
rect 36234 327922 36290 327978
rect 36358 327922 36414 327978
rect 36482 327922 36538 327978
rect 36606 327922 36662 327978
rect 36234 310294 36290 310350
rect 36358 310294 36414 310350
rect 36482 310294 36538 310350
rect 36606 310294 36662 310350
rect 36234 310170 36290 310226
rect 36358 310170 36414 310226
rect 36482 310170 36538 310226
rect 36606 310170 36662 310226
rect 36234 310046 36290 310102
rect 36358 310046 36414 310102
rect 36482 310046 36538 310102
rect 36606 310046 36662 310102
rect 36234 309922 36290 309978
rect 36358 309922 36414 309978
rect 36482 309922 36538 309978
rect 36606 309922 36662 309978
rect 36234 292294 36290 292350
rect 36358 292294 36414 292350
rect 36482 292294 36538 292350
rect 36606 292294 36662 292350
rect 36234 292170 36290 292226
rect 36358 292170 36414 292226
rect 36482 292170 36538 292226
rect 36606 292170 36662 292226
rect 36234 292046 36290 292102
rect 36358 292046 36414 292102
rect 36482 292046 36538 292102
rect 36606 292046 36662 292102
rect 36234 291922 36290 291978
rect 36358 291922 36414 291978
rect 36482 291922 36538 291978
rect 36606 291922 36662 291978
rect 36234 274294 36290 274350
rect 36358 274294 36414 274350
rect 36482 274294 36538 274350
rect 36606 274294 36662 274350
rect 36234 274170 36290 274226
rect 36358 274170 36414 274226
rect 36482 274170 36538 274226
rect 36606 274170 36662 274226
rect 36234 274046 36290 274102
rect 36358 274046 36414 274102
rect 36482 274046 36538 274102
rect 36606 274046 36662 274102
rect 36234 273922 36290 273978
rect 36358 273922 36414 273978
rect 36482 273922 36538 273978
rect 36606 273922 36662 273978
rect 36234 256294 36290 256350
rect 36358 256294 36414 256350
rect 36482 256294 36538 256350
rect 36606 256294 36662 256350
rect 36234 256170 36290 256226
rect 36358 256170 36414 256226
rect 36482 256170 36538 256226
rect 36606 256170 36662 256226
rect 36234 256046 36290 256102
rect 36358 256046 36414 256102
rect 36482 256046 36538 256102
rect 36606 256046 36662 256102
rect 36234 255922 36290 255978
rect 36358 255922 36414 255978
rect 36482 255922 36538 255978
rect 36606 255922 36662 255978
rect 35196 241082 35252 241138
rect 9234 226294 9290 226350
rect 9358 226294 9414 226350
rect 9482 226294 9538 226350
rect 9606 226294 9662 226350
rect 9234 226170 9290 226226
rect 9358 226170 9414 226226
rect 9482 226170 9538 226226
rect 9606 226170 9662 226226
rect 9234 226046 9290 226102
rect 9358 226046 9414 226102
rect 9482 226046 9538 226102
rect 9606 226046 9662 226102
rect 9234 225922 9290 225978
rect 9358 225922 9414 225978
rect 9482 225922 9538 225978
rect 9606 225922 9662 225978
rect 9234 208294 9290 208350
rect 9358 208294 9414 208350
rect 9482 208294 9538 208350
rect 9606 208294 9662 208350
rect 9234 208170 9290 208226
rect 9358 208170 9414 208226
rect 9482 208170 9538 208226
rect 9606 208170 9662 208226
rect 9234 208046 9290 208102
rect 9358 208046 9414 208102
rect 9482 208046 9538 208102
rect 9606 208046 9662 208102
rect 9234 207922 9290 207978
rect 9358 207922 9414 207978
rect 9482 207922 9538 207978
rect 9606 207922 9662 207978
rect 9234 190294 9290 190350
rect 9358 190294 9414 190350
rect 9482 190294 9538 190350
rect 9606 190294 9662 190350
rect 9234 190170 9290 190226
rect 9358 190170 9414 190226
rect 9482 190170 9538 190226
rect 9606 190170 9662 190226
rect 9234 190046 9290 190102
rect 9358 190046 9414 190102
rect 9482 190046 9538 190102
rect 9606 190046 9662 190102
rect 9234 189922 9290 189978
rect 9358 189922 9414 189978
rect 9482 189922 9538 189978
rect 9606 189922 9662 189978
rect 9234 172294 9290 172350
rect 9358 172294 9414 172350
rect 9482 172294 9538 172350
rect 9606 172294 9662 172350
rect 9234 172170 9290 172226
rect 9358 172170 9414 172226
rect 9482 172170 9538 172226
rect 9606 172170 9662 172226
rect 9234 172046 9290 172102
rect 9358 172046 9414 172102
rect 9482 172046 9538 172102
rect 9606 172046 9662 172102
rect 9234 171922 9290 171978
rect 9358 171922 9414 171978
rect 9482 171922 9538 171978
rect 9606 171922 9662 171978
rect 9234 154294 9290 154350
rect 9358 154294 9414 154350
rect 9482 154294 9538 154350
rect 9606 154294 9662 154350
rect 9234 154170 9290 154226
rect 9358 154170 9414 154226
rect 9482 154170 9538 154226
rect 9606 154170 9662 154226
rect 9234 154046 9290 154102
rect 9358 154046 9414 154102
rect 9482 154046 9538 154102
rect 9606 154046 9662 154102
rect 9234 153922 9290 153978
rect 9358 153922 9414 153978
rect 9482 153922 9538 153978
rect 9606 153922 9662 153978
rect 9234 136294 9290 136350
rect 9358 136294 9414 136350
rect 9482 136294 9538 136350
rect 9606 136294 9662 136350
rect 9234 136170 9290 136226
rect 9358 136170 9414 136226
rect 9482 136170 9538 136226
rect 9606 136170 9662 136226
rect 9234 136046 9290 136102
rect 9358 136046 9414 136102
rect 9482 136046 9538 136102
rect 9606 136046 9662 136102
rect 9234 135922 9290 135978
rect 9358 135922 9414 135978
rect 9482 135922 9538 135978
rect 9606 135922 9662 135978
rect 9234 118294 9290 118350
rect 9358 118294 9414 118350
rect 9482 118294 9538 118350
rect 9606 118294 9662 118350
rect 9234 118170 9290 118226
rect 9358 118170 9414 118226
rect 9482 118170 9538 118226
rect 9606 118170 9662 118226
rect 9234 118046 9290 118102
rect 9358 118046 9414 118102
rect 9482 118046 9538 118102
rect 9606 118046 9662 118102
rect 9234 117922 9290 117978
rect 9358 117922 9414 117978
rect 9482 117922 9538 117978
rect 9606 117922 9662 117978
rect 9234 100294 9290 100350
rect 9358 100294 9414 100350
rect 9482 100294 9538 100350
rect 9606 100294 9662 100350
rect 9234 100170 9290 100226
rect 9358 100170 9414 100226
rect 9482 100170 9538 100226
rect 9606 100170 9662 100226
rect 9234 100046 9290 100102
rect 9358 100046 9414 100102
rect 9482 100046 9538 100102
rect 9606 100046 9662 100102
rect 9234 99922 9290 99978
rect 9358 99922 9414 99978
rect 9482 99922 9538 99978
rect 9606 99922 9662 99978
rect 9234 82294 9290 82350
rect 9358 82294 9414 82350
rect 9482 82294 9538 82350
rect 9606 82294 9662 82350
rect 9234 82170 9290 82226
rect 9358 82170 9414 82226
rect 9482 82170 9538 82226
rect 9606 82170 9662 82226
rect 9234 82046 9290 82102
rect 9358 82046 9414 82102
rect 9482 82046 9538 82102
rect 9606 82046 9662 82102
rect 9234 81922 9290 81978
rect 9358 81922 9414 81978
rect 9482 81922 9538 81978
rect 9606 81922 9662 81978
rect 9234 64294 9290 64350
rect 9358 64294 9414 64350
rect 9482 64294 9538 64350
rect 9606 64294 9662 64350
rect 9234 64170 9290 64226
rect 9358 64170 9414 64226
rect 9482 64170 9538 64226
rect 9606 64170 9662 64226
rect 9234 64046 9290 64102
rect 9358 64046 9414 64102
rect 9482 64046 9538 64102
rect 9606 64046 9662 64102
rect 9234 63922 9290 63978
rect 9358 63922 9414 63978
rect 9482 63922 9538 63978
rect 9606 63922 9662 63978
rect 9234 46294 9290 46350
rect 9358 46294 9414 46350
rect 9482 46294 9538 46350
rect 9606 46294 9662 46350
rect 9234 46170 9290 46226
rect 9358 46170 9414 46226
rect 9482 46170 9538 46226
rect 9606 46170 9662 46226
rect 9234 46046 9290 46102
rect 9358 46046 9414 46102
rect 9482 46046 9538 46102
rect 9606 46046 9662 46102
rect 9234 45922 9290 45978
rect 9358 45922 9414 45978
rect 9482 45922 9538 45978
rect 9606 45922 9662 45978
rect 9234 28294 9290 28350
rect 9358 28294 9414 28350
rect 9482 28294 9538 28350
rect 9606 28294 9662 28350
rect 9234 28170 9290 28226
rect 9358 28170 9414 28226
rect 9482 28170 9538 28226
rect 9606 28170 9662 28226
rect 9234 28046 9290 28102
rect 9358 28046 9414 28102
rect 9482 28046 9538 28102
rect 9606 28046 9662 28102
rect 9234 27922 9290 27978
rect 9358 27922 9414 27978
rect 9482 27922 9538 27978
rect 9606 27922 9662 27978
rect 9234 10294 9290 10350
rect 9358 10294 9414 10350
rect 9482 10294 9538 10350
rect 9606 10294 9662 10350
rect 9234 10170 9290 10226
rect 9358 10170 9414 10226
rect 9482 10170 9538 10226
rect 9606 10170 9662 10226
rect 9234 10046 9290 10102
rect 9358 10046 9414 10102
rect 9482 10046 9538 10102
rect 9606 10046 9662 10102
rect 9234 9922 9290 9978
rect 9358 9922 9414 9978
rect 9482 9922 9538 9978
rect 9606 9922 9662 9978
rect 16716 234242 16772 234298
rect 25116 231002 25172 231058
rect 18396 227582 18452 227638
rect 20076 224162 20132 224218
rect 35084 230282 35140 230338
rect 34972 4742 35028 4798
rect 36234 238294 36290 238350
rect 36358 238294 36414 238350
rect 36482 238294 36538 238350
rect 36606 238294 36662 238350
rect 36234 238170 36290 238226
rect 36358 238170 36414 238226
rect 36482 238170 36538 238226
rect 36606 238170 36662 238226
rect 36234 238046 36290 238102
rect 36358 238046 36414 238102
rect 36482 238046 36538 238102
rect 36606 238046 36662 238102
rect 36234 237922 36290 237978
rect 36358 237922 36414 237978
rect 36482 237922 36538 237978
rect 36606 237922 36662 237978
rect 36234 220294 36290 220350
rect 36358 220294 36414 220350
rect 36482 220294 36538 220350
rect 36606 220294 36662 220350
rect 36234 220170 36290 220226
rect 36358 220170 36414 220226
rect 36482 220170 36538 220226
rect 36606 220170 36662 220226
rect 36234 220046 36290 220102
rect 36358 220046 36414 220102
rect 36482 220046 36538 220102
rect 36606 220046 36662 220102
rect 36234 219922 36290 219978
rect 36358 219922 36414 219978
rect 36482 219922 36538 219978
rect 36606 219922 36662 219978
rect 39954 598116 40010 598172
rect 40078 598116 40134 598172
rect 40202 598116 40258 598172
rect 40326 598116 40382 598172
rect 39954 597992 40010 598048
rect 40078 597992 40134 598048
rect 40202 597992 40258 598048
rect 40326 597992 40382 598048
rect 39954 597868 40010 597924
rect 40078 597868 40134 597924
rect 40202 597868 40258 597924
rect 40326 597868 40382 597924
rect 39954 597744 40010 597800
rect 40078 597744 40134 597800
rect 40202 597744 40258 597800
rect 40326 597744 40382 597800
rect 39954 586294 40010 586350
rect 40078 586294 40134 586350
rect 40202 586294 40258 586350
rect 40326 586294 40382 586350
rect 39954 586170 40010 586226
rect 40078 586170 40134 586226
rect 40202 586170 40258 586226
rect 40326 586170 40382 586226
rect 39954 586046 40010 586102
rect 40078 586046 40134 586102
rect 40202 586046 40258 586102
rect 40326 586046 40382 586102
rect 39954 585922 40010 585978
rect 40078 585922 40134 585978
rect 40202 585922 40258 585978
rect 40326 585922 40382 585978
rect 39954 568294 40010 568350
rect 40078 568294 40134 568350
rect 40202 568294 40258 568350
rect 40326 568294 40382 568350
rect 39954 568170 40010 568226
rect 40078 568170 40134 568226
rect 40202 568170 40258 568226
rect 40326 568170 40382 568226
rect 39954 568046 40010 568102
rect 40078 568046 40134 568102
rect 40202 568046 40258 568102
rect 40326 568046 40382 568102
rect 39954 567922 40010 567978
rect 40078 567922 40134 567978
rect 40202 567922 40258 567978
rect 40326 567922 40382 567978
rect 39954 550294 40010 550350
rect 40078 550294 40134 550350
rect 40202 550294 40258 550350
rect 40326 550294 40382 550350
rect 39954 550170 40010 550226
rect 40078 550170 40134 550226
rect 40202 550170 40258 550226
rect 40326 550170 40382 550226
rect 39954 550046 40010 550102
rect 40078 550046 40134 550102
rect 40202 550046 40258 550102
rect 40326 550046 40382 550102
rect 39954 549922 40010 549978
rect 40078 549922 40134 549978
rect 40202 549922 40258 549978
rect 40326 549922 40382 549978
rect 39954 532294 40010 532350
rect 40078 532294 40134 532350
rect 40202 532294 40258 532350
rect 40326 532294 40382 532350
rect 39954 532170 40010 532226
rect 40078 532170 40134 532226
rect 40202 532170 40258 532226
rect 40326 532170 40382 532226
rect 39954 532046 40010 532102
rect 40078 532046 40134 532102
rect 40202 532046 40258 532102
rect 40326 532046 40382 532102
rect 39954 531922 40010 531978
rect 40078 531922 40134 531978
rect 40202 531922 40258 531978
rect 40326 531922 40382 531978
rect 66954 597156 67010 597212
rect 67078 597156 67134 597212
rect 67202 597156 67258 597212
rect 67326 597156 67382 597212
rect 66954 597032 67010 597088
rect 67078 597032 67134 597088
rect 67202 597032 67258 597088
rect 67326 597032 67382 597088
rect 66954 596908 67010 596964
rect 67078 596908 67134 596964
rect 67202 596908 67258 596964
rect 67326 596908 67382 596964
rect 66954 596784 67010 596840
rect 67078 596784 67134 596840
rect 67202 596784 67258 596840
rect 67326 596784 67382 596840
rect 66954 580294 67010 580350
rect 67078 580294 67134 580350
rect 67202 580294 67258 580350
rect 67326 580294 67382 580350
rect 66954 580170 67010 580226
rect 67078 580170 67134 580226
rect 67202 580170 67258 580226
rect 67326 580170 67382 580226
rect 66954 580046 67010 580102
rect 67078 580046 67134 580102
rect 67202 580046 67258 580102
rect 67326 580046 67382 580102
rect 66954 579922 67010 579978
rect 67078 579922 67134 579978
rect 67202 579922 67258 579978
rect 67326 579922 67382 579978
rect 66954 562294 67010 562350
rect 67078 562294 67134 562350
rect 67202 562294 67258 562350
rect 67326 562294 67382 562350
rect 66954 562170 67010 562226
rect 67078 562170 67134 562226
rect 67202 562170 67258 562226
rect 67326 562170 67382 562226
rect 66954 562046 67010 562102
rect 67078 562046 67134 562102
rect 67202 562046 67258 562102
rect 67326 562046 67382 562102
rect 66954 561922 67010 561978
rect 67078 561922 67134 561978
rect 67202 561922 67258 561978
rect 67326 561922 67382 561978
rect 66954 544294 67010 544350
rect 67078 544294 67134 544350
rect 67202 544294 67258 544350
rect 67326 544294 67382 544350
rect 66954 544170 67010 544226
rect 67078 544170 67134 544226
rect 67202 544170 67258 544226
rect 67326 544170 67382 544226
rect 66954 544046 67010 544102
rect 67078 544046 67134 544102
rect 67202 544046 67258 544102
rect 67326 544046 67382 544102
rect 66954 543922 67010 543978
rect 67078 543922 67134 543978
rect 67202 543922 67258 543978
rect 67326 543922 67382 543978
rect 70674 598116 70730 598172
rect 70798 598116 70854 598172
rect 70922 598116 70978 598172
rect 71046 598116 71102 598172
rect 70674 597992 70730 598048
rect 70798 597992 70854 598048
rect 70922 597992 70978 598048
rect 71046 597992 71102 598048
rect 70674 597868 70730 597924
rect 70798 597868 70854 597924
rect 70922 597868 70978 597924
rect 71046 597868 71102 597924
rect 70674 597744 70730 597800
rect 70798 597744 70854 597800
rect 70922 597744 70978 597800
rect 71046 597744 71102 597800
rect 70674 586294 70730 586350
rect 70798 586294 70854 586350
rect 70922 586294 70978 586350
rect 71046 586294 71102 586350
rect 70674 586170 70730 586226
rect 70798 586170 70854 586226
rect 70922 586170 70978 586226
rect 71046 586170 71102 586226
rect 70674 586046 70730 586102
rect 70798 586046 70854 586102
rect 70922 586046 70978 586102
rect 71046 586046 71102 586102
rect 70674 585922 70730 585978
rect 70798 585922 70854 585978
rect 70922 585922 70978 585978
rect 71046 585922 71102 585978
rect 70674 568294 70730 568350
rect 70798 568294 70854 568350
rect 70922 568294 70978 568350
rect 71046 568294 71102 568350
rect 70674 568170 70730 568226
rect 70798 568170 70854 568226
rect 70922 568170 70978 568226
rect 71046 568170 71102 568226
rect 70674 568046 70730 568102
rect 70798 568046 70854 568102
rect 70922 568046 70978 568102
rect 71046 568046 71102 568102
rect 70674 567922 70730 567978
rect 70798 567922 70854 567978
rect 70922 567922 70978 567978
rect 71046 567922 71102 567978
rect 70674 550294 70730 550350
rect 70798 550294 70854 550350
rect 70922 550294 70978 550350
rect 71046 550294 71102 550350
rect 70674 550170 70730 550226
rect 70798 550170 70854 550226
rect 70922 550170 70978 550226
rect 71046 550170 71102 550226
rect 70674 550046 70730 550102
rect 70798 550046 70854 550102
rect 70922 550046 70978 550102
rect 71046 550046 71102 550102
rect 70674 549922 70730 549978
rect 70798 549922 70854 549978
rect 70922 549922 70978 549978
rect 71046 549922 71102 549978
rect 97674 597156 97730 597212
rect 97798 597156 97854 597212
rect 97922 597156 97978 597212
rect 98046 597156 98102 597212
rect 97674 597032 97730 597088
rect 97798 597032 97854 597088
rect 97922 597032 97978 597088
rect 98046 597032 98102 597088
rect 97674 596908 97730 596964
rect 97798 596908 97854 596964
rect 97922 596908 97978 596964
rect 98046 596908 98102 596964
rect 97674 596784 97730 596840
rect 97798 596784 97854 596840
rect 97922 596784 97978 596840
rect 98046 596784 98102 596840
rect 97674 580294 97730 580350
rect 97798 580294 97854 580350
rect 97922 580294 97978 580350
rect 98046 580294 98102 580350
rect 97674 580170 97730 580226
rect 97798 580170 97854 580226
rect 97922 580170 97978 580226
rect 98046 580170 98102 580226
rect 97674 580046 97730 580102
rect 97798 580046 97854 580102
rect 97922 580046 97978 580102
rect 98046 580046 98102 580102
rect 97674 579922 97730 579978
rect 97798 579922 97854 579978
rect 97922 579922 97978 579978
rect 98046 579922 98102 579978
rect 97674 562294 97730 562350
rect 97798 562294 97854 562350
rect 97922 562294 97978 562350
rect 98046 562294 98102 562350
rect 97674 562170 97730 562226
rect 97798 562170 97854 562226
rect 97922 562170 97978 562226
rect 98046 562170 98102 562226
rect 97674 562046 97730 562102
rect 97798 562046 97854 562102
rect 97922 562046 97978 562102
rect 98046 562046 98102 562102
rect 97674 561922 97730 561978
rect 97798 561922 97854 561978
rect 97922 561922 97978 561978
rect 98046 561922 98102 561978
rect 97674 544294 97730 544350
rect 97798 544294 97854 544350
rect 97922 544294 97978 544350
rect 98046 544294 98102 544350
rect 97674 544170 97730 544226
rect 97798 544170 97854 544226
rect 97922 544170 97978 544226
rect 98046 544170 98102 544226
rect 97674 544046 97730 544102
rect 97798 544046 97854 544102
rect 97922 544046 97978 544102
rect 98046 544046 98102 544102
rect 97674 543922 97730 543978
rect 97798 543922 97854 543978
rect 97922 543922 97978 543978
rect 98046 543922 98102 543978
rect 101394 598116 101450 598172
rect 101518 598116 101574 598172
rect 101642 598116 101698 598172
rect 101766 598116 101822 598172
rect 101394 597992 101450 598048
rect 101518 597992 101574 598048
rect 101642 597992 101698 598048
rect 101766 597992 101822 598048
rect 101394 597868 101450 597924
rect 101518 597868 101574 597924
rect 101642 597868 101698 597924
rect 101766 597868 101822 597924
rect 101394 597744 101450 597800
rect 101518 597744 101574 597800
rect 101642 597744 101698 597800
rect 101766 597744 101822 597800
rect 101394 586294 101450 586350
rect 101518 586294 101574 586350
rect 101642 586294 101698 586350
rect 101766 586294 101822 586350
rect 101394 586170 101450 586226
rect 101518 586170 101574 586226
rect 101642 586170 101698 586226
rect 101766 586170 101822 586226
rect 101394 586046 101450 586102
rect 101518 586046 101574 586102
rect 101642 586046 101698 586102
rect 101766 586046 101822 586102
rect 101394 585922 101450 585978
rect 101518 585922 101574 585978
rect 101642 585922 101698 585978
rect 101766 585922 101822 585978
rect 101394 568294 101450 568350
rect 101518 568294 101574 568350
rect 101642 568294 101698 568350
rect 101766 568294 101822 568350
rect 101394 568170 101450 568226
rect 101518 568170 101574 568226
rect 101642 568170 101698 568226
rect 101766 568170 101822 568226
rect 101394 568046 101450 568102
rect 101518 568046 101574 568102
rect 101642 568046 101698 568102
rect 101766 568046 101822 568102
rect 101394 567922 101450 567978
rect 101518 567922 101574 567978
rect 101642 567922 101698 567978
rect 101766 567922 101822 567978
rect 128394 597156 128450 597212
rect 128518 597156 128574 597212
rect 128642 597156 128698 597212
rect 128766 597156 128822 597212
rect 128394 597032 128450 597088
rect 128518 597032 128574 597088
rect 128642 597032 128698 597088
rect 128766 597032 128822 597088
rect 128394 596908 128450 596964
rect 128518 596908 128574 596964
rect 128642 596908 128698 596964
rect 128766 596908 128822 596964
rect 128394 596784 128450 596840
rect 128518 596784 128574 596840
rect 128642 596784 128698 596840
rect 128766 596784 128822 596840
rect 128394 580294 128450 580350
rect 128518 580294 128574 580350
rect 128642 580294 128698 580350
rect 128766 580294 128822 580350
rect 128394 580170 128450 580226
rect 128518 580170 128574 580226
rect 128642 580170 128698 580226
rect 128766 580170 128822 580226
rect 128394 580046 128450 580102
rect 128518 580046 128574 580102
rect 128642 580046 128698 580102
rect 128766 580046 128822 580102
rect 128394 579922 128450 579978
rect 128518 579922 128574 579978
rect 128642 579922 128698 579978
rect 128766 579922 128822 579978
rect 128394 562294 128450 562350
rect 128518 562294 128574 562350
rect 128642 562294 128698 562350
rect 128766 562294 128822 562350
rect 128394 562170 128450 562226
rect 128518 562170 128574 562226
rect 128642 562170 128698 562226
rect 128766 562170 128822 562226
rect 128394 562046 128450 562102
rect 128518 562046 128574 562102
rect 128642 562046 128698 562102
rect 128766 562046 128822 562102
rect 117336 561932 117392 561988
rect 117460 561932 117516 561988
rect 117584 561932 117640 561988
rect 117708 561932 117764 561988
rect 117832 561932 117888 561988
rect 117956 561932 118012 561988
rect 118080 561932 118136 561988
rect 118204 561932 118260 561988
rect 118328 561932 118384 561988
rect 118452 561932 118508 561988
rect 118576 561932 118632 561988
rect 118700 561932 118756 561988
rect 118824 561932 118880 561988
rect 118948 561932 119004 561988
rect 119072 561932 119128 561988
rect 119196 561932 119252 561988
rect 119320 561932 119376 561988
rect 119444 561932 119500 561988
rect 119568 561932 119624 561988
rect 119692 561932 119748 561988
rect 119816 561932 119872 561988
rect 119940 561932 119996 561988
rect 120064 561932 120120 561988
rect 120188 561932 120244 561988
rect 120312 561932 120368 561988
rect 120436 561932 120492 561988
rect 120560 561932 120616 561988
rect 120684 561932 120740 561988
rect 120808 561932 120864 561988
rect 120932 561932 120988 561988
rect 121056 561932 121112 561988
rect 121180 561932 121236 561988
rect 121304 561932 121360 561988
rect 121428 561932 121484 561988
rect 121552 561932 121608 561988
rect 121676 561932 121732 561988
rect 121800 561932 121856 561988
rect 121924 561932 121980 561988
rect 122048 561932 122104 561988
rect 122172 561932 122228 561988
rect 122296 561932 122352 561988
rect 122420 561932 122476 561988
rect 122544 561932 122600 561988
rect 122668 561932 122724 561988
rect 122792 561932 122848 561988
rect 122916 561932 122972 561988
rect 123040 561932 123096 561988
rect 123164 561932 123220 561988
rect 123288 561932 123344 561988
rect 123412 561932 123468 561988
rect 123536 561932 123592 561988
rect 123660 561932 123716 561988
rect 123784 561932 123840 561988
rect 123908 561932 123964 561988
rect 124032 561932 124088 561988
rect 124156 561932 124212 561988
rect 124280 561932 124336 561988
rect 124404 561932 124460 561988
rect 124528 561932 124584 561988
rect 128394 561922 128450 561978
rect 128518 561922 128574 561978
rect 128642 561922 128698 561978
rect 128766 561922 128822 561978
rect 101394 550294 101450 550350
rect 101518 550294 101574 550350
rect 101642 550294 101698 550350
rect 101766 550294 101822 550350
rect 101394 550170 101450 550226
rect 101518 550170 101574 550226
rect 101642 550170 101698 550226
rect 101766 550170 101822 550226
rect 101394 550046 101450 550102
rect 101518 550046 101574 550102
rect 101642 550046 101698 550102
rect 101766 550046 101822 550102
rect 101394 549922 101450 549978
rect 101518 549922 101574 549978
rect 101642 549922 101698 549978
rect 101766 549922 101822 549978
rect 128394 544294 128450 544350
rect 128518 544294 128574 544350
rect 128642 544294 128698 544350
rect 128766 544294 128822 544350
rect 128394 544170 128450 544226
rect 128518 544170 128574 544226
rect 128642 544170 128698 544226
rect 128766 544170 128822 544226
rect 104066 544007 104122 544063
rect 104190 544007 104246 544063
rect 104314 544007 104370 544063
rect 104438 544007 104494 544063
rect 104562 544007 104618 544063
rect 104686 544007 104742 544063
rect 104810 544007 104866 544063
rect 104934 544007 104990 544063
rect 105058 544007 105114 544063
rect 105182 544007 105238 544063
rect 105306 544007 105362 544063
rect 105430 544007 105486 544063
rect 105554 544007 105610 544063
rect 105678 544007 105734 544063
rect 105802 544007 105858 544063
rect 105926 544007 105982 544063
rect 106050 544007 106106 544063
rect 106174 544007 106230 544063
rect 106298 544007 106354 544063
rect 106422 544007 106478 544063
rect 106546 544007 106602 544063
rect 106670 544007 106726 544063
rect 106794 544007 106850 544063
rect 106918 544007 106974 544063
rect 107042 544007 107098 544063
rect 107166 544007 107222 544063
rect 107290 544007 107346 544063
rect 107414 544007 107470 544063
rect 107538 544007 107594 544063
rect 107662 544007 107718 544063
rect 107786 544007 107842 544063
rect 107910 544007 107966 544063
rect 108034 544007 108090 544063
rect 108158 544007 108214 544063
rect 108282 544007 108338 544063
rect 108406 544007 108462 544063
rect 108530 544007 108586 544063
rect 108654 544007 108710 544063
rect 108778 544007 108834 544063
rect 108902 544007 108958 544063
rect 109026 544007 109082 544063
rect 109150 544007 109206 544063
rect 109274 544007 109330 544063
rect 109398 544007 109454 544063
rect 109522 544007 109578 544063
rect 109646 544007 109702 544063
rect 109770 544007 109826 544063
rect 109894 544007 109950 544063
rect 110018 544007 110074 544063
rect 110142 544007 110198 544063
rect 110266 544007 110322 544063
rect 110390 544007 110446 544063
rect 110514 544007 110570 544063
rect 110638 544007 110694 544063
rect 110762 544007 110818 544063
rect 110886 544007 110942 544063
rect 111010 544007 111066 544063
rect 111134 544007 111190 544063
rect 111258 544007 111314 544063
rect 111382 544007 111438 544063
rect 111506 544007 111562 544063
rect 111630 544007 111686 544063
rect 111754 544007 111810 544063
rect 111878 544007 111934 544063
rect 112002 544007 112058 544063
rect 112126 544007 112182 544063
rect 112250 544007 112306 544063
rect 112374 544007 112430 544063
rect 112498 544007 112554 544063
rect 112622 544007 112678 544063
rect 112746 544007 112802 544063
rect 112870 544007 112926 544063
rect 112994 544007 113050 544063
rect 113118 544007 113174 544063
rect 113242 544007 113298 544063
rect 113366 544007 113422 544063
rect 113490 544007 113546 544063
rect 113614 544007 113670 544063
rect 113738 544007 113794 544063
rect 113862 544007 113918 544063
rect 113986 544007 114042 544063
rect 114110 544007 114166 544063
rect 114234 544007 114290 544063
rect 114358 544007 114414 544063
rect 114482 544007 114538 544063
rect 114606 544007 114662 544063
rect 114730 544007 114786 544063
rect 114854 544007 114910 544063
rect 114978 544007 115034 544063
rect 115102 544007 115158 544063
rect 115226 544007 115282 544063
rect 115350 544007 115406 544063
rect 115474 544007 115530 544063
rect 115598 544007 115654 544063
rect 115722 544007 115778 544063
rect 115846 544007 115902 544063
rect 115970 544007 116026 544063
rect 116094 544007 116150 544063
rect 116218 544007 116274 544063
rect 116342 544007 116398 544063
rect 116466 544007 116522 544063
rect 116590 544007 116646 544063
rect 116714 544007 116770 544063
rect 116838 544007 116894 544063
rect 116962 544007 117018 544063
rect 117086 544007 117142 544063
rect 117210 544007 117266 544063
rect 117334 544007 117390 544063
rect 117458 544007 117514 544063
rect 117582 544007 117638 544063
rect 117706 544007 117762 544063
rect 117830 544007 117886 544063
rect 117954 544007 118010 544063
rect 118078 544007 118134 544063
rect 118202 544007 118258 544063
rect 118326 544007 118382 544063
rect 118450 544007 118506 544063
rect 118574 544007 118630 544063
rect 118698 544007 118754 544063
rect 118822 544007 118878 544063
rect 118946 544007 119002 544063
rect 119070 544007 119126 544063
rect 119194 544007 119250 544063
rect 119318 544007 119374 544063
rect 119442 544007 119498 544063
rect 119566 544007 119622 544063
rect 119690 544007 119746 544063
rect 119814 544007 119870 544063
rect 119938 544007 119994 544063
rect 120062 544007 120118 544063
rect 120186 544007 120242 544063
rect 120310 544007 120366 544063
rect 120434 544007 120490 544063
rect 120558 544007 120614 544063
rect 120682 544007 120738 544063
rect 120806 544007 120862 544063
rect 120930 544007 120986 544063
rect 121054 544007 121110 544063
rect 121178 544007 121234 544063
rect 121302 544007 121358 544063
rect 121426 544007 121482 544063
rect 121550 544007 121606 544063
rect 121674 544007 121730 544063
rect 121798 544007 121854 544063
rect 104066 543883 104122 543939
rect 104190 543883 104246 543939
rect 104314 543883 104370 543939
rect 104438 543883 104494 543939
rect 104562 543883 104618 543939
rect 104686 543883 104742 543939
rect 104810 543883 104866 543939
rect 104934 543883 104990 543939
rect 105058 543883 105114 543939
rect 105182 543883 105238 543939
rect 105306 543883 105362 543939
rect 105430 543883 105486 543939
rect 105554 543883 105610 543939
rect 105678 543883 105734 543939
rect 105802 543883 105858 543939
rect 105926 543883 105982 543939
rect 106050 543883 106106 543939
rect 106174 543883 106230 543939
rect 106298 543883 106354 543939
rect 106422 543883 106478 543939
rect 106546 543883 106602 543939
rect 106670 543883 106726 543939
rect 106794 543883 106850 543939
rect 106918 543883 106974 543939
rect 107042 543883 107098 543939
rect 107166 543883 107222 543939
rect 107290 543883 107346 543939
rect 107414 543883 107470 543939
rect 107538 543883 107594 543939
rect 107662 543883 107718 543939
rect 107786 543883 107842 543939
rect 107910 543883 107966 543939
rect 108034 543883 108090 543939
rect 108158 543883 108214 543939
rect 108282 543883 108338 543939
rect 108406 543883 108462 543939
rect 108530 543883 108586 543939
rect 108654 543883 108710 543939
rect 108778 543883 108834 543939
rect 108902 543883 108958 543939
rect 109026 543883 109082 543939
rect 109150 543883 109206 543939
rect 109274 543883 109330 543939
rect 109398 543883 109454 543939
rect 109522 543883 109578 543939
rect 109646 543883 109702 543939
rect 109770 543883 109826 543939
rect 109894 543883 109950 543939
rect 110018 543883 110074 543939
rect 110142 543883 110198 543939
rect 110266 543883 110322 543939
rect 110390 543883 110446 543939
rect 110514 543883 110570 543939
rect 110638 543883 110694 543939
rect 110762 543883 110818 543939
rect 110886 543883 110942 543939
rect 111010 543883 111066 543939
rect 111134 543883 111190 543939
rect 111258 543883 111314 543939
rect 111382 543883 111438 543939
rect 111506 543883 111562 543939
rect 111630 543883 111686 543939
rect 111754 543883 111810 543939
rect 111878 543883 111934 543939
rect 112002 543883 112058 543939
rect 112126 543883 112182 543939
rect 112250 543883 112306 543939
rect 112374 543883 112430 543939
rect 112498 543883 112554 543939
rect 112622 543883 112678 543939
rect 112746 543883 112802 543939
rect 112870 543883 112926 543939
rect 112994 543883 113050 543939
rect 113118 543883 113174 543939
rect 113242 543883 113298 543939
rect 113366 543883 113422 543939
rect 113490 543883 113546 543939
rect 113614 543883 113670 543939
rect 113738 543883 113794 543939
rect 113862 543883 113918 543939
rect 113986 543883 114042 543939
rect 114110 543883 114166 543939
rect 114234 543883 114290 543939
rect 114358 543883 114414 543939
rect 114482 543883 114538 543939
rect 114606 543883 114662 543939
rect 114730 543883 114786 543939
rect 114854 543883 114910 543939
rect 114978 543883 115034 543939
rect 115102 543883 115158 543939
rect 115226 543883 115282 543939
rect 115350 543883 115406 543939
rect 115474 543883 115530 543939
rect 115598 543883 115654 543939
rect 115722 543883 115778 543939
rect 115846 543883 115902 543939
rect 115970 543883 116026 543939
rect 116094 543883 116150 543939
rect 116218 543883 116274 543939
rect 116342 543883 116398 543939
rect 116466 543883 116522 543939
rect 116590 543883 116646 543939
rect 116714 543883 116770 543939
rect 116838 543883 116894 543939
rect 116962 543883 117018 543939
rect 117086 543883 117142 543939
rect 117210 543883 117266 543939
rect 117334 543883 117390 543939
rect 117458 543883 117514 543939
rect 117582 543883 117638 543939
rect 117706 543883 117762 543939
rect 117830 543883 117886 543939
rect 117954 543883 118010 543939
rect 118078 543883 118134 543939
rect 118202 543883 118258 543939
rect 118326 543883 118382 543939
rect 118450 543883 118506 543939
rect 118574 543883 118630 543939
rect 118698 543883 118754 543939
rect 118822 543883 118878 543939
rect 118946 543883 119002 543939
rect 119070 543883 119126 543939
rect 119194 543883 119250 543939
rect 119318 543883 119374 543939
rect 119442 543883 119498 543939
rect 119566 543883 119622 543939
rect 119690 543883 119746 543939
rect 119814 543883 119870 543939
rect 119938 543883 119994 543939
rect 120062 543883 120118 543939
rect 120186 543883 120242 543939
rect 120310 543883 120366 543939
rect 120434 543883 120490 543939
rect 120558 543883 120614 543939
rect 120682 543883 120738 543939
rect 120806 543883 120862 543939
rect 120930 543883 120986 543939
rect 121054 543883 121110 543939
rect 121178 543883 121234 543939
rect 121302 543883 121358 543939
rect 121426 543883 121482 543939
rect 121550 543883 121606 543939
rect 121674 543883 121730 543939
rect 121798 543883 121854 543939
rect 128394 544046 128450 544102
rect 128518 544046 128574 544102
rect 128642 544046 128698 544102
rect 128766 544046 128822 544102
rect 128394 543922 128450 543978
rect 128518 543922 128574 543978
rect 128642 543922 128698 543978
rect 128766 543922 128822 543978
rect 132114 598116 132170 598172
rect 132238 598116 132294 598172
rect 132362 598116 132418 598172
rect 132486 598116 132542 598172
rect 132114 597992 132170 598048
rect 132238 597992 132294 598048
rect 132362 597992 132418 598048
rect 132486 597992 132542 598048
rect 132114 597868 132170 597924
rect 132238 597868 132294 597924
rect 132362 597868 132418 597924
rect 132486 597868 132542 597924
rect 132114 597744 132170 597800
rect 132238 597744 132294 597800
rect 132362 597744 132418 597800
rect 132486 597744 132542 597800
rect 132114 586294 132170 586350
rect 132238 586294 132294 586350
rect 132362 586294 132418 586350
rect 132486 586294 132542 586350
rect 132114 586170 132170 586226
rect 132238 586170 132294 586226
rect 132362 586170 132418 586226
rect 132486 586170 132542 586226
rect 132114 586046 132170 586102
rect 132238 586046 132294 586102
rect 132362 586046 132418 586102
rect 132486 586046 132542 586102
rect 132114 585922 132170 585978
rect 132238 585922 132294 585978
rect 132362 585922 132418 585978
rect 132486 585922 132542 585978
rect 132114 568294 132170 568350
rect 132238 568294 132294 568350
rect 132362 568294 132418 568350
rect 132486 568294 132542 568350
rect 132114 568170 132170 568226
rect 132238 568170 132294 568226
rect 132362 568170 132418 568226
rect 132486 568170 132542 568226
rect 132114 568046 132170 568102
rect 132238 568046 132294 568102
rect 132362 568046 132418 568102
rect 132486 568046 132542 568102
rect 132114 567922 132170 567978
rect 132238 567922 132294 567978
rect 132362 567922 132418 567978
rect 132486 567922 132542 567978
rect 132114 550294 132170 550350
rect 132238 550294 132294 550350
rect 132362 550294 132418 550350
rect 132486 550294 132542 550350
rect 132114 550170 132170 550226
rect 132238 550170 132294 550226
rect 132362 550170 132418 550226
rect 132486 550170 132542 550226
rect 132114 550046 132170 550102
rect 132238 550046 132294 550102
rect 132362 550046 132418 550102
rect 132486 550046 132542 550102
rect 132114 549922 132170 549978
rect 132238 549922 132294 549978
rect 132362 549922 132418 549978
rect 132486 549922 132542 549978
rect 159114 597156 159170 597212
rect 159238 597156 159294 597212
rect 159362 597156 159418 597212
rect 159486 597156 159542 597212
rect 159114 597032 159170 597088
rect 159238 597032 159294 597088
rect 159362 597032 159418 597088
rect 159486 597032 159542 597088
rect 159114 596908 159170 596964
rect 159238 596908 159294 596964
rect 159362 596908 159418 596964
rect 159486 596908 159542 596964
rect 159114 596784 159170 596840
rect 159238 596784 159294 596840
rect 159362 596784 159418 596840
rect 159486 596784 159542 596840
rect 159114 580294 159170 580350
rect 159238 580294 159294 580350
rect 159362 580294 159418 580350
rect 159486 580294 159542 580350
rect 159114 580170 159170 580226
rect 159238 580170 159294 580226
rect 159362 580170 159418 580226
rect 159486 580170 159542 580226
rect 159114 580046 159170 580102
rect 159238 580046 159294 580102
rect 159362 580046 159418 580102
rect 159486 580046 159542 580102
rect 159114 579922 159170 579978
rect 159238 579922 159294 579978
rect 159362 579922 159418 579978
rect 159486 579922 159542 579978
rect 159114 562294 159170 562350
rect 159238 562294 159294 562350
rect 159362 562294 159418 562350
rect 159486 562294 159542 562350
rect 159114 562170 159170 562226
rect 159238 562170 159294 562226
rect 159362 562170 159418 562226
rect 159486 562170 159542 562226
rect 159114 562046 159170 562102
rect 159238 562046 159294 562102
rect 159362 562046 159418 562102
rect 159486 562046 159542 562102
rect 159114 561922 159170 561978
rect 159238 561922 159294 561978
rect 159362 561922 159418 561978
rect 159486 561922 159542 561978
rect 159114 544294 159170 544350
rect 159238 544294 159294 544350
rect 159362 544294 159418 544350
rect 159486 544294 159542 544350
rect 159114 544170 159170 544226
rect 159238 544170 159294 544226
rect 159362 544170 159418 544226
rect 159486 544170 159542 544226
rect 159114 544046 159170 544102
rect 159238 544046 159294 544102
rect 159362 544046 159418 544102
rect 159486 544046 159542 544102
rect 159114 543922 159170 543978
rect 159238 543922 159294 543978
rect 159362 543922 159418 543978
rect 159486 543922 159542 543978
rect 71876 532332 71932 532388
rect 72000 532332 72056 532388
rect 72124 532332 72180 532388
rect 72248 532332 72304 532388
rect 72372 532332 72428 532388
rect 72496 532332 72552 532388
rect 72620 532332 72676 532388
rect 72744 532332 72800 532388
rect 72868 532332 72924 532388
rect 72992 532332 73048 532388
rect 73116 532332 73172 532388
rect 73240 532332 73296 532388
rect 73364 532332 73420 532388
rect 73488 532332 73544 532388
rect 73612 532332 73668 532388
rect 73736 532332 73792 532388
rect 73860 532332 73916 532388
rect 73984 532332 74040 532388
rect 74108 532332 74164 532388
rect 74232 532332 74288 532388
rect 74356 532332 74412 532388
rect 74480 532332 74536 532388
rect 74604 532332 74660 532388
rect 74728 532332 74784 532388
rect 74852 532332 74908 532388
rect 74976 532332 75032 532388
rect 75100 532332 75156 532388
rect 75224 532332 75280 532388
rect 75348 532332 75404 532388
rect 75472 532332 75528 532388
rect 75596 532332 75652 532388
rect 75720 532332 75776 532388
rect 75844 532332 75900 532388
rect 75968 532332 76024 532388
rect 76092 532332 76148 532388
rect 76216 532332 76272 532388
rect 76340 532332 76396 532388
rect 76464 532332 76520 532388
rect 76588 532332 76644 532388
rect 76712 532332 76768 532388
rect 76836 532332 76892 532388
rect 76960 532332 77016 532388
rect 77084 532332 77140 532388
rect 77208 532332 77264 532388
rect 77332 532332 77388 532388
rect 77456 532332 77512 532388
rect 77580 532332 77636 532388
rect 77704 532332 77760 532388
rect 77828 532332 77884 532388
rect 77952 532332 78008 532388
rect 78076 532332 78132 532388
rect 78200 532332 78256 532388
rect 78324 532332 78380 532388
rect 78448 532332 78504 532388
rect 78572 532332 78628 532388
rect 78696 532332 78752 532388
rect 78820 532332 78876 532388
rect 78944 532332 79000 532388
rect 79068 532332 79124 532388
rect 79192 532332 79248 532388
rect 79316 532332 79372 532388
rect 79440 532332 79496 532388
rect 79564 532332 79620 532388
rect 79688 532332 79744 532388
rect 79812 532332 79868 532388
rect 79936 532332 79992 532388
rect 80060 532332 80116 532388
rect 80184 532332 80240 532388
rect 80308 532332 80364 532388
rect 80432 532332 80488 532388
rect 80556 532332 80612 532388
rect 80680 532332 80736 532388
rect 80804 532332 80860 532388
rect 80928 532332 80984 532388
rect 81052 532332 81108 532388
rect 81176 532332 81232 532388
rect 81300 532332 81356 532388
rect 81424 532332 81480 532388
rect 81548 532332 81604 532388
rect 81672 532332 81728 532388
rect 81796 532332 81852 532388
rect 81920 532332 81976 532388
rect 82044 532332 82100 532388
rect 82168 532332 82224 532388
rect 82292 532332 82348 532388
rect 82416 532332 82472 532388
rect 82540 532332 82596 532388
rect 82664 532332 82720 532388
rect 82788 532332 82844 532388
rect 159114 526294 159170 526350
rect 159238 526294 159294 526350
rect 159362 526294 159418 526350
rect 159486 526294 159542 526350
rect 94310 526092 94366 526148
rect 94434 526092 94490 526148
rect 94558 526092 94614 526148
rect 94682 526092 94738 526148
rect 94806 526092 94862 526148
rect 94930 526092 94986 526148
rect 95054 526092 95110 526148
rect 95178 526092 95234 526148
rect 95302 526092 95358 526148
rect 95426 526092 95482 526148
rect 95550 526092 95606 526148
rect 95674 526092 95730 526148
rect 95798 526092 95854 526148
rect 95922 526092 95978 526148
rect 96046 526092 96102 526148
rect 96170 526092 96226 526148
rect 96294 526092 96350 526148
rect 96418 526092 96474 526148
rect 96542 526092 96598 526148
rect 96666 526092 96722 526148
rect 96790 526092 96846 526148
rect 96914 526092 96970 526148
rect 97038 526092 97094 526148
rect 97162 526092 97218 526148
rect 97286 526092 97342 526148
rect 97410 526092 97466 526148
rect 97534 526092 97590 526148
rect 97658 526092 97714 526148
rect 97782 526092 97838 526148
rect 97906 526092 97962 526148
rect 98030 526092 98086 526148
rect 98154 526092 98210 526148
rect 98278 526092 98334 526148
rect 98402 526092 98458 526148
rect 98526 526092 98582 526148
rect 98650 526092 98706 526148
rect 98774 526092 98830 526148
rect 98898 526092 98954 526148
rect 99022 526092 99078 526148
rect 99146 526092 99202 526148
rect 99270 526092 99326 526148
rect 99394 526092 99450 526148
rect 99518 526092 99574 526148
rect 99642 526092 99698 526148
rect 99766 526092 99822 526148
rect 99890 526092 99946 526148
rect 100014 526092 100070 526148
rect 100138 526092 100194 526148
rect 100262 526092 100318 526148
rect 100386 526092 100442 526148
rect 100510 526092 100566 526148
rect 100634 526092 100690 526148
rect 100758 526092 100814 526148
rect 100882 526092 100938 526148
rect 101006 526092 101062 526148
rect 101130 526092 101186 526148
rect 101254 526092 101310 526148
rect 101378 526092 101434 526148
rect 101502 526092 101558 526148
rect 101626 526092 101682 526148
rect 101750 526092 101806 526148
rect 101874 526092 101930 526148
rect 101998 526092 102054 526148
rect 102122 526092 102178 526148
rect 102246 526092 102302 526148
rect 102370 526092 102426 526148
rect 102494 526092 102550 526148
rect 102618 526092 102674 526148
rect 102742 526092 102798 526148
rect 102866 526092 102922 526148
rect 102990 526092 103046 526148
rect 103114 526092 103170 526148
rect 103238 526092 103294 526148
rect 103362 526092 103418 526148
rect 103486 526092 103542 526148
rect 103610 526092 103666 526148
rect 103734 526092 103790 526148
rect 103858 526092 103914 526148
rect 103982 526092 104038 526148
rect 104106 526092 104162 526148
rect 104230 526092 104286 526148
rect 104354 526092 104410 526148
rect 104478 526092 104534 526148
rect 104602 526092 104658 526148
rect 104726 526092 104782 526148
rect 104850 526092 104906 526148
rect 104974 526092 105030 526148
rect 105098 526092 105154 526148
rect 105222 526092 105278 526148
rect 105346 526092 105402 526148
rect 105470 526092 105526 526148
rect 105594 526092 105650 526148
rect 105718 526092 105774 526148
rect 105842 526092 105898 526148
rect 105966 526092 106022 526148
rect 106090 526092 106146 526148
rect 106214 526092 106270 526148
rect 106338 526092 106394 526148
rect 106462 526092 106518 526148
rect 106586 526092 106642 526148
rect 106710 526092 106766 526148
rect 106834 526092 106890 526148
rect 106958 526092 107014 526148
rect 107082 526092 107138 526148
rect 107206 526092 107262 526148
rect 107330 526092 107386 526148
rect 107454 526092 107510 526148
rect 107578 526092 107634 526148
rect 107702 526092 107758 526148
rect 107826 526092 107882 526148
rect 107950 526092 108006 526148
rect 108074 526092 108130 526148
rect 108198 526092 108254 526148
rect 108322 526092 108378 526148
rect 108446 526092 108502 526148
rect 108570 526092 108626 526148
rect 108694 526092 108750 526148
rect 108818 526092 108874 526148
rect 108942 526092 108998 526148
rect 109066 526092 109122 526148
rect 109190 526092 109246 526148
rect 109314 526092 109370 526148
rect 109438 526092 109494 526148
rect 109562 526092 109618 526148
rect 109686 526092 109742 526148
rect 109810 526092 109866 526148
rect 109934 526092 109990 526148
rect 110058 526092 110114 526148
rect 110182 526092 110238 526148
rect 110306 526092 110362 526148
rect 110430 526092 110486 526148
rect 110554 526092 110610 526148
rect 110678 526092 110734 526148
rect 110802 526092 110858 526148
rect 110926 526092 110982 526148
rect 111050 526092 111106 526148
rect 111174 526092 111230 526148
rect 111298 526092 111354 526148
rect 111422 526092 111478 526148
rect 111546 526092 111602 526148
rect 111670 526092 111726 526148
rect 111794 526092 111850 526148
rect 111918 526092 111974 526148
rect 112042 526092 112098 526148
rect 112166 526092 112222 526148
rect 112290 526092 112346 526148
rect 112414 526092 112470 526148
rect 112538 526092 112594 526148
rect 112662 526092 112718 526148
rect 112786 526092 112842 526148
rect 112910 526092 112966 526148
rect 113034 526092 113090 526148
rect 113158 526092 113214 526148
rect 113282 526092 113338 526148
rect 113406 526092 113462 526148
rect 113530 526092 113586 526148
rect 113654 526092 113710 526148
rect 113778 526092 113834 526148
rect 113902 526092 113958 526148
rect 114026 526092 114082 526148
rect 114150 526092 114206 526148
rect 114274 526092 114330 526148
rect 159114 526170 159170 526226
rect 159238 526170 159294 526226
rect 159362 526170 159418 526226
rect 159486 526170 159542 526226
rect 159114 526046 159170 526102
rect 159238 526046 159294 526102
rect 159362 526046 159418 526102
rect 159486 526046 159542 526102
rect 39954 514294 40010 514350
rect 40078 514294 40134 514350
rect 40202 514294 40258 514350
rect 40326 514294 40382 514350
rect 39954 514170 40010 514226
rect 40078 514170 40134 514226
rect 40202 514170 40258 514226
rect 40326 514170 40382 514226
rect 159114 525922 159170 525978
rect 159238 525922 159294 525978
rect 159362 525922 159418 525978
rect 159486 525922 159542 525978
rect 39954 514046 40010 514102
rect 40078 514046 40134 514102
rect 40202 514046 40258 514102
rect 40326 514046 40382 514102
rect 39954 513922 40010 513978
rect 40078 513922 40134 513978
rect 40202 513922 40258 513978
rect 40326 513922 40382 513978
rect 60844 514074 60900 514130
rect 60968 514074 61024 514130
rect 61092 514074 61148 514130
rect 61216 514074 61272 514130
rect 61340 514074 61396 514130
rect 61464 514074 61520 514130
rect 61588 514074 61644 514130
rect 61712 514074 61768 514130
rect 61836 514074 61892 514130
rect 61960 514074 62016 514130
rect 62084 514074 62140 514130
rect 62208 514074 62264 514130
rect 62332 514074 62388 514130
rect 62456 514074 62512 514130
rect 62580 514074 62636 514130
rect 62704 514074 62760 514130
rect 62828 514074 62884 514130
rect 62952 514074 63008 514130
rect 63076 514074 63132 514130
rect 63200 514074 63256 514130
rect 63324 514074 63380 514130
rect 63448 514074 63504 514130
rect 63572 514074 63628 514130
rect 63696 514074 63752 514130
rect 63820 514074 63876 514130
rect 63944 514074 64000 514130
rect 64068 514074 64124 514130
rect 64192 514074 64248 514130
rect 64316 514074 64372 514130
rect 64440 514074 64496 514130
rect 64564 514074 64620 514130
rect 64688 514074 64744 514130
rect 64812 514074 64868 514130
rect 64936 514074 64992 514130
rect 65060 514074 65116 514130
rect 65184 514074 65240 514130
rect 65308 514074 65364 514130
rect 65432 514074 65488 514130
rect 65556 514074 65612 514130
rect 65680 514074 65736 514130
rect 65804 514074 65860 514130
rect 65928 514074 65984 514130
rect 66052 514074 66108 514130
rect 66176 514074 66232 514130
rect 66300 514074 66356 514130
rect 60844 513950 60900 514006
rect 60968 513950 61024 514006
rect 61092 513950 61148 514006
rect 61216 513950 61272 514006
rect 61340 513950 61396 514006
rect 61464 513950 61520 514006
rect 61588 513950 61644 514006
rect 61712 513950 61768 514006
rect 61836 513950 61892 514006
rect 61960 513950 62016 514006
rect 62084 513950 62140 514006
rect 62208 513950 62264 514006
rect 62332 513950 62388 514006
rect 62456 513950 62512 514006
rect 62580 513950 62636 514006
rect 62704 513950 62760 514006
rect 62828 513950 62884 514006
rect 62952 513950 63008 514006
rect 63076 513950 63132 514006
rect 63200 513950 63256 514006
rect 63324 513950 63380 514006
rect 63448 513950 63504 514006
rect 63572 513950 63628 514006
rect 63696 513950 63752 514006
rect 63820 513950 63876 514006
rect 63944 513950 64000 514006
rect 64068 513950 64124 514006
rect 64192 513950 64248 514006
rect 64316 513950 64372 514006
rect 64440 513950 64496 514006
rect 64564 513950 64620 514006
rect 64688 513950 64744 514006
rect 64812 513950 64868 514006
rect 64936 513950 64992 514006
rect 65060 513950 65116 514006
rect 65184 513950 65240 514006
rect 65308 513950 65364 514006
rect 65432 513950 65488 514006
rect 65556 513950 65612 514006
rect 65680 513950 65736 514006
rect 65804 513950 65860 514006
rect 65928 513950 65984 514006
rect 66052 513950 66108 514006
rect 66176 513950 66232 514006
rect 66300 513950 66356 514006
rect 87884 508332 87940 508388
rect 88008 508332 88064 508388
rect 88132 508332 88188 508388
rect 88256 508332 88312 508388
rect 88380 508332 88436 508388
rect 88504 508332 88560 508388
rect 88628 508332 88684 508388
rect 88752 508332 88808 508388
rect 88876 508332 88932 508388
rect 89000 508332 89056 508388
rect 89124 508332 89180 508388
rect 89248 508332 89304 508388
rect 89372 508332 89428 508388
rect 89496 508332 89552 508388
rect 89620 508332 89676 508388
rect 89744 508332 89800 508388
rect 89868 508332 89924 508388
rect 89992 508332 90048 508388
rect 90116 508332 90172 508388
rect 90240 508332 90296 508388
rect 90364 508332 90420 508388
rect 90488 508332 90544 508388
rect 90612 508332 90668 508388
rect 90736 508332 90792 508388
rect 90860 508332 90916 508388
rect 90984 508332 91040 508388
rect 91108 508332 91164 508388
rect 91232 508332 91288 508388
rect 91356 508332 91412 508388
rect 91480 508332 91536 508388
rect 91604 508332 91660 508388
rect 91728 508332 91784 508388
rect 91852 508332 91908 508388
rect 91976 508332 92032 508388
rect 92100 508332 92156 508388
rect 92224 508332 92280 508388
rect 92348 508332 92404 508388
rect 92472 508332 92528 508388
rect 92596 508332 92652 508388
rect 92720 508332 92776 508388
rect 92844 508332 92900 508388
rect 92968 508332 93024 508388
rect 93092 508332 93148 508388
rect 93216 508332 93272 508388
rect 93340 508332 93396 508388
rect 93464 508332 93520 508388
rect 93588 508332 93644 508388
rect 93712 508332 93768 508388
rect 93836 508332 93892 508388
rect 93960 508332 94016 508388
rect 94084 508332 94140 508388
rect 94208 508332 94264 508388
rect 94332 508332 94388 508388
rect 94456 508332 94512 508388
rect 94580 508332 94636 508388
rect 94704 508332 94760 508388
rect 94828 508332 94884 508388
rect 94952 508332 95008 508388
rect 95076 508332 95132 508388
rect 95200 508332 95256 508388
rect 95324 508332 95380 508388
rect 95448 508332 95504 508388
rect 95572 508332 95628 508388
rect 95696 508332 95752 508388
rect 95820 508332 95876 508388
rect 95944 508332 96000 508388
rect 96068 508332 96124 508388
rect 96192 508332 96248 508388
rect 96316 508332 96372 508388
rect 96440 508332 96496 508388
rect 96564 508332 96620 508388
rect 96688 508332 96744 508388
rect 96812 508332 96868 508388
rect 96936 508332 96992 508388
rect 97060 508332 97116 508388
rect 97184 508332 97240 508388
rect 97308 508332 97364 508388
rect 97432 508332 97488 508388
rect 97556 508332 97612 508388
rect 97680 508332 97736 508388
rect 97804 508332 97860 508388
rect 97928 508332 97984 508388
rect 98052 508332 98108 508388
rect 98176 508332 98232 508388
rect 98300 508332 98356 508388
rect 159114 508294 159170 508350
rect 159238 508294 159294 508350
rect 159362 508294 159418 508350
rect 159486 508294 159542 508350
rect 159114 508170 159170 508226
rect 159238 508170 159294 508226
rect 159362 508170 159418 508226
rect 159486 508170 159542 508226
rect 87724 508012 87780 508068
rect 87848 508012 87904 508068
rect 87972 508012 88028 508068
rect 88096 508012 88152 508068
rect 88220 508012 88276 508068
rect 88344 508012 88400 508068
rect 88468 508012 88524 508068
rect 88592 508012 88648 508068
rect 88716 508012 88772 508068
rect 88840 508012 88896 508068
rect 88964 508012 89020 508068
rect 89088 508012 89144 508068
rect 89212 508012 89268 508068
rect 89336 508012 89392 508068
rect 89460 508012 89516 508068
rect 89584 508012 89640 508068
rect 89708 508012 89764 508068
rect 89832 508012 89888 508068
rect 89956 508012 90012 508068
rect 90080 508012 90136 508068
rect 90204 508012 90260 508068
rect 90328 508012 90384 508068
rect 90452 508012 90508 508068
rect 90576 508012 90632 508068
rect 90700 508012 90756 508068
rect 90824 508012 90880 508068
rect 90948 508012 91004 508068
rect 91072 508012 91128 508068
rect 91196 508012 91252 508068
rect 91320 508012 91376 508068
rect 91444 508012 91500 508068
rect 91568 508012 91624 508068
rect 91692 508012 91748 508068
rect 91816 508012 91872 508068
rect 91940 508012 91996 508068
rect 92064 508012 92120 508068
rect 92188 508012 92244 508068
rect 92312 508012 92368 508068
rect 92436 508012 92492 508068
rect 92560 508012 92616 508068
rect 92684 508012 92740 508068
rect 92808 508012 92864 508068
rect 92932 508012 92988 508068
rect 93056 508012 93112 508068
rect 93180 508012 93236 508068
rect 93304 508012 93360 508068
rect 93428 508012 93484 508068
rect 93552 508012 93608 508068
rect 93676 508012 93732 508068
rect 93800 508012 93856 508068
rect 93924 508012 93980 508068
rect 94048 508012 94104 508068
rect 94172 508012 94228 508068
rect 94296 508012 94352 508068
rect 94420 508012 94476 508068
rect 94544 508012 94600 508068
rect 94668 508012 94724 508068
rect 94792 508012 94848 508068
rect 94916 508012 94972 508068
rect 95040 508012 95096 508068
rect 95164 508012 95220 508068
rect 95288 508012 95344 508068
rect 95412 508012 95468 508068
rect 95536 508012 95592 508068
rect 95660 508012 95716 508068
rect 95784 508012 95840 508068
rect 95908 508012 95964 508068
rect 96032 508012 96088 508068
rect 96156 508012 96212 508068
rect 96280 508012 96336 508068
rect 96404 508012 96460 508068
rect 96528 508012 96584 508068
rect 96652 508012 96708 508068
rect 96776 508012 96832 508068
rect 96900 508012 96956 508068
rect 97024 508012 97080 508068
rect 97148 508012 97204 508068
rect 97272 508012 97328 508068
rect 97396 508012 97452 508068
rect 97520 508012 97576 508068
rect 97644 508012 97700 508068
rect 97768 508012 97824 508068
rect 97892 508012 97948 508068
rect 98016 508012 98072 508068
rect 98140 508012 98196 508068
rect 159114 508046 159170 508102
rect 159238 508046 159294 508102
rect 159362 508046 159418 508102
rect 159486 508046 159542 508102
rect 159114 507922 159170 507978
rect 159238 507922 159294 507978
rect 159362 507922 159418 507978
rect 159486 507922 159542 507978
rect 39954 496294 40010 496350
rect 40078 496294 40134 496350
rect 40202 496294 40258 496350
rect 40326 496294 40382 496350
rect 61956 496332 62012 496388
rect 62080 496332 62136 496388
rect 62204 496332 62260 496388
rect 62328 496332 62384 496388
rect 62452 496332 62508 496388
rect 62576 496332 62632 496388
rect 62700 496332 62756 496388
rect 62824 496332 62880 496388
rect 62948 496332 63004 496388
rect 63072 496332 63128 496388
rect 63196 496332 63252 496388
rect 63320 496332 63376 496388
rect 63444 496332 63500 496388
rect 63568 496332 63624 496388
rect 63692 496332 63748 496388
rect 63816 496332 63872 496388
rect 63940 496332 63996 496388
rect 64064 496332 64120 496388
rect 64188 496332 64244 496388
rect 64312 496332 64368 496388
rect 64436 496332 64492 496388
rect 64560 496332 64616 496388
rect 64684 496332 64740 496388
rect 64808 496332 64864 496388
rect 64932 496332 64988 496388
rect 65056 496332 65112 496388
rect 65180 496332 65236 496388
rect 65304 496332 65360 496388
rect 65428 496332 65484 496388
rect 65552 496332 65608 496388
rect 65676 496332 65732 496388
rect 65800 496332 65856 496388
rect 65924 496332 65980 496388
rect 66048 496332 66104 496388
rect 66172 496332 66228 496388
rect 66296 496332 66352 496388
rect 66420 496332 66476 496388
rect 66544 496332 66600 496388
rect 66668 496332 66724 496388
rect 66792 496332 66848 496388
rect 66916 496332 66972 496388
rect 67040 496332 67096 496388
rect 67164 496332 67220 496388
rect 67288 496332 67344 496388
rect 67412 496332 67468 496388
rect 67536 496332 67592 496388
rect 67660 496332 67716 496388
rect 67784 496332 67840 496388
rect 67908 496332 67964 496388
rect 39954 496170 40010 496226
rect 40078 496170 40134 496226
rect 40202 496170 40258 496226
rect 40326 496170 40382 496226
rect 39954 496046 40010 496102
rect 40078 496046 40134 496102
rect 40202 496046 40258 496102
rect 40326 496046 40382 496102
rect 39954 495922 40010 495978
rect 40078 495922 40134 495978
rect 40202 495922 40258 495978
rect 40326 495922 40382 495978
rect 62116 496007 62172 496063
rect 62240 496007 62296 496063
rect 62364 496007 62420 496063
rect 62488 496007 62544 496063
rect 62612 496007 62668 496063
rect 62736 496007 62792 496063
rect 62860 496007 62916 496063
rect 62984 496007 63040 496063
rect 63108 496007 63164 496063
rect 63232 496007 63288 496063
rect 63356 496007 63412 496063
rect 63480 496007 63536 496063
rect 63604 496007 63660 496063
rect 63728 496007 63784 496063
rect 63852 496007 63908 496063
rect 63976 496007 64032 496063
rect 64100 496007 64156 496063
rect 64224 496007 64280 496063
rect 64348 496007 64404 496063
rect 64472 496007 64528 496063
rect 64596 496007 64652 496063
rect 64720 496007 64776 496063
rect 64844 496007 64900 496063
rect 64968 496007 65024 496063
rect 65092 496007 65148 496063
rect 65216 496007 65272 496063
rect 65340 496007 65396 496063
rect 65464 496007 65520 496063
rect 65588 496007 65644 496063
rect 65712 496007 65768 496063
rect 65836 496007 65892 496063
rect 65960 496007 66016 496063
rect 66084 496007 66140 496063
rect 66208 496007 66264 496063
rect 66332 496007 66388 496063
rect 66456 496007 66512 496063
rect 66580 496007 66636 496063
rect 66704 496007 66760 496063
rect 66828 496007 66884 496063
rect 66952 496007 67008 496063
rect 67076 496007 67132 496063
rect 67200 496007 67256 496063
rect 67324 496007 67380 496063
rect 67448 496007 67504 496063
rect 67572 496007 67628 496063
rect 67696 496007 67752 496063
rect 67820 496007 67876 496063
rect 67944 496007 68000 496063
rect 68068 496007 68124 496063
rect 62116 495883 62172 495939
rect 62240 495883 62296 495939
rect 62364 495883 62420 495939
rect 62488 495883 62544 495939
rect 62612 495883 62668 495939
rect 62736 495883 62792 495939
rect 62860 495883 62916 495939
rect 62984 495883 63040 495939
rect 63108 495883 63164 495939
rect 63232 495883 63288 495939
rect 63356 495883 63412 495939
rect 63480 495883 63536 495939
rect 63604 495883 63660 495939
rect 63728 495883 63784 495939
rect 63852 495883 63908 495939
rect 63976 495883 64032 495939
rect 64100 495883 64156 495939
rect 64224 495883 64280 495939
rect 64348 495883 64404 495939
rect 64472 495883 64528 495939
rect 64596 495883 64652 495939
rect 64720 495883 64776 495939
rect 64844 495883 64900 495939
rect 64968 495883 65024 495939
rect 65092 495883 65148 495939
rect 65216 495883 65272 495939
rect 65340 495883 65396 495939
rect 65464 495883 65520 495939
rect 65588 495883 65644 495939
rect 65712 495883 65768 495939
rect 65836 495883 65892 495939
rect 65960 495883 66016 495939
rect 66084 495883 66140 495939
rect 66208 495883 66264 495939
rect 66332 495883 66388 495939
rect 66456 495883 66512 495939
rect 66580 495883 66636 495939
rect 66704 495883 66760 495939
rect 66828 495883 66884 495939
rect 66952 495883 67008 495939
rect 67076 495883 67132 495939
rect 67200 495883 67256 495939
rect 67324 495883 67380 495939
rect 67448 495883 67504 495939
rect 67572 495883 67628 495939
rect 67696 495883 67752 495939
rect 67820 495883 67876 495939
rect 67944 495883 68000 495939
rect 68068 495883 68124 495939
rect 82894 490357 82950 490413
rect 83018 490357 83074 490413
rect 82894 490233 82950 490289
rect 83018 490233 83074 490289
rect 83142 490357 83198 490413
rect 83266 490357 83322 490413
rect 83390 490357 83446 490413
rect 83514 490357 83570 490413
rect 83142 490233 83198 490289
rect 83266 490233 83322 490289
rect 83390 490233 83446 490289
rect 83514 490233 83570 490289
rect 83638 490357 83694 490413
rect 83762 490357 83818 490413
rect 83886 490357 83942 490413
rect 84010 490357 84066 490413
rect 83638 490233 83694 490289
rect 83762 490233 83818 490289
rect 83886 490233 83942 490289
rect 84010 490233 84066 490289
rect 84134 490357 84190 490413
rect 84258 490357 84314 490413
rect 84382 490357 84438 490413
rect 84506 490357 84562 490413
rect 84134 490233 84190 490289
rect 84258 490233 84314 490289
rect 84382 490233 84438 490289
rect 84506 490233 84562 490289
rect 84630 490357 84686 490413
rect 84754 490357 84810 490413
rect 84878 490357 84934 490413
rect 85002 490357 85058 490413
rect 84630 490233 84686 490289
rect 84754 490233 84810 490289
rect 84878 490233 84934 490289
rect 85002 490233 85058 490289
rect 85126 490357 85182 490413
rect 85250 490357 85306 490413
rect 85374 490357 85430 490413
rect 85498 490357 85554 490413
rect 85126 490233 85182 490289
rect 85250 490233 85306 490289
rect 85374 490233 85430 490289
rect 85498 490233 85554 490289
rect 85622 490357 85678 490413
rect 85746 490357 85802 490413
rect 85870 490357 85926 490413
rect 85994 490357 86050 490413
rect 85622 490233 85678 490289
rect 85746 490233 85802 490289
rect 85870 490233 85926 490289
rect 85994 490233 86050 490289
rect 86118 490357 86174 490413
rect 86242 490357 86298 490413
rect 86366 490357 86422 490413
rect 86490 490357 86546 490413
rect 86118 490233 86174 490289
rect 86242 490233 86298 490289
rect 86366 490233 86422 490289
rect 86490 490233 86546 490289
rect 128394 490294 128450 490350
rect 128518 490294 128574 490350
rect 128642 490294 128698 490350
rect 128766 490294 128822 490350
rect 128394 490170 128450 490226
rect 128518 490170 128574 490226
rect 128642 490170 128698 490226
rect 128766 490170 128822 490226
rect 128394 490046 128450 490102
rect 128518 490046 128574 490102
rect 128642 490046 128698 490102
rect 128766 490046 128822 490102
rect 82734 489932 82790 489988
rect 82858 489932 82914 489988
rect 82982 489932 83038 489988
rect 83106 489932 83162 489988
rect 83230 489932 83286 489988
rect 83354 489932 83410 489988
rect 83478 489932 83534 489988
rect 83602 489932 83658 489988
rect 83726 489932 83782 489988
rect 83850 489932 83906 489988
rect 83974 489932 84030 489988
rect 84098 489932 84154 489988
rect 84222 489932 84278 489988
rect 84346 489932 84402 489988
rect 84470 489932 84526 489988
rect 84594 489932 84650 489988
rect 84718 489932 84774 489988
rect 84842 489932 84898 489988
rect 84966 489932 85022 489988
rect 85090 489932 85146 489988
rect 85214 489932 85270 489988
rect 85338 489932 85394 489988
rect 85462 489932 85518 489988
rect 85586 489932 85642 489988
rect 85710 489932 85766 489988
rect 85834 489932 85890 489988
rect 85958 489932 86014 489988
rect 86082 489932 86138 489988
rect 86206 489932 86262 489988
rect 86330 489932 86386 489988
rect 128394 489922 128450 489978
rect 128518 489922 128574 489978
rect 128642 489922 128698 489978
rect 128766 489922 128822 489978
rect 39954 478294 40010 478350
rect 40078 478294 40134 478350
rect 40202 478294 40258 478350
rect 40326 478294 40382 478350
rect 39954 478170 40010 478226
rect 40078 478170 40134 478226
rect 40202 478170 40258 478226
rect 40326 478170 40382 478226
rect 39954 478046 40010 478102
rect 40078 478046 40134 478102
rect 40202 478046 40258 478102
rect 40326 478046 40382 478102
rect 39954 477922 40010 477978
rect 40078 477922 40134 477978
rect 40202 477922 40258 477978
rect 40326 477922 40382 477978
rect 39954 460294 40010 460350
rect 40078 460294 40134 460350
rect 40202 460294 40258 460350
rect 40326 460294 40382 460350
rect 39954 460170 40010 460226
rect 40078 460170 40134 460226
rect 40202 460170 40258 460226
rect 40326 460170 40382 460226
rect 39954 460046 40010 460102
rect 40078 460046 40134 460102
rect 40202 460046 40258 460102
rect 40326 460046 40382 460102
rect 39954 459922 40010 459978
rect 40078 459922 40134 459978
rect 40202 459922 40258 459978
rect 40326 459922 40382 459978
rect 39954 442294 40010 442350
rect 40078 442294 40134 442350
rect 40202 442294 40258 442350
rect 40326 442294 40382 442350
rect 39954 442170 40010 442226
rect 40078 442170 40134 442226
rect 40202 442170 40258 442226
rect 40326 442170 40382 442226
rect 39954 442046 40010 442102
rect 40078 442046 40134 442102
rect 40202 442046 40258 442102
rect 40326 442046 40382 442102
rect 39954 441922 40010 441978
rect 40078 441922 40134 441978
rect 40202 441922 40258 441978
rect 40326 441922 40382 441978
rect 39954 424294 40010 424350
rect 40078 424294 40134 424350
rect 40202 424294 40258 424350
rect 40326 424294 40382 424350
rect 39954 424170 40010 424226
rect 40078 424170 40134 424226
rect 40202 424170 40258 424226
rect 40326 424170 40382 424226
rect 39954 424046 40010 424102
rect 40078 424046 40134 424102
rect 40202 424046 40258 424102
rect 40326 424046 40382 424102
rect 39954 423922 40010 423978
rect 40078 423922 40134 423978
rect 40202 423922 40258 423978
rect 40326 423922 40382 423978
rect 39954 406294 40010 406350
rect 40078 406294 40134 406350
rect 40202 406294 40258 406350
rect 40326 406294 40382 406350
rect 39954 406170 40010 406226
rect 40078 406170 40134 406226
rect 40202 406170 40258 406226
rect 40326 406170 40382 406226
rect 39954 406046 40010 406102
rect 40078 406046 40134 406102
rect 40202 406046 40258 406102
rect 40326 406046 40382 406102
rect 39954 405922 40010 405978
rect 40078 405922 40134 405978
rect 40202 405922 40258 405978
rect 40326 405922 40382 405978
rect 39954 388294 40010 388350
rect 40078 388294 40134 388350
rect 40202 388294 40258 388350
rect 40326 388294 40382 388350
rect 39954 388170 40010 388226
rect 40078 388170 40134 388226
rect 40202 388170 40258 388226
rect 40326 388170 40382 388226
rect 39954 388046 40010 388102
rect 40078 388046 40134 388102
rect 40202 388046 40258 388102
rect 40326 388046 40382 388102
rect 39954 387922 40010 387978
rect 40078 387922 40134 387978
rect 40202 387922 40258 387978
rect 40326 387922 40382 387978
rect 39954 370294 40010 370350
rect 40078 370294 40134 370350
rect 40202 370294 40258 370350
rect 40326 370294 40382 370350
rect 39954 370170 40010 370226
rect 40078 370170 40134 370226
rect 40202 370170 40258 370226
rect 40326 370170 40382 370226
rect 39954 370046 40010 370102
rect 40078 370046 40134 370102
rect 40202 370046 40258 370102
rect 40326 370046 40382 370102
rect 39954 369922 40010 369978
rect 40078 369922 40134 369978
rect 40202 369922 40258 369978
rect 40326 369922 40382 369978
rect 66954 472294 67010 472350
rect 67078 472294 67134 472350
rect 67202 472294 67258 472350
rect 67326 472294 67382 472350
rect 66954 472170 67010 472226
rect 67078 472170 67134 472226
rect 67202 472170 67258 472226
rect 67326 472170 67382 472226
rect 66954 472046 67010 472102
rect 67078 472046 67134 472102
rect 67202 472046 67258 472102
rect 67326 472046 67382 472102
rect 66954 471922 67010 471978
rect 67078 471922 67134 471978
rect 67202 471922 67258 471978
rect 67326 471922 67382 471978
rect 66954 454294 67010 454350
rect 67078 454294 67134 454350
rect 67202 454294 67258 454350
rect 67326 454294 67382 454350
rect 66954 454170 67010 454226
rect 67078 454170 67134 454226
rect 67202 454170 67258 454226
rect 67326 454170 67382 454226
rect 66954 454046 67010 454102
rect 67078 454046 67134 454102
rect 67202 454046 67258 454102
rect 67326 454046 67382 454102
rect 66954 453922 67010 453978
rect 67078 453922 67134 453978
rect 67202 453922 67258 453978
rect 67326 453922 67382 453978
rect 66954 436294 67010 436350
rect 67078 436294 67134 436350
rect 67202 436294 67258 436350
rect 67326 436294 67382 436350
rect 66954 436170 67010 436226
rect 67078 436170 67134 436226
rect 67202 436170 67258 436226
rect 67326 436170 67382 436226
rect 66954 436046 67010 436102
rect 67078 436046 67134 436102
rect 67202 436046 67258 436102
rect 67326 436046 67382 436102
rect 66954 435922 67010 435978
rect 67078 435922 67134 435978
rect 67202 435922 67258 435978
rect 67326 435922 67382 435978
rect 66954 418294 67010 418350
rect 67078 418294 67134 418350
rect 67202 418294 67258 418350
rect 67326 418294 67382 418350
rect 66954 418170 67010 418226
rect 67078 418170 67134 418226
rect 67202 418170 67258 418226
rect 67326 418170 67382 418226
rect 66954 418046 67010 418102
rect 67078 418046 67134 418102
rect 67202 418046 67258 418102
rect 67326 418046 67382 418102
rect 66954 417922 67010 417978
rect 67078 417922 67134 417978
rect 67202 417922 67258 417978
rect 67326 417922 67382 417978
rect 66954 400294 67010 400350
rect 67078 400294 67134 400350
rect 67202 400294 67258 400350
rect 67326 400294 67382 400350
rect 66954 400170 67010 400226
rect 67078 400170 67134 400226
rect 67202 400170 67258 400226
rect 67326 400170 67382 400226
rect 66954 400046 67010 400102
rect 67078 400046 67134 400102
rect 67202 400046 67258 400102
rect 67326 400046 67382 400102
rect 66954 399922 67010 399978
rect 67078 399922 67134 399978
rect 67202 399922 67258 399978
rect 67326 399922 67382 399978
rect 66954 382294 67010 382350
rect 67078 382294 67134 382350
rect 67202 382294 67258 382350
rect 67326 382294 67382 382350
rect 66954 382170 67010 382226
rect 67078 382170 67134 382226
rect 67202 382170 67258 382226
rect 67326 382170 67382 382226
rect 66954 382046 67010 382102
rect 67078 382046 67134 382102
rect 67202 382046 67258 382102
rect 67326 382046 67382 382102
rect 66954 381922 67010 381978
rect 67078 381922 67134 381978
rect 67202 381922 67258 381978
rect 67326 381922 67382 381978
rect 39954 352294 40010 352350
rect 40078 352294 40134 352350
rect 40202 352294 40258 352350
rect 40326 352294 40382 352350
rect 39954 352170 40010 352226
rect 40078 352170 40134 352226
rect 40202 352170 40258 352226
rect 40326 352170 40382 352226
rect 39954 352046 40010 352102
rect 40078 352046 40134 352102
rect 40202 352046 40258 352102
rect 40326 352046 40382 352102
rect 39954 351922 40010 351978
rect 40078 351922 40134 351978
rect 40202 351922 40258 351978
rect 40326 351922 40382 351978
rect 39954 334294 40010 334350
rect 40078 334294 40134 334350
rect 40202 334294 40258 334350
rect 40326 334294 40382 334350
rect 39954 334170 40010 334226
rect 40078 334170 40134 334226
rect 40202 334170 40258 334226
rect 40326 334170 40382 334226
rect 39954 334046 40010 334102
rect 40078 334046 40134 334102
rect 40202 334046 40258 334102
rect 40326 334046 40382 334102
rect 39954 333922 40010 333978
rect 40078 333922 40134 333978
rect 40202 333922 40258 333978
rect 40326 333922 40382 333978
rect 39954 316294 40010 316350
rect 40078 316294 40134 316350
rect 40202 316294 40258 316350
rect 40326 316294 40382 316350
rect 39954 316170 40010 316226
rect 40078 316170 40134 316226
rect 40202 316170 40258 316226
rect 40326 316170 40382 316226
rect 39954 316046 40010 316102
rect 40078 316046 40134 316102
rect 40202 316046 40258 316102
rect 40326 316046 40382 316102
rect 39954 315922 40010 315978
rect 40078 315922 40134 315978
rect 40202 315922 40258 315978
rect 40326 315922 40382 315978
rect 63756 366362 63812 366418
rect 66954 364294 67010 364350
rect 67078 364294 67134 364350
rect 67202 364294 67258 364350
rect 67326 364294 67382 364350
rect 66954 364170 67010 364226
rect 67078 364170 67134 364226
rect 67202 364170 67258 364226
rect 67326 364170 67382 364226
rect 66954 364046 67010 364102
rect 67078 364046 67134 364102
rect 67202 364046 67258 364102
rect 67326 364046 67382 364102
rect 66954 363922 67010 363978
rect 67078 363922 67134 363978
rect 67202 363922 67258 363978
rect 67326 363922 67382 363978
rect 66954 346294 67010 346350
rect 67078 346294 67134 346350
rect 67202 346294 67258 346350
rect 67326 346294 67382 346350
rect 66954 346170 67010 346226
rect 67078 346170 67134 346226
rect 67202 346170 67258 346226
rect 67326 346170 67382 346226
rect 66954 346046 67010 346102
rect 67078 346046 67134 346102
rect 67202 346046 67258 346102
rect 67326 346046 67382 346102
rect 66954 345922 67010 345978
rect 67078 345922 67134 345978
rect 67202 345922 67258 345978
rect 67326 345922 67382 345978
rect 66954 328294 67010 328350
rect 67078 328294 67134 328350
rect 67202 328294 67258 328350
rect 67326 328294 67382 328350
rect 66954 328170 67010 328226
rect 67078 328170 67134 328226
rect 67202 328170 67258 328226
rect 67326 328170 67382 328226
rect 66954 328046 67010 328102
rect 67078 328046 67134 328102
rect 67202 328046 67258 328102
rect 67326 328046 67382 328102
rect 66954 327922 67010 327978
rect 67078 327922 67134 327978
rect 67202 327922 67258 327978
rect 67326 327922 67382 327978
rect 66954 310294 67010 310350
rect 67078 310294 67134 310350
rect 67202 310294 67258 310350
rect 67326 310294 67382 310350
rect 66954 310170 67010 310226
rect 67078 310170 67134 310226
rect 67202 310170 67258 310226
rect 67326 310170 67382 310226
rect 66954 310046 67010 310102
rect 67078 310046 67134 310102
rect 67202 310046 67258 310102
rect 67326 310046 67382 310102
rect 66954 309922 67010 309978
rect 67078 309922 67134 309978
rect 67202 309922 67258 309978
rect 67326 309922 67382 309978
rect 39954 298294 40010 298350
rect 40078 298294 40134 298350
rect 40202 298294 40258 298350
rect 40326 298294 40382 298350
rect 39954 298170 40010 298226
rect 40078 298170 40134 298226
rect 40202 298170 40258 298226
rect 40326 298170 40382 298226
rect 39954 298046 40010 298102
rect 40078 298046 40134 298102
rect 40202 298046 40258 298102
rect 40326 298046 40382 298102
rect 70674 478294 70730 478350
rect 70798 478294 70854 478350
rect 70922 478294 70978 478350
rect 71046 478294 71102 478350
rect 70674 478170 70730 478226
rect 70798 478170 70854 478226
rect 70922 478170 70978 478226
rect 71046 478170 71102 478226
rect 77956 478252 78012 478308
rect 78080 478252 78136 478308
rect 78204 478252 78260 478308
rect 78328 478252 78384 478308
rect 78452 478252 78508 478308
rect 78576 478252 78632 478308
rect 78700 478252 78756 478308
rect 78824 478252 78880 478308
rect 78948 478252 79004 478308
rect 70674 478046 70730 478102
rect 70798 478046 70854 478102
rect 70922 478046 70978 478102
rect 71046 478046 71102 478102
rect 70674 477922 70730 477978
rect 70798 477922 70854 477978
rect 70922 477922 70978 477978
rect 71046 477922 71102 477978
rect 78586 477932 78642 477988
rect 78710 477932 78766 477988
rect 78834 477932 78890 477988
rect 78958 477932 79014 477988
rect 70674 460294 70730 460350
rect 70798 460294 70854 460350
rect 70922 460294 70978 460350
rect 71046 460294 71102 460350
rect 70674 460170 70730 460226
rect 70798 460170 70854 460226
rect 70922 460170 70978 460226
rect 71046 460170 71102 460226
rect 70674 460046 70730 460102
rect 70798 460046 70854 460102
rect 70922 460046 70978 460102
rect 71046 460046 71102 460102
rect 70674 459922 70730 459978
rect 70798 459922 70854 459978
rect 70922 459922 70978 459978
rect 71046 459922 71102 459978
rect 70674 442294 70730 442350
rect 70798 442294 70854 442350
rect 70922 442294 70978 442350
rect 71046 442294 71102 442350
rect 70674 442170 70730 442226
rect 70798 442170 70854 442226
rect 70922 442170 70978 442226
rect 71046 442170 71102 442226
rect 70674 442046 70730 442102
rect 70798 442046 70854 442102
rect 70922 442046 70978 442102
rect 71046 442046 71102 442102
rect 70674 441922 70730 441978
rect 70798 441922 70854 441978
rect 70922 441922 70978 441978
rect 71046 441922 71102 441978
rect 70674 424294 70730 424350
rect 70798 424294 70854 424350
rect 70922 424294 70978 424350
rect 71046 424294 71102 424350
rect 70674 424170 70730 424226
rect 70798 424170 70854 424226
rect 70922 424170 70978 424226
rect 71046 424170 71102 424226
rect 70674 424046 70730 424102
rect 70798 424046 70854 424102
rect 70922 424046 70978 424102
rect 71046 424046 71102 424102
rect 70674 423922 70730 423978
rect 70798 423922 70854 423978
rect 70922 423922 70978 423978
rect 71046 423922 71102 423978
rect 70674 406294 70730 406350
rect 70798 406294 70854 406350
rect 70922 406294 70978 406350
rect 71046 406294 71102 406350
rect 70674 406170 70730 406226
rect 70798 406170 70854 406226
rect 70922 406170 70978 406226
rect 71046 406170 71102 406226
rect 70674 406046 70730 406102
rect 70798 406046 70854 406102
rect 70922 406046 70978 406102
rect 71046 406046 71102 406102
rect 70674 405922 70730 405978
rect 70798 405922 70854 405978
rect 70922 405922 70978 405978
rect 71046 405922 71102 405978
rect 70674 388294 70730 388350
rect 70798 388294 70854 388350
rect 70922 388294 70978 388350
rect 71046 388294 71102 388350
rect 70674 388170 70730 388226
rect 70798 388170 70854 388226
rect 70922 388170 70978 388226
rect 71046 388170 71102 388226
rect 70674 388046 70730 388102
rect 70798 388046 70854 388102
rect 70922 388046 70978 388102
rect 71046 388046 71102 388102
rect 70674 387922 70730 387978
rect 70798 387922 70854 387978
rect 70922 387922 70978 387978
rect 71046 387922 71102 387978
rect 70674 370294 70730 370350
rect 70798 370294 70854 370350
rect 70922 370294 70978 370350
rect 71046 370294 71102 370350
rect 70674 370170 70730 370226
rect 70798 370170 70854 370226
rect 70922 370170 70978 370226
rect 71046 370170 71102 370226
rect 70674 370046 70730 370102
rect 70798 370046 70854 370102
rect 70922 370046 70978 370102
rect 71046 370046 71102 370102
rect 70674 369922 70730 369978
rect 70798 369922 70854 369978
rect 70922 369922 70978 369978
rect 71046 369922 71102 369978
rect 97674 472294 97730 472350
rect 97798 472294 97854 472350
rect 97922 472294 97978 472350
rect 98046 472294 98102 472350
rect 97674 472170 97730 472226
rect 97798 472170 97854 472226
rect 97922 472170 97978 472226
rect 98046 472170 98102 472226
rect 97674 472046 97730 472102
rect 97798 472046 97854 472102
rect 97922 472046 97978 472102
rect 98046 472046 98102 472102
rect 97674 471922 97730 471978
rect 97798 471922 97854 471978
rect 97922 471922 97978 471978
rect 98046 471922 98102 471978
rect 97674 454294 97730 454350
rect 97798 454294 97854 454350
rect 97922 454294 97978 454350
rect 98046 454294 98102 454350
rect 97674 454170 97730 454226
rect 97798 454170 97854 454226
rect 97922 454170 97978 454226
rect 98046 454170 98102 454226
rect 97674 454046 97730 454102
rect 97798 454046 97854 454102
rect 97922 454046 97978 454102
rect 98046 454046 98102 454102
rect 97674 453922 97730 453978
rect 97798 453922 97854 453978
rect 97922 453922 97978 453978
rect 98046 453922 98102 453978
rect 97674 436294 97730 436350
rect 97798 436294 97854 436350
rect 97922 436294 97978 436350
rect 98046 436294 98102 436350
rect 97674 436170 97730 436226
rect 97798 436170 97854 436226
rect 97922 436170 97978 436226
rect 98046 436170 98102 436226
rect 97674 436046 97730 436102
rect 97798 436046 97854 436102
rect 97922 436046 97978 436102
rect 98046 436046 98102 436102
rect 97674 435922 97730 435978
rect 97798 435922 97854 435978
rect 97922 435922 97978 435978
rect 98046 435922 98102 435978
rect 97674 418294 97730 418350
rect 97798 418294 97854 418350
rect 97922 418294 97978 418350
rect 98046 418294 98102 418350
rect 97674 418170 97730 418226
rect 97798 418170 97854 418226
rect 97922 418170 97978 418226
rect 98046 418170 98102 418226
rect 97674 418046 97730 418102
rect 97798 418046 97854 418102
rect 97922 418046 97978 418102
rect 98046 418046 98102 418102
rect 97674 417922 97730 417978
rect 97798 417922 97854 417978
rect 97922 417922 97978 417978
rect 98046 417922 98102 417978
rect 97674 400294 97730 400350
rect 97798 400294 97854 400350
rect 97922 400294 97978 400350
rect 98046 400294 98102 400350
rect 97674 400170 97730 400226
rect 97798 400170 97854 400226
rect 97922 400170 97978 400226
rect 98046 400170 98102 400226
rect 97674 400046 97730 400102
rect 97798 400046 97854 400102
rect 97922 400046 97978 400102
rect 98046 400046 98102 400102
rect 97674 399922 97730 399978
rect 97798 399922 97854 399978
rect 97922 399922 97978 399978
rect 98046 399922 98102 399978
rect 101394 460294 101450 460350
rect 101518 460294 101574 460350
rect 101642 460294 101698 460350
rect 101766 460294 101822 460350
rect 101394 460170 101450 460226
rect 101518 460170 101574 460226
rect 101642 460170 101698 460226
rect 101766 460170 101822 460226
rect 101394 460046 101450 460102
rect 101518 460046 101574 460102
rect 101642 460046 101698 460102
rect 101766 460046 101822 460102
rect 101394 459922 101450 459978
rect 101518 459922 101574 459978
rect 101642 459922 101698 459978
rect 101766 459922 101822 459978
rect 101394 442294 101450 442350
rect 101518 442294 101574 442350
rect 101642 442294 101698 442350
rect 101766 442294 101822 442350
rect 101394 442170 101450 442226
rect 101518 442170 101574 442226
rect 101642 442170 101698 442226
rect 101766 442170 101822 442226
rect 101394 442046 101450 442102
rect 101518 442046 101574 442102
rect 101642 442046 101698 442102
rect 101766 442046 101822 442102
rect 101394 441922 101450 441978
rect 101518 441922 101574 441978
rect 101642 441922 101698 441978
rect 101766 441922 101822 441978
rect 101394 424294 101450 424350
rect 101518 424294 101574 424350
rect 101642 424294 101698 424350
rect 101766 424294 101822 424350
rect 101394 424170 101450 424226
rect 101518 424170 101574 424226
rect 101642 424170 101698 424226
rect 101766 424170 101822 424226
rect 101394 424046 101450 424102
rect 101518 424046 101574 424102
rect 101642 424046 101698 424102
rect 101766 424046 101822 424102
rect 101394 423922 101450 423978
rect 101518 423922 101574 423978
rect 101642 423922 101698 423978
rect 101766 423922 101822 423978
rect 101394 406294 101450 406350
rect 101518 406294 101574 406350
rect 101642 406294 101698 406350
rect 101766 406294 101822 406350
rect 101394 406170 101450 406226
rect 101518 406170 101574 406226
rect 101642 406170 101698 406226
rect 101766 406170 101822 406226
rect 101394 406046 101450 406102
rect 101518 406046 101574 406102
rect 101642 406046 101698 406102
rect 101766 406046 101822 406102
rect 101394 405922 101450 405978
rect 101518 405922 101574 405978
rect 101642 405922 101698 405978
rect 101766 405922 101822 405978
rect 101394 388294 101450 388350
rect 101518 388294 101574 388350
rect 101642 388294 101698 388350
rect 101766 388294 101822 388350
rect 101394 388170 101450 388226
rect 101518 388170 101574 388226
rect 101642 388170 101698 388226
rect 101766 388170 101822 388226
rect 101394 388046 101450 388102
rect 101518 388046 101574 388102
rect 101642 388046 101698 388102
rect 101766 388046 101822 388102
rect 101394 387922 101450 387978
rect 101518 387922 101574 387978
rect 101642 387922 101698 387978
rect 101766 387922 101822 387978
rect 97674 382294 97730 382350
rect 97798 382294 97854 382350
rect 97922 382294 97978 382350
rect 98046 382294 98102 382350
rect 97674 382170 97730 382226
rect 97798 382170 97854 382226
rect 97922 382170 97978 382226
rect 98046 382170 98102 382226
rect 97674 382046 97730 382102
rect 97798 382046 97854 382102
rect 97922 382046 97978 382102
rect 98046 382046 98102 382102
rect 97674 381922 97730 381978
rect 97798 381922 97854 381978
rect 97922 381922 97978 381978
rect 98046 381922 98102 381978
rect 93996 367082 94052 367138
rect 70674 352294 70730 352350
rect 70798 352294 70854 352350
rect 70922 352294 70978 352350
rect 71046 352294 71102 352350
rect 70674 352170 70730 352226
rect 70798 352170 70854 352226
rect 70922 352170 70978 352226
rect 71046 352170 71102 352226
rect 70674 352046 70730 352102
rect 70798 352046 70854 352102
rect 70922 352046 70978 352102
rect 71046 352046 71102 352102
rect 70674 351922 70730 351978
rect 70798 351922 70854 351978
rect 70922 351922 70978 351978
rect 71046 351922 71102 351978
rect 70674 334294 70730 334350
rect 70798 334294 70854 334350
rect 70922 334294 70978 334350
rect 71046 334294 71102 334350
rect 70674 334170 70730 334226
rect 70798 334170 70854 334226
rect 70922 334170 70978 334226
rect 71046 334170 71102 334226
rect 70674 334046 70730 334102
rect 70798 334046 70854 334102
rect 70922 334046 70978 334102
rect 71046 334046 71102 334102
rect 70674 333922 70730 333978
rect 70798 333922 70854 333978
rect 70922 333922 70978 333978
rect 71046 333922 71102 333978
rect 70674 316294 70730 316350
rect 70798 316294 70854 316350
rect 70922 316294 70978 316350
rect 71046 316294 71102 316350
rect 70674 316170 70730 316226
rect 70798 316170 70854 316226
rect 70922 316170 70978 316226
rect 71046 316170 71102 316226
rect 70674 316046 70730 316102
rect 70798 316046 70854 316102
rect 70922 316046 70978 316102
rect 71046 316046 71102 316102
rect 70674 315922 70730 315978
rect 70798 315922 70854 315978
rect 70922 315922 70978 315978
rect 71046 315922 71102 315978
rect 78876 365822 78932 365878
rect 97674 364294 97730 364350
rect 97798 364294 97854 364350
rect 97922 364294 97978 364350
rect 98046 364294 98102 364350
rect 97674 364170 97730 364226
rect 97798 364170 97854 364226
rect 97922 364170 97978 364226
rect 98046 364170 98102 364226
rect 97674 364046 97730 364102
rect 97798 364046 97854 364102
rect 97922 364046 97978 364102
rect 98046 364046 98102 364102
rect 97674 363922 97730 363978
rect 97798 363922 97854 363978
rect 97922 363922 97978 363978
rect 98046 363922 98102 363978
rect 97674 346294 97730 346350
rect 97798 346294 97854 346350
rect 97922 346294 97978 346350
rect 98046 346294 98102 346350
rect 97674 346170 97730 346226
rect 97798 346170 97854 346226
rect 97922 346170 97978 346226
rect 98046 346170 98102 346226
rect 97674 346046 97730 346102
rect 97798 346046 97854 346102
rect 97922 346046 97978 346102
rect 98046 346046 98102 346102
rect 97674 345922 97730 345978
rect 97798 345922 97854 345978
rect 97922 345922 97978 345978
rect 98046 345922 98102 345978
rect 97674 328294 97730 328350
rect 97798 328294 97854 328350
rect 97922 328294 97978 328350
rect 98046 328294 98102 328350
rect 97674 328170 97730 328226
rect 97798 328170 97854 328226
rect 97922 328170 97978 328226
rect 98046 328170 98102 328226
rect 97674 328046 97730 328102
rect 97798 328046 97854 328102
rect 97922 328046 97978 328102
rect 98046 328046 98102 328102
rect 97674 327922 97730 327978
rect 97798 327922 97854 327978
rect 97922 327922 97978 327978
rect 98046 327922 98102 327978
rect 97674 310294 97730 310350
rect 97798 310294 97854 310350
rect 97922 310294 97978 310350
rect 98046 310294 98102 310350
rect 97674 310170 97730 310226
rect 97798 310170 97854 310226
rect 97922 310170 97978 310226
rect 98046 310170 98102 310226
rect 97674 310046 97730 310102
rect 97798 310046 97854 310102
rect 97922 310046 97978 310102
rect 98046 310046 98102 310102
rect 97674 309922 97730 309978
rect 97798 309922 97854 309978
rect 97922 309922 97978 309978
rect 98046 309922 98102 309978
rect 70674 298366 70730 298422
rect 70798 298366 70854 298422
rect 70922 298366 70978 298422
rect 71046 298366 71102 298422
rect 70674 298242 70730 298298
rect 70798 298242 70854 298298
rect 70922 298242 70978 298298
rect 71046 298242 71102 298298
rect 70674 298118 70730 298174
rect 70798 298118 70854 298174
rect 70922 298118 70978 298174
rect 71046 298118 71102 298174
rect 39954 297922 40010 297978
rect 40078 297922 40134 297978
rect 40202 297922 40258 297978
rect 40326 297922 40382 297978
rect 44518 292294 44574 292350
rect 44642 292294 44698 292350
rect 44518 292170 44574 292226
rect 44642 292170 44698 292226
rect 44518 292046 44574 292102
rect 44642 292046 44698 292102
rect 44518 291922 44574 291978
rect 44642 291922 44698 291978
rect 75238 292294 75294 292350
rect 75362 292294 75418 292350
rect 75238 292170 75294 292226
rect 75362 292170 75418 292226
rect 75238 292046 75294 292102
rect 75362 292046 75418 292102
rect 75238 291922 75294 291978
rect 75362 291922 75418 291978
rect 97674 292294 97730 292350
rect 97798 292294 97854 292350
rect 97922 292294 97978 292350
rect 98046 292294 98102 292350
rect 97674 292170 97730 292226
rect 97798 292170 97854 292226
rect 97922 292170 97978 292226
rect 98046 292170 98102 292226
rect 97674 292046 97730 292102
rect 97798 292046 97854 292102
rect 97922 292046 97978 292102
rect 98046 292046 98102 292102
rect 97674 291922 97730 291978
rect 97798 291922 97854 291978
rect 97922 291922 97978 291978
rect 98046 291922 98102 291978
rect 39954 280294 40010 280350
rect 40078 280294 40134 280350
rect 40202 280294 40258 280350
rect 40326 280294 40382 280350
rect 39954 280170 40010 280226
rect 40078 280170 40134 280226
rect 40202 280170 40258 280226
rect 40326 280170 40382 280226
rect 39954 280046 40010 280102
rect 40078 280046 40134 280102
rect 40202 280046 40258 280102
rect 40326 280046 40382 280102
rect 39954 279922 40010 279978
rect 40078 279922 40134 279978
rect 40202 279922 40258 279978
rect 40326 279922 40382 279978
rect 59878 280294 59934 280350
rect 60002 280294 60058 280350
rect 59878 280170 59934 280226
rect 60002 280170 60058 280226
rect 59878 280046 59934 280102
rect 60002 280046 60058 280102
rect 59878 279922 59934 279978
rect 60002 279922 60058 279978
rect 90598 280294 90654 280350
rect 90722 280294 90778 280350
rect 90598 280170 90654 280226
rect 90722 280170 90778 280226
rect 90598 280046 90654 280102
rect 90722 280046 90778 280102
rect 90598 279922 90654 279978
rect 90722 279922 90778 279978
rect 44518 274294 44574 274350
rect 44642 274294 44698 274350
rect 44518 274170 44574 274226
rect 44642 274170 44698 274226
rect 44518 274046 44574 274102
rect 44642 274046 44698 274102
rect 44518 273922 44574 273978
rect 44642 273922 44698 273978
rect 75238 274294 75294 274350
rect 75362 274294 75418 274350
rect 75238 274170 75294 274226
rect 75362 274170 75418 274226
rect 75238 274046 75294 274102
rect 75362 274046 75418 274102
rect 75238 273922 75294 273978
rect 75362 273922 75418 273978
rect 97674 274294 97730 274350
rect 97798 274294 97854 274350
rect 97922 274294 97978 274350
rect 98046 274294 98102 274350
rect 97674 274170 97730 274226
rect 97798 274170 97854 274226
rect 97922 274170 97978 274226
rect 98046 274170 98102 274226
rect 97674 274046 97730 274102
rect 97798 274046 97854 274102
rect 97922 274046 97978 274102
rect 98046 274046 98102 274102
rect 97674 273922 97730 273978
rect 97798 273922 97854 273978
rect 97922 273922 97978 273978
rect 98046 273922 98102 273978
rect 39954 262294 40010 262350
rect 40078 262294 40134 262350
rect 40202 262294 40258 262350
rect 40326 262294 40382 262350
rect 39954 262170 40010 262226
rect 40078 262170 40134 262226
rect 40202 262170 40258 262226
rect 40326 262170 40382 262226
rect 39954 262046 40010 262102
rect 40078 262046 40134 262102
rect 40202 262046 40258 262102
rect 40326 262046 40382 262102
rect 39954 261922 40010 261978
rect 40078 261922 40134 261978
rect 40202 261922 40258 261978
rect 40326 261922 40382 261978
rect 59878 262294 59934 262350
rect 60002 262294 60058 262350
rect 59878 262170 59934 262226
rect 60002 262170 60058 262226
rect 59878 262046 59934 262102
rect 60002 262046 60058 262102
rect 59878 261922 59934 261978
rect 60002 261922 60058 261978
rect 90598 262294 90654 262350
rect 90722 262294 90778 262350
rect 90598 262170 90654 262226
rect 90722 262170 90778 262226
rect 90598 262046 90654 262102
rect 90722 262046 90778 262102
rect 90598 261922 90654 261978
rect 90722 261922 90778 261978
rect 44518 256294 44574 256350
rect 44642 256294 44698 256350
rect 44518 256170 44574 256226
rect 44642 256170 44698 256226
rect 44518 256046 44574 256102
rect 44642 256046 44698 256102
rect 44518 255922 44574 255978
rect 44642 255922 44698 255978
rect 75238 256294 75294 256350
rect 75362 256294 75418 256350
rect 75238 256170 75294 256226
rect 75362 256170 75418 256226
rect 75238 256046 75294 256102
rect 75362 256046 75418 256102
rect 75238 255922 75294 255978
rect 75362 255922 75418 255978
rect 97674 256294 97730 256350
rect 97798 256294 97854 256350
rect 97922 256294 97978 256350
rect 98046 256294 98102 256350
rect 97674 256170 97730 256226
rect 97798 256170 97854 256226
rect 97922 256170 97978 256226
rect 98046 256170 98102 256226
rect 97674 256046 97730 256102
rect 97798 256046 97854 256102
rect 97922 256046 97978 256102
rect 98046 256046 98102 256102
rect 97674 255922 97730 255978
rect 97798 255922 97854 255978
rect 97922 255922 97978 255978
rect 98046 255922 98102 255978
rect 39954 244294 40010 244350
rect 40078 244294 40134 244350
rect 40202 244294 40258 244350
rect 40326 244294 40382 244350
rect 39954 244170 40010 244226
rect 40078 244170 40134 244226
rect 40202 244170 40258 244226
rect 40326 244170 40382 244226
rect 39954 244046 40010 244102
rect 40078 244046 40134 244102
rect 40202 244046 40258 244102
rect 40326 244046 40382 244102
rect 39954 243922 40010 243978
rect 40078 243922 40134 243978
rect 40202 243922 40258 243978
rect 40326 243922 40382 243978
rect 46172 247022 46228 247078
rect 59878 244294 59934 244350
rect 60002 244294 60058 244350
rect 59878 244170 59934 244226
rect 60002 244170 60058 244226
rect 59878 244046 59934 244102
rect 60002 244046 60058 244102
rect 59878 243922 59934 243978
rect 60002 243922 60058 243978
rect 39954 226294 40010 226350
rect 40078 226294 40134 226350
rect 40202 226294 40258 226350
rect 40326 226294 40382 226350
rect 39954 226170 40010 226226
rect 40078 226170 40134 226226
rect 40202 226170 40258 226226
rect 40326 226170 40382 226226
rect 39954 226046 40010 226102
rect 40078 226046 40134 226102
rect 40202 226046 40258 226102
rect 40326 226046 40382 226102
rect 39954 225922 40010 225978
rect 40078 225922 40134 225978
rect 40202 225922 40258 225978
rect 40326 225922 40382 225978
rect 36234 202294 36290 202350
rect 36358 202294 36414 202350
rect 36482 202294 36538 202350
rect 36606 202294 36662 202350
rect 36234 202170 36290 202226
rect 36358 202170 36414 202226
rect 36482 202170 36538 202226
rect 36606 202170 36662 202226
rect 36234 202046 36290 202102
rect 36358 202046 36414 202102
rect 36482 202046 36538 202102
rect 36606 202046 36662 202102
rect 36234 201922 36290 201978
rect 36358 201922 36414 201978
rect 36482 201922 36538 201978
rect 36606 201922 36662 201978
rect 36234 184294 36290 184350
rect 36358 184294 36414 184350
rect 36482 184294 36538 184350
rect 36606 184294 36662 184350
rect 36234 184170 36290 184226
rect 36358 184170 36414 184226
rect 36482 184170 36538 184226
rect 36606 184170 36662 184226
rect 36234 184046 36290 184102
rect 36358 184046 36414 184102
rect 36482 184046 36538 184102
rect 36606 184046 36662 184102
rect 36234 183922 36290 183978
rect 36358 183922 36414 183978
rect 36482 183922 36538 183978
rect 36606 183922 36662 183978
rect 36234 166294 36290 166350
rect 36358 166294 36414 166350
rect 36482 166294 36538 166350
rect 36606 166294 36662 166350
rect 36234 166170 36290 166226
rect 36358 166170 36414 166226
rect 36482 166170 36538 166226
rect 36606 166170 36662 166226
rect 36234 166046 36290 166102
rect 36358 166046 36414 166102
rect 36482 166046 36538 166102
rect 36606 166046 36662 166102
rect 36234 165922 36290 165978
rect 36358 165922 36414 165978
rect 36482 165922 36538 165978
rect 36606 165922 36662 165978
rect 36234 148294 36290 148350
rect 36358 148294 36414 148350
rect 36482 148294 36538 148350
rect 36606 148294 36662 148350
rect 36234 148170 36290 148226
rect 36358 148170 36414 148226
rect 36482 148170 36538 148226
rect 36606 148170 36662 148226
rect 36234 148046 36290 148102
rect 36358 148046 36414 148102
rect 36482 148046 36538 148102
rect 36606 148046 36662 148102
rect 36234 147922 36290 147978
rect 36358 147922 36414 147978
rect 36482 147922 36538 147978
rect 36606 147922 36662 147978
rect 36234 130294 36290 130350
rect 36358 130294 36414 130350
rect 36482 130294 36538 130350
rect 36606 130294 36662 130350
rect 36234 130170 36290 130226
rect 36358 130170 36414 130226
rect 36482 130170 36538 130226
rect 36606 130170 36662 130226
rect 36234 130046 36290 130102
rect 36358 130046 36414 130102
rect 36482 130046 36538 130102
rect 36606 130046 36662 130102
rect 36234 129922 36290 129978
rect 36358 129922 36414 129978
rect 36482 129922 36538 129978
rect 36606 129922 36662 129978
rect 36234 112294 36290 112350
rect 36358 112294 36414 112350
rect 36482 112294 36538 112350
rect 36606 112294 36662 112350
rect 36234 112170 36290 112226
rect 36358 112170 36414 112226
rect 36482 112170 36538 112226
rect 36606 112170 36662 112226
rect 36234 112046 36290 112102
rect 36358 112046 36414 112102
rect 36482 112046 36538 112102
rect 36606 112046 36662 112102
rect 36234 111922 36290 111978
rect 36358 111922 36414 111978
rect 36482 111922 36538 111978
rect 36606 111922 36662 111978
rect 36234 94294 36290 94350
rect 36358 94294 36414 94350
rect 36482 94294 36538 94350
rect 36606 94294 36662 94350
rect 36234 94170 36290 94226
rect 36358 94170 36414 94226
rect 36482 94170 36538 94226
rect 36606 94170 36662 94226
rect 36234 94046 36290 94102
rect 36358 94046 36414 94102
rect 36482 94046 36538 94102
rect 36606 94046 36662 94102
rect 36234 93922 36290 93978
rect 36358 93922 36414 93978
rect 36482 93922 36538 93978
rect 36606 93922 36662 93978
rect 36234 76294 36290 76350
rect 36358 76294 36414 76350
rect 36482 76294 36538 76350
rect 36606 76294 36662 76350
rect 36234 76170 36290 76226
rect 36358 76170 36414 76226
rect 36482 76170 36538 76226
rect 36606 76170 36662 76226
rect 36234 76046 36290 76102
rect 36358 76046 36414 76102
rect 36482 76046 36538 76102
rect 36606 76046 36662 76102
rect 36234 75922 36290 75978
rect 36358 75922 36414 75978
rect 36482 75922 36538 75978
rect 36606 75922 36662 75978
rect 36234 58294 36290 58350
rect 36358 58294 36414 58350
rect 36482 58294 36538 58350
rect 36606 58294 36662 58350
rect 36234 58170 36290 58226
rect 36358 58170 36414 58226
rect 36482 58170 36538 58226
rect 36606 58170 36662 58226
rect 36234 58046 36290 58102
rect 36358 58046 36414 58102
rect 36482 58046 36538 58102
rect 36606 58046 36662 58102
rect 36234 57922 36290 57978
rect 36358 57922 36414 57978
rect 36482 57922 36538 57978
rect 36606 57922 36662 57978
rect 36234 40294 36290 40350
rect 36358 40294 36414 40350
rect 36482 40294 36538 40350
rect 36606 40294 36662 40350
rect 36234 40170 36290 40226
rect 36358 40170 36414 40226
rect 36482 40170 36538 40226
rect 36606 40170 36662 40226
rect 36234 40046 36290 40102
rect 36358 40046 36414 40102
rect 36482 40046 36538 40102
rect 36606 40046 36662 40102
rect 36234 39922 36290 39978
rect 36358 39922 36414 39978
rect 36482 39922 36538 39978
rect 36606 39922 36662 39978
rect 36234 22294 36290 22350
rect 36358 22294 36414 22350
rect 36482 22294 36538 22350
rect 36606 22294 36662 22350
rect 36234 22170 36290 22226
rect 36358 22170 36414 22226
rect 36482 22170 36538 22226
rect 36606 22170 36662 22226
rect 36234 22046 36290 22102
rect 36358 22046 36414 22102
rect 36482 22046 36538 22102
rect 36606 22046 36662 22102
rect 36234 21922 36290 21978
rect 36358 21922 36414 21978
rect 36482 21922 36538 21978
rect 36606 21922 36662 21978
rect 39676 4922 39732 4978
rect 39954 208294 40010 208350
rect 40078 208294 40134 208350
rect 40202 208294 40258 208350
rect 40326 208294 40382 208350
rect 39954 208170 40010 208226
rect 40078 208170 40134 208226
rect 40202 208170 40258 208226
rect 40326 208170 40382 208226
rect 39954 208046 40010 208102
rect 40078 208046 40134 208102
rect 40202 208046 40258 208102
rect 40326 208046 40382 208102
rect 39954 207922 40010 207978
rect 40078 207922 40134 207978
rect 40202 207922 40258 207978
rect 40326 207922 40382 207978
rect 39954 190294 40010 190350
rect 40078 190294 40134 190350
rect 40202 190294 40258 190350
rect 40326 190294 40382 190350
rect 39954 190170 40010 190226
rect 40078 190170 40134 190226
rect 40202 190170 40258 190226
rect 40326 190170 40382 190226
rect 39954 190046 40010 190102
rect 40078 190046 40134 190102
rect 40202 190046 40258 190102
rect 40326 190046 40382 190102
rect 39954 189922 40010 189978
rect 40078 189922 40134 189978
rect 40202 189922 40258 189978
rect 40326 189922 40382 189978
rect 39954 172294 40010 172350
rect 40078 172294 40134 172350
rect 40202 172294 40258 172350
rect 40326 172294 40382 172350
rect 39954 172170 40010 172226
rect 40078 172170 40134 172226
rect 40202 172170 40258 172226
rect 40326 172170 40382 172226
rect 39954 172046 40010 172102
rect 40078 172046 40134 172102
rect 40202 172046 40258 172102
rect 40326 172046 40382 172102
rect 39954 171922 40010 171978
rect 40078 171922 40134 171978
rect 40202 171922 40258 171978
rect 40326 171922 40382 171978
rect 39954 154294 40010 154350
rect 40078 154294 40134 154350
rect 40202 154294 40258 154350
rect 40326 154294 40382 154350
rect 39954 154170 40010 154226
rect 40078 154170 40134 154226
rect 40202 154170 40258 154226
rect 40326 154170 40382 154226
rect 39954 154046 40010 154102
rect 40078 154046 40134 154102
rect 40202 154046 40258 154102
rect 40326 154046 40382 154102
rect 39954 153922 40010 153978
rect 40078 153922 40134 153978
rect 40202 153922 40258 153978
rect 40326 153922 40382 153978
rect 39954 136294 40010 136350
rect 40078 136294 40134 136350
rect 40202 136294 40258 136350
rect 40326 136294 40382 136350
rect 39954 136170 40010 136226
rect 40078 136170 40134 136226
rect 40202 136170 40258 136226
rect 40326 136170 40382 136226
rect 39954 136046 40010 136102
rect 40078 136046 40134 136102
rect 40202 136046 40258 136102
rect 40326 136046 40382 136102
rect 39954 135922 40010 135978
rect 40078 135922 40134 135978
rect 40202 135922 40258 135978
rect 40326 135922 40382 135978
rect 39954 118294 40010 118350
rect 40078 118294 40134 118350
rect 40202 118294 40258 118350
rect 40326 118294 40382 118350
rect 39954 118170 40010 118226
rect 40078 118170 40134 118226
rect 40202 118170 40258 118226
rect 40326 118170 40382 118226
rect 39954 118046 40010 118102
rect 40078 118046 40134 118102
rect 40202 118046 40258 118102
rect 40326 118046 40382 118102
rect 39954 117922 40010 117978
rect 40078 117922 40134 117978
rect 40202 117922 40258 117978
rect 40326 117922 40382 117978
rect 39954 100294 40010 100350
rect 40078 100294 40134 100350
rect 40202 100294 40258 100350
rect 40326 100294 40382 100350
rect 39954 100170 40010 100226
rect 40078 100170 40134 100226
rect 40202 100170 40258 100226
rect 40326 100170 40382 100226
rect 39954 100046 40010 100102
rect 40078 100046 40134 100102
rect 40202 100046 40258 100102
rect 40326 100046 40382 100102
rect 39954 99922 40010 99978
rect 40078 99922 40134 99978
rect 40202 99922 40258 99978
rect 40326 99922 40382 99978
rect 39954 82294 40010 82350
rect 40078 82294 40134 82350
rect 40202 82294 40258 82350
rect 40326 82294 40382 82350
rect 39954 82170 40010 82226
rect 40078 82170 40134 82226
rect 40202 82170 40258 82226
rect 40326 82170 40382 82226
rect 39954 82046 40010 82102
rect 40078 82046 40134 82102
rect 40202 82046 40258 82102
rect 40326 82046 40382 82102
rect 39954 81922 40010 81978
rect 40078 81922 40134 81978
rect 40202 81922 40258 81978
rect 40326 81922 40382 81978
rect 39954 64294 40010 64350
rect 40078 64294 40134 64350
rect 40202 64294 40258 64350
rect 40326 64294 40382 64350
rect 39954 64170 40010 64226
rect 40078 64170 40134 64226
rect 40202 64170 40258 64226
rect 40326 64170 40382 64226
rect 39954 64046 40010 64102
rect 40078 64046 40134 64102
rect 40202 64046 40258 64102
rect 40326 64046 40382 64102
rect 39954 63922 40010 63978
rect 40078 63922 40134 63978
rect 40202 63922 40258 63978
rect 40326 63922 40382 63978
rect 39954 46294 40010 46350
rect 40078 46294 40134 46350
rect 40202 46294 40258 46350
rect 40326 46294 40382 46350
rect 39954 46170 40010 46226
rect 40078 46170 40134 46226
rect 40202 46170 40258 46226
rect 40326 46170 40382 46226
rect 39954 46046 40010 46102
rect 40078 46046 40134 46102
rect 40202 46046 40258 46102
rect 40326 46046 40382 46102
rect 39954 45922 40010 45978
rect 40078 45922 40134 45978
rect 40202 45922 40258 45978
rect 40326 45922 40382 45978
rect 39954 28294 40010 28350
rect 40078 28294 40134 28350
rect 40202 28294 40258 28350
rect 40326 28294 40382 28350
rect 39954 28170 40010 28226
rect 40078 28170 40134 28226
rect 40202 28170 40258 28226
rect 40326 28170 40382 28226
rect 39954 28046 40010 28102
rect 40078 28046 40134 28102
rect 40202 28046 40258 28102
rect 40326 28046 40382 28102
rect 39954 27922 40010 27978
rect 40078 27922 40134 27978
rect 40202 27922 40258 27978
rect 40326 27922 40382 27978
rect 39954 10294 40010 10350
rect 40078 10294 40134 10350
rect 40202 10294 40258 10350
rect 40326 10294 40382 10350
rect 39954 10170 40010 10226
rect 40078 10170 40134 10226
rect 40202 10170 40258 10226
rect 40326 10170 40382 10226
rect 39954 10046 40010 10102
rect 40078 10046 40134 10102
rect 40202 10046 40258 10102
rect 40326 10046 40382 10102
rect 39954 9922 40010 9978
rect 40078 9922 40134 9978
rect 40202 9922 40258 9978
rect 40326 9922 40382 9978
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 9234 -1176 9290 -1120
rect 9358 -1176 9414 -1120
rect 9482 -1176 9538 -1120
rect 9606 -1176 9662 -1120
rect 9234 -1300 9290 -1244
rect 9358 -1300 9414 -1244
rect 9482 -1300 9538 -1244
rect 9606 -1300 9662 -1244
rect 9234 -1424 9290 -1368
rect 9358 -1424 9414 -1368
rect 9482 -1424 9538 -1368
rect 9606 -1424 9662 -1368
rect 9234 -1548 9290 -1492
rect 9358 -1548 9414 -1492
rect 9482 -1548 9538 -1492
rect 9606 -1548 9662 -1492
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 41356 234422 41412 234478
rect 44518 202294 44574 202350
rect 44642 202294 44698 202350
rect 44518 202170 44574 202226
rect 44642 202170 44698 202226
rect 44518 202046 44574 202102
rect 44642 202046 44698 202102
rect 44518 201922 44574 201978
rect 44642 201922 44698 201978
rect 44518 184294 44574 184350
rect 44642 184294 44698 184350
rect 44518 184170 44574 184226
rect 44642 184170 44698 184226
rect 44518 184046 44574 184102
rect 44642 184046 44698 184102
rect 44518 183922 44574 183978
rect 44642 183922 44698 183978
rect 44518 166294 44574 166350
rect 44642 166294 44698 166350
rect 44518 166170 44574 166226
rect 44642 166170 44698 166226
rect 44518 166046 44574 166102
rect 44642 166046 44698 166102
rect 44518 165922 44574 165978
rect 44642 165922 44698 165978
rect 44518 148294 44574 148350
rect 44642 148294 44698 148350
rect 44518 148170 44574 148226
rect 44642 148170 44698 148226
rect 44518 148046 44574 148102
rect 44642 148046 44698 148102
rect 44518 147922 44574 147978
rect 44642 147922 44698 147978
rect 44518 130294 44574 130350
rect 44642 130294 44698 130350
rect 44518 130170 44574 130226
rect 44642 130170 44698 130226
rect 44518 130046 44574 130102
rect 44642 130046 44698 130102
rect 44518 129922 44574 129978
rect 44642 129922 44698 129978
rect 44518 112294 44574 112350
rect 44642 112294 44698 112350
rect 44518 112170 44574 112226
rect 44642 112170 44698 112226
rect 44518 112046 44574 112102
rect 44642 112046 44698 112102
rect 44518 111922 44574 111978
rect 44642 111922 44698 111978
rect 44518 94294 44574 94350
rect 44642 94294 44698 94350
rect 44518 94170 44574 94226
rect 44642 94170 44698 94226
rect 44518 94046 44574 94102
rect 44642 94046 44698 94102
rect 44518 93922 44574 93978
rect 44642 93922 44698 93978
rect 44518 76294 44574 76350
rect 44642 76294 44698 76350
rect 44518 76170 44574 76226
rect 44642 76170 44698 76226
rect 44518 76046 44574 76102
rect 44642 76046 44698 76102
rect 44518 75922 44574 75978
rect 44642 75922 44698 75978
rect 44518 58294 44574 58350
rect 44642 58294 44698 58350
rect 44518 58170 44574 58226
rect 44642 58170 44698 58226
rect 44518 58046 44574 58102
rect 44642 58046 44698 58102
rect 44518 57922 44574 57978
rect 44642 57922 44698 57978
rect 66954 238294 67010 238350
rect 67078 238294 67134 238350
rect 67202 238294 67258 238350
rect 67326 238294 67382 238350
rect 66954 238170 67010 238226
rect 67078 238170 67134 238226
rect 67202 238170 67258 238226
rect 67326 238170 67382 238226
rect 66954 238046 67010 238102
rect 67078 238046 67134 238102
rect 67202 238046 67258 238102
rect 67326 238046 67382 238102
rect 66954 237922 67010 237978
rect 67078 237922 67134 237978
rect 67202 237922 67258 237978
rect 67326 237922 67382 237978
rect 49644 206522 49700 206578
rect 49532 164582 49588 164638
rect 66954 220294 67010 220350
rect 67078 220294 67134 220350
rect 67202 220294 67258 220350
rect 67326 220294 67382 220350
rect 66954 220170 67010 220226
rect 67078 220170 67134 220226
rect 67202 220170 67258 220226
rect 67326 220170 67382 220226
rect 66954 220046 67010 220102
rect 67078 220046 67134 220102
rect 67202 220046 67258 220102
rect 67326 220046 67382 220102
rect 66954 219922 67010 219978
rect 67078 219922 67134 219978
rect 67202 219922 67258 219978
rect 67326 219922 67382 219978
rect 70674 244294 70730 244350
rect 70798 244294 70854 244350
rect 70922 244294 70978 244350
rect 71046 244294 71102 244350
rect 70674 244170 70730 244226
rect 70798 244170 70854 244226
rect 70922 244170 70978 244226
rect 71046 244170 71102 244226
rect 70674 244046 70730 244102
rect 70798 244046 70854 244102
rect 70922 244046 70978 244102
rect 71046 244046 71102 244102
rect 70674 243922 70730 243978
rect 70798 243922 70854 243978
rect 70922 243922 70978 243978
rect 71046 243922 71102 243978
rect 90598 244294 90654 244350
rect 90722 244294 90778 244350
rect 90598 244170 90654 244226
rect 90722 244170 90778 244226
rect 90598 244046 90654 244102
rect 90722 244046 90778 244102
rect 90598 243922 90654 243978
rect 90722 243922 90778 243978
rect 97674 238294 97730 238350
rect 97798 238294 97854 238350
rect 97922 238294 97978 238350
rect 98046 238294 98102 238350
rect 76972 237662 77028 237718
rect 97674 238170 97730 238226
rect 97798 238170 97854 238226
rect 97922 238170 97978 238226
rect 98046 238170 98102 238226
rect 97674 238046 97730 238102
rect 97798 238046 97854 238102
rect 97922 238046 97978 238102
rect 98046 238046 98102 238102
rect 97674 237922 97730 237978
rect 97798 237922 97854 237978
rect 97922 237922 97978 237978
rect 98046 237922 98102 237978
rect 72940 237482 72996 237538
rect 70674 226294 70730 226350
rect 70798 226294 70854 226350
rect 70922 226294 70978 226350
rect 71046 226294 71102 226350
rect 70674 226170 70730 226226
rect 70798 226170 70854 226226
rect 70922 226170 70978 226226
rect 71046 226170 71102 226226
rect 70674 226046 70730 226102
rect 70798 226046 70854 226102
rect 70922 226046 70978 226102
rect 71046 226046 71102 226102
rect 70674 225922 70730 225978
rect 70798 225922 70854 225978
rect 70922 225922 70978 225978
rect 71046 225922 71102 225978
rect 99932 237482 99988 237538
rect 128394 472294 128450 472350
rect 128518 472294 128574 472350
rect 128642 472294 128698 472350
rect 128766 472294 128822 472350
rect 128394 472170 128450 472226
rect 128518 472170 128574 472226
rect 128642 472170 128698 472226
rect 128766 472170 128822 472226
rect 128394 472046 128450 472102
rect 128518 472046 128574 472102
rect 128642 472046 128698 472102
rect 128766 472046 128822 472102
rect 128394 471922 128450 471978
rect 128518 471922 128574 471978
rect 128642 471922 128698 471978
rect 128766 471922 128822 471978
rect 128394 454294 128450 454350
rect 128518 454294 128574 454350
rect 128642 454294 128698 454350
rect 128766 454294 128822 454350
rect 128394 454170 128450 454226
rect 128518 454170 128574 454226
rect 128642 454170 128698 454226
rect 128766 454170 128822 454226
rect 128394 454046 128450 454102
rect 128518 454046 128574 454102
rect 128642 454046 128698 454102
rect 128766 454046 128822 454102
rect 128394 453922 128450 453978
rect 128518 453922 128574 453978
rect 128642 453922 128698 453978
rect 128766 453922 128822 453978
rect 128394 436294 128450 436350
rect 128518 436294 128574 436350
rect 128642 436294 128698 436350
rect 128766 436294 128822 436350
rect 128394 436170 128450 436226
rect 128518 436170 128574 436226
rect 128642 436170 128698 436226
rect 128766 436170 128822 436226
rect 128394 436046 128450 436102
rect 128518 436046 128574 436102
rect 128642 436046 128698 436102
rect 128766 436046 128822 436102
rect 128394 435922 128450 435978
rect 128518 435922 128574 435978
rect 128642 435922 128698 435978
rect 128766 435922 128822 435978
rect 128394 418294 128450 418350
rect 128518 418294 128574 418350
rect 128642 418294 128698 418350
rect 128766 418294 128822 418350
rect 128394 418170 128450 418226
rect 128518 418170 128574 418226
rect 128642 418170 128698 418226
rect 128766 418170 128822 418226
rect 128394 418046 128450 418102
rect 128518 418046 128574 418102
rect 128642 418046 128698 418102
rect 128766 418046 128822 418102
rect 128394 417922 128450 417978
rect 128518 417922 128574 417978
rect 128642 417922 128698 417978
rect 128766 417922 128822 417978
rect 128394 400294 128450 400350
rect 128518 400294 128574 400350
rect 128642 400294 128698 400350
rect 128766 400294 128822 400350
rect 128394 400170 128450 400226
rect 128518 400170 128574 400226
rect 128642 400170 128698 400226
rect 128766 400170 128822 400226
rect 128394 400046 128450 400102
rect 128518 400046 128574 400102
rect 128642 400046 128698 400102
rect 128766 400046 128822 400102
rect 128394 399922 128450 399978
rect 128518 399922 128574 399978
rect 128642 399922 128698 399978
rect 128766 399922 128822 399978
rect 101394 370294 101450 370350
rect 101518 370294 101574 370350
rect 101642 370294 101698 370350
rect 101766 370294 101822 370350
rect 101394 370170 101450 370226
rect 101518 370170 101574 370226
rect 101642 370170 101698 370226
rect 101766 370170 101822 370226
rect 101394 370046 101450 370102
rect 101518 370046 101574 370102
rect 101642 370046 101698 370102
rect 101766 370046 101822 370102
rect 101394 369922 101450 369978
rect 101518 369922 101574 369978
rect 101642 369922 101698 369978
rect 101766 369922 101822 369978
rect 101394 352294 101450 352350
rect 101518 352294 101574 352350
rect 101642 352294 101698 352350
rect 101766 352294 101822 352350
rect 101394 352170 101450 352226
rect 101518 352170 101574 352226
rect 101642 352170 101698 352226
rect 101766 352170 101822 352226
rect 101394 352046 101450 352102
rect 101518 352046 101574 352102
rect 101642 352046 101698 352102
rect 101766 352046 101822 352102
rect 101394 351922 101450 351978
rect 101518 351922 101574 351978
rect 101642 351922 101698 351978
rect 101766 351922 101822 351978
rect 101394 334294 101450 334350
rect 101518 334294 101574 334350
rect 101642 334294 101698 334350
rect 101766 334294 101822 334350
rect 101394 334170 101450 334226
rect 101518 334170 101574 334226
rect 101642 334170 101698 334226
rect 101766 334170 101822 334226
rect 101394 334046 101450 334102
rect 101518 334046 101574 334102
rect 101642 334046 101698 334102
rect 101766 334046 101822 334102
rect 101394 333922 101450 333978
rect 101518 333922 101574 333978
rect 101642 333922 101698 333978
rect 101766 333922 101822 333978
rect 101394 316294 101450 316350
rect 101518 316294 101574 316350
rect 101642 316294 101698 316350
rect 101766 316294 101822 316350
rect 101394 316170 101450 316226
rect 101518 316170 101574 316226
rect 101642 316170 101698 316226
rect 101766 316170 101822 316226
rect 101394 316046 101450 316102
rect 101518 316046 101574 316102
rect 101642 316046 101698 316102
rect 101766 316046 101822 316102
rect 101394 315922 101450 315978
rect 101518 315922 101574 315978
rect 101642 315922 101698 315978
rect 101766 315922 101822 315978
rect 101394 298294 101450 298350
rect 101518 298294 101574 298350
rect 101642 298294 101698 298350
rect 101766 298294 101822 298350
rect 101394 298170 101450 298226
rect 101518 298170 101574 298226
rect 101642 298170 101698 298226
rect 101766 298170 101822 298226
rect 101394 298046 101450 298102
rect 101518 298046 101574 298102
rect 101642 298046 101698 298102
rect 101766 298046 101822 298102
rect 101394 297922 101450 297978
rect 101518 297922 101574 297978
rect 101642 297922 101698 297978
rect 101766 297922 101822 297978
rect 101394 280294 101450 280350
rect 101518 280294 101574 280350
rect 101642 280294 101698 280350
rect 101766 280294 101822 280350
rect 101394 280170 101450 280226
rect 101518 280170 101574 280226
rect 101642 280170 101698 280226
rect 101766 280170 101822 280226
rect 101394 280046 101450 280102
rect 101518 280046 101574 280102
rect 101642 280046 101698 280102
rect 101766 280046 101822 280102
rect 101394 279922 101450 279978
rect 101518 279922 101574 279978
rect 101642 279922 101698 279978
rect 101766 279922 101822 279978
rect 101394 262294 101450 262350
rect 101518 262294 101574 262350
rect 101642 262294 101698 262350
rect 101766 262294 101822 262350
rect 101394 262170 101450 262226
rect 101518 262170 101574 262226
rect 101642 262170 101698 262226
rect 101766 262170 101822 262226
rect 101394 262046 101450 262102
rect 101518 262046 101574 262102
rect 101642 262046 101698 262102
rect 101766 262046 101822 262102
rect 101394 261922 101450 261978
rect 101518 261922 101574 261978
rect 101642 261922 101698 261978
rect 101766 261922 101822 261978
rect 101394 244294 101450 244350
rect 101518 244294 101574 244350
rect 101642 244294 101698 244350
rect 101766 244294 101822 244350
rect 101394 244170 101450 244226
rect 101518 244170 101574 244226
rect 101642 244170 101698 244226
rect 101766 244170 101822 244226
rect 101394 244046 101450 244102
rect 101518 244046 101574 244102
rect 101642 244046 101698 244102
rect 101766 244046 101822 244102
rect 101394 243922 101450 243978
rect 101518 243922 101574 243978
rect 101642 243922 101698 243978
rect 101766 243922 101822 243978
rect 97674 220294 97730 220350
rect 97798 220294 97854 220350
rect 97922 220294 97978 220350
rect 98046 220294 98102 220350
rect 97674 220170 97730 220226
rect 97798 220170 97854 220226
rect 97922 220170 97978 220226
rect 98046 220170 98102 220226
rect 97674 220046 97730 220102
rect 97798 220046 97854 220102
rect 97922 220046 97978 220102
rect 98046 220046 98102 220102
rect 97674 219922 97730 219978
rect 97798 219922 97854 219978
rect 97922 219922 97978 219978
rect 98046 219922 98102 219978
rect 128394 382294 128450 382350
rect 128518 382294 128574 382350
rect 128642 382294 128698 382350
rect 128766 382294 128822 382350
rect 128394 382170 128450 382226
rect 128518 382170 128574 382226
rect 128642 382170 128698 382226
rect 128766 382170 128822 382226
rect 128394 382046 128450 382102
rect 128518 382046 128574 382102
rect 128642 382046 128698 382102
rect 128766 382046 128822 382102
rect 128394 381922 128450 381978
rect 128518 381922 128574 381978
rect 128642 381922 128698 381978
rect 128766 381922 128822 381978
rect 128394 364294 128450 364350
rect 128518 364294 128574 364350
rect 128642 364294 128698 364350
rect 128766 364294 128822 364350
rect 128394 364170 128450 364226
rect 128518 364170 128574 364226
rect 128642 364170 128698 364226
rect 128766 364170 128822 364226
rect 128394 364046 128450 364102
rect 128518 364046 128574 364102
rect 128642 364046 128698 364102
rect 128766 364046 128822 364102
rect 128394 363922 128450 363978
rect 128518 363922 128574 363978
rect 128642 363922 128698 363978
rect 128766 363922 128822 363978
rect 128394 346294 128450 346350
rect 128518 346294 128574 346350
rect 128642 346294 128698 346350
rect 128766 346294 128822 346350
rect 128394 346170 128450 346226
rect 128518 346170 128574 346226
rect 128642 346170 128698 346226
rect 128766 346170 128822 346226
rect 128394 346046 128450 346102
rect 128518 346046 128574 346102
rect 128642 346046 128698 346102
rect 128766 346046 128822 346102
rect 128394 345922 128450 345978
rect 128518 345922 128574 345978
rect 128642 345922 128698 345978
rect 128766 345922 128822 345978
rect 128394 328294 128450 328350
rect 128518 328294 128574 328350
rect 128642 328294 128698 328350
rect 128766 328294 128822 328350
rect 128394 328170 128450 328226
rect 128518 328170 128574 328226
rect 128642 328170 128698 328226
rect 128766 328170 128822 328226
rect 128394 328046 128450 328102
rect 128518 328046 128574 328102
rect 128642 328046 128698 328102
rect 128766 328046 128822 328102
rect 128394 327922 128450 327978
rect 128518 327922 128574 327978
rect 128642 327922 128698 327978
rect 128766 327922 128822 327978
rect 128394 310294 128450 310350
rect 128518 310294 128574 310350
rect 128642 310294 128698 310350
rect 128766 310294 128822 310350
rect 128394 310170 128450 310226
rect 128518 310170 128574 310226
rect 128642 310170 128698 310226
rect 128766 310170 128822 310226
rect 128394 310046 128450 310102
rect 128518 310046 128574 310102
rect 128642 310046 128698 310102
rect 128766 310046 128822 310102
rect 128394 309922 128450 309978
rect 128518 309922 128574 309978
rect 128642 309922 128698 309978
rect 128766 309922 128822 309978
rect 128394 292294 128450 292350
rect 128518 292294 128574 292350
rect 128642 292294 128698 292350
rect 128766 292294 128822 292350
rect 128394 292170 128450 292226
rect 128518 292170 128574 292226
rect 128642 292170 128698 292226
rect 128766 292170 128822 292226
rect 128394 292046 128450 292102
rect 128518 292046 128574 292102
rect 128642 292046 128698 292102
rect 128766 292046 128822 292102
rect 128394 291922 128450 291978
rect 128518 291922 128574 291978
rect 128642 291922 128698 291978
rect 128766 291922 128822 291978
rect 110012 237662 110068 237718
rect 101394 226294 101450 226350
rect 101518 226294 101574 226350
rect 101642 226294 101698 226350
rect 101766 226294 101822 226350
rect 101394 226170 101450 226226
rect 101518 226170 101574 226226
rect 101642 226170 101698 226226
rect 101766 226170 101822 226226
rect 101394 226046 101450 226102
rect 101518 226046 101574 226102
rect 101642 226046 101698 226102
rect 101766 226046 101822 226102
rect 101394 225922 101450 225978
rect 101518 225922 101574 225978
rect 101642 225922 101698 225978
rect 101766 225922 101822 225978
rect 128394 274294 128450 274350
rect 128518 274294 128574 274350
rect 128642 274294 128698 274350
rect 128766 274294 128822 274350
rect 128394 274170 128450 274226
rect 128518 274170 128574 274226
rect 128642 274170 128698 274226
rect 128766 274170 128822 274226
rect 128394 274046 128450 274102
rect 128518 274046 128574 274102
rect 128642 274046 128698 274102
rect 128766 274046 128822 274102
rect 128394 273922 128450 273978
rect 128518 273922 128574 273978
rect 128642 273922 128698 273978
rect 128766 273922 128822 273978
rect 128394 256294 128450 256350
rect 128518 256294 128574 256350
rect 128642 256294 128698 256350
rect 128766 256294 128822 256350
rect 128394 256170 128450 256226
rect 128518 256170 128574 256226
rect 128642 256170 128698 256226
rect 128766 256170 128822 256226
rect 128394 256046 128450 256102
rect 128518 256046 128574 256102
rect 128642 256046 128698 256102
rect 128766 256046 128822 256102
rect 128394 255922 128450 255978
rect 128518 255922 128574 255978
rect 128642 255922 128698 255978
rect 128766 255922 128822 255978
rect 128394 238294 128450 238350
rect 128518 238294 128574 238350
rect 128642 238294 128698 238350
rect 128766 238294 128822 238350
rect 128394 238170 128450 238226
rect 128518 238170 128574 238226
rect 128642 238170 128698 238226
rect 128766 238170 128822 238226
rect 128394 238046 128450 238102
rect 128518 238046 128574 238102
rect 128642 238046 128698 238102
rect 128766 238046 128822 238102
rect 128394 237922 128450 237978
rect 128518 237922 128574 237978
rect 128642 237922 128698 237978
rect 128766 237922 128822 237978
rect 128394 220294 128450 220350
rect 128518 220294 128574 220350
rect 128642 220294 128698 220350
rect 128766 220294 128822 220350
rect 128394 220170 128450 220226
rect 128518 220170 128574 220226
rect 128642 220170 128698 220226
rect 128766 220170 128822 220226
rect 128394 220046 128450 220102
rect 128518 220046 128574 220102
rect 128642 220046 128698 220102
rect 128766 220046 128822 220102
rect 128394 219922 128450 219978
rect 128518 219922 128574 219978
rect 128642 219922 128698 219978
rect 128766 219922 128822 219978
rect 132114 478294 132170 478350
rect 132238 478294 132294 478350
rect 132362 478294 132418 478350
rect 132486 478294 132542 478350
rect 132114 478170 132170 478226
rect 132238 478170 132294 478226
rect 132362 478170 132418 478226
rect 132486 478170 132542 478226
rect 132114 478046 132170 478102
rect 132238 478046 132294 478102
rect 132362 478046 132418 478102
rect 132486 478046 132542 478102
rect 132114 477922 132170 477978
rect 132238 477922 132294 477978
rect 132362 477922 132418 477978
rect 132486 477922 132542 477978
rect 132114 460294 132170 460350
rect 132238 460294 132294 460350
rect 132362 460294 132418 460350
rect 132486 460294 132542 460350
rect 132114 460170 132170 460226
rect 132238 460170 132294 460226
rect 132362 460170 132418 460226
rect 132486 460170 132542 460226
rect 132114 460046 132170 460102
rect 132238 460046 132294 460102
rect 132362 460046 132418 460102
rect 132486 460046 132542 460102
rect 132114 459922 132170 459978
rect 132238 459922 132294 459978
rect 132362 459922 132418 459978
rect 132486 459922 132542 459978
rect 132114 442294 132170 442350
rect 132238 442294 132294 442350
rect 132362 442294 132418 442350
rect 132486 442294 132542 442350
rect 132114 442170 132170 442226
rect 132238 442170 132294 442226
rect 132362 442170 132418 442226
rect 132486 442170 132542 442226
rect 132114 442046 132170 442102
rect 132238 442046 132294 442102
rect 132362 442046 132418 442102
rect 132486 442046 132542 442102
rect 132114 441922 132170 441978
rect 132238 441922 132294 441978
rect 132362 441922 132418 441978
rect 132486 441922 132542 441978
rect 132114 424294 132170 424350
rect 132238 424294 132294 424350
rect 132362 424294 132418 424350
rect 132486 424294 132542 424350
rect 132114 424170 132170 424226
rect 132238 424170 132294 424226
rect 132362 424170 132418 424226
rect 132486 424170 132542 424226
rect 132114 424046 132170 424102
rect 132238 424046 132294 424102
rect 132362 424046 132418 424102
rect 132486 424046 132542 424102
rect 132114 423922 132170 423978
rect 132238 423922 132294 423978
rect 132362 423922 132418 423978
rect 132486 423922 132542 423978
rect 132114 406294 132170 406350
rect 132238 406294 132294 406350
rect 132362 406294 132418 406350
rect 132486 406294 132542 406350
rect 132114 406170 132170 406226
rect 132238 406170 132294 406226
rect 132362 406170 132418 406226
rect 132486 406170 132542 406226
rect 132114 406046 132170 406102
rect 132238 406046 132294 406102
rect 132362 406046 132418 406102
rect 132486 406046 132542 406102
rect 132114 405922 132170 405978
rect 132238 405922 132294 405978
rect 132362 405922 132418 405978
rect 132486 405922 132542 405978
rect 132114 388294 132170 388350
rect 132238 388294 132294 388350
rect 132362 388294 132418 388350
rect 132486 388294 132542 388350
rect 132114 388170 132170 388226
rect 132238 388170 132294 388226
rect 132362 388170 132418 388226
rect 132486 388170 132542 388226
rect 132114 388046 132170 388102
rect 132238 388046 132294 388102
rect 132362 388046 132418 388102
rect 132486 388046 132542 388102
rect 132114 387922 132170 387978
rect 132238 387922 132294 387978
rect 132362 387922 132418 387978
rect 132486 387922 132542 387978
rect 132114 370294 132170 370350
rect 132238 370294 132294 370350
rect 132362 370294 132418 370350
rect 132486 370294 132542 370350
rect 132114 370170 132170 370226
rect 132238 370170 132294 370226
rect 132362 370170 132418 370226
rect 132486 370170 132542 370226
rect 132114 370046 132170 370102
rect 132238 370046 132294 370102
rect 132362 370046 132418 370102
rect 132486 370046 132542 370102
rect 132114 369922 132170 369978
rect 132238 369922 132294 369978
rect 132362 369922 132418 369978
rect 132486 369922 132542 369978
rect 159114 490294 159170 490350
rect 159238 490294 159294 490350
rect 159362 490294 159418 490350
rect 159486 490294 159542 490350
rect 159114 490170 159170 490226
rect 159238 490170 159294 490226
rect 159362 490170 159418 490226
rect 159486 490170 159542 490226
rect 159114 490046 159170 490102
rect 159238 490046 159294 490102
rect 159362 490046 159418 490102
rect 159486 490046 159542 490102
rect 159114 489922 159170 489978
rect 159238 489922 159294 489978
rect 159362 489922 159418 489978
rect 159486 489922 159542 489978
rect 159114 472294 159170 472350
rect 159238 472294 159294 472350
rect 159362 472294 159418 472350
rect 159486 472294 159542 472350
rect 159114 472170 159170 472226
rect 159238 472170 159294 472226
rect 159362 472170 159418 472226
rect 159486 472170 159542 472226
rect 159114 472046 159170 472102
rect 159238 472046 159294 472102
rect 159362 472046 159418 472102
rect 159486 472046 159542 472102
rect 159114 471922 159170 471978
rect 159238 471922 159294 471978
rect 159362 471922 159418 471978
rect 159486 471922 159542 471978
rect 159114 454294 159170 454350
rect 159238 454294 159294 454350
rect 159362 454294 159418 454350
rect 159486 454294 159542 454350
rect 159114 454170 159170 454226
rect 159238 454170 159294 454226
rect 159362 454170 159418 454226
rect 159486 454170 159542 454226
rect 159114 454046 159170 454102
rect 159238 454046 159294 454102
rect 159362 454046 159418 454102
rect 159486 454046 159542 454102
rect 159114 453922 159170 453978
rect 159238 453922 159294 453978
rect 159362 453922 159418 453978
rect 159486 453922 159542 453978
rect 159114 436294 159170 436350
rect 159238 436294 159294 436350
rect 159362 436294 159418 436350
rect 159486 436294 159542 436350
rect 159114 436170 159170 436226
rect 159238 436170 159294 436226
rect 159362 436170 159418 436226
rect 159486 436170 159542 436226
rect 159114 436046 159170 436102
rect 159238 436046 159294 436102
rect 159362 436046 159418 436102
rect 159486 436046 159542 436102
rect 159114 435922 159170 435978
rect 159238 435922 159294 435978
rect 159362 435922 159418 435978
rect 159486 435922 159542 435978
rect 159114 418294 159170 418350
rect 159238 418294 159294 418350
rect 159362 418294 159418 418350
rect 159486 418294 159542 418350
rect 159114 418170 159170 418226
rect 159238 418170 159294 418226
rect 159362 418170 159418 418226
rect 159486 418170 159542 418226
rect 159114 418046 159170 418102
rect 159238 418046 159294 418102
rect 159362 418046 159418 418102
rect 159486 418046 159542 418102
rect 159114 417922 159170 417978
rect 159238 417922 159294 417978
rect 159362 417922 159418 417978
rect 159486 417922 159542 417978
rect 159114 400294 159170 400350
rect 159238 400294 159294 400350
rect 159362 400294 159418 400350
rect 159486 400294 159542 400350
rect 159114 400170 159170 400226
rect 159238 400170 159294 400226
rect 159362 400170 159418 400226
rect 159486 400170 159542 400226
rect 159114 400046 159170 400102
rect 159238 400046 159294 400102
rect 159362 400046 159418 400102
rect 159486 400046 159542 400102
rect 159114 399922 159170 399978
rect 159238 399922 159294 399978
rect 159362 399922 159418 399978
rect 159486 399922 159542 399978
rect 159114 382294 159170 382350
rect 159238 382294 159294 382350
rect 159362 382294 159418 382350
rect 159486 382294 159542 382350
rect 159114 382170 159170 382226
rect 159238 382170 159294 382226
rect 159362 382170 159418 382226
rect 159486 382170 159542 382226
rect 159114 382046 159170 382102
rect 159238 382046 159294 382102
rect 159362 382046 159418 382102
rect 159486 382046 159542 382102
rect 159114 381922 159170 381978
rect 159238 381922 159294 381978
rect 159362 381922 159418 381978
rect 159486 381922 159542 381978
rect 159114 364360 159170 364416
rect 159238 364360 159294 364416
rect 159362 364360 159418 364416
rect 159486 364360 159542 364416
rect 159114 364236 159170 364292
rect 159238 364236 159294 364292
rect 159362 364236 159418 364292
rect 159486 364236 159542 364292
rect 162834 598116 162890 598172
rect 162958 598116 163014 598172
rect 163082 598116 163138 598172
rect 163206 598116 163262 598172
rect 162834 597992 162890 598048
rect 162958 597992 163014 598048
rect 163082 597992 163138 598048
rect 163206 597992 163262 598048
rect 162834 597868 162890 597924
rect 162958 597868 163014 597924
rect 163082 597868 163138 597924
rect 163206 597868 163262 597924
rect 162834 597744 162890 597800
rect 162958 597744 163014 597800
rect 163082 597744 163138 597800
rect 163206 597744 163262 597800
rect 162834 586294 162890 586350
rect 162958 586294 163014 586350
rect 163082 586294 163138 586350
rect 163206 586294 163262 586350
rect 162834 586170 162890 586226
rect 162958 586170 163014 586226
rect 163082 586170 163138 586226
rect 163206 586170 163262 586226
rect 162834 586046 162890 586102
rect 162958 586046 163014 586102
rect 163082 586046 163138 586102
rect 163206 586046 163262 586102
rect 162834 585922 162890 585978
rect 162958 585922 163014 585978
rect 163082 585922 163138 585978
rect 163206 585922 163262 585978
rect 189834 597156 189890 597212
rect 189958 597156 190014 597212
rect 190082 597156 190138 597212
rect 190206 597156 190262 597212
rect 189834 597032 189890 597088
rect 189958 597032 190014 597088
rect 190082 597032 190138 597088
rect 190206 597032 190262 597088
rect 189834 596908 189890 596964
rect 189958 596908 190014 596964
rect 190082 596908 190138 596964
rect 190206 596908 190262 596964
rect 189834 596784 189890 596840
rect 189958 596784 190014 596840
rect 190082 596784 190138 596840
rect 190206 596784 190262 596840
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 189834 580294 189890 580350
rect 189958 580294 190014 580350
rect 190082 580294 190138 580350
rect 190206 580294 190262 580350
rect 189834 580170 189890 580226
rect 189958 580170 190014 580226
rect 190082 580170 190138 580226
rect 190206 580170 190262 580226
rect 189834 580046 189890 580102
rect 189958 580046 190014 580102
rect 190082 580046 190138 580102
rect 190206 580046 190262 580102
rect 189834 579922 189890 579978
rect 189958 579922 190014 579978
rect 190082 579922 190138 579978
rect 190206 579922 190262 579978
rect 162834 568294 162890 568350
rect 162958 568294 163014 568350
rect 163082 568294 163138 568350
rect 163206 568294 163262 568350
rect 162834 568170 162890 568226
rect 162958 568170 163014 568226
rect 163082 568170 163138 568226
rect 163206 568170 163262 568226
rect 162834 568046 162890 568102
rect 162958 568046 163014 568102
rect 163082 568046 163138 568102
rect 163206 568046 163262 568102
rect 162834 567922 162890 567978
rect 162958 567922 163014 567978
rect 163082 567922 163138 567978
rect 163206 567922 163262 567978
rect 162834 550294 162890 550350
rect 162958 550294 163014 550350
rect 163082 550294 163138 550350
rect 163206 550294 163262 550350
rect 162834 550170 162890 550226
rect 162958 550170 163014 550226
rect 163082 550170 163138 550226
rect 163206 550170 163262 550226
rect 162834 550046 162890 550102
rect 162958 550046 163014 550102
rect 163082 550046 163138 550102
rect 163206 550046 163262 550102
rect 162834 549922 162890 549978
rect 162958 549922 163014 549978
rect 163082 549922 163138 549978
rect 163206 549922 163262 549978
rect 162834 532294 162890 532350
rect 162958 532294 163014 532350
rect 163082 532294 163138 532350
rect 163206 532294 163262 532350
rect 162834 532170 162890 532226
rect 162958 532170 163014 532226
rect 163082 532170 163138 532226
rect 163206 532170 163262 532226
rect 162834 532046 162890 532102
rect 162958 532046 163014 532102
rect 163082 532046 163138 532102
rect 163206 532046 163262 532102
rect 162834 531922 162890 531978
rect 162958 531922 163014 531978
rect 163082 531922 163138 531978
rect 163206 531922 163262 531978
rect 162834 514294 162890 514350
rect 162958 514294 163014 514350
rect 163082 514294 163138 514350
rect 163206 514294 163262 514350
rect 162834 514170 162890 514226
rect 162958 514170 163014 514226
rect 163082 514170 163138 514226
rect 163206 514170 163262 514226
rect 162834 514046 162890 514102
rect 162958 514046 163014 514102
rect 163082 514046 163138 514102
rect 163206 514046 163262 514102
rect 162834 513922 162890 513978
rect 162958 513922 163014 513978
rect 163082 513922 163138 513978
rect 163206 513922 163262 513978
rect 162834 496294 162890 496350
rect 162958 496294 163014 496350
rect 163082 496294 163138 496350
rect 163206 496294 163262 496350
rect 162834 496170 162890 496226
rect 162958 496170 163014 496226
rect 163082 496170 163138 496226
rect 163206 496170 163262 496226
rect 162834 496046 162890 496102
rect 162958 496046 163014 496102
rect 163082 496046 163138 496102
rect 163206 496046 163262 496102
rect 162834 495922 162890 495978
rect 162958 495922 163014 495978
rect 163082 495922 163138 495978
rect 163206 495922 163262 495978
rect 162834 478294 162890 478350
rect 162958 478294 163014 478350
rect 163082 478294 163138 478350
rect 163206 478294 163262 478350
rect 162834 478170 162890 478226
rect 162958 478170 163014 478226
rect 163082 478170 163138 478226
rect 163206 478170 163262 478226
rect 162834 478046 162890 478102
rect 162958 478046 163014 478102
rect 163082 478046 163138 478102
rect 163206 478046 163262 478102
rect 162834 477922 162890 477978
rect 162958 477922 163014 477978
rect 163082 477922 163138 477978
rect 163206 477922 163262 477978
rect 162834 460294 162890 460350
rect 162958 460294 163014 460350
rect 163082 460294 163138 460350
rect 163206 460294 163262 460350
rect 162834 460170 162890 460226
rect 162958 460170 163014 460226
rect 163082 460170 163138 460226
rect 163206 460170 163262 460226
rect 162834 460046 162890 460102
rect 162958 460046 163014 460102
rect 163082 460046 163138 460102
rect 163206 460046 163262 460102
rect 162834 459922 162890 459978
rect 162958 459922 163014 459978
rect 163082 459922 163138 459978
rect 163206 459922 163262 459978
rect 162834 442294 162890 442350
rect 162958 442294 163014 442350
rect 163082 442294 163138 442350
rect 163206 442294 163262 442350
rect 162834 442170 162890 442226
rect 162958 442170 163014 442226
rect 163082 442170 163138 442226
rect 163206 442170 163262 442226
rect 162834 442046 162890 442102
rect 162958 442046 163014 442102
rect 163082 442046 163138 442102
rect 163206 442046 163262 442102
rect 162834 441922 162890 441978
rect 162958 441922 163014 441978
rect 163082 441922 163138 441978
rect 163206 441922 163262 441978
rect 162834 424294 162890 424350
rect 162958 424294 163014 424350
rect 163082 424294 163138 424350
rect 163206 424294 163262 424350
rect 162834 424170 162890 424226
rect 162958 424170 163014 424226
rect 163082 424170 163138 424226
rect 163206 424170 163262 424226
rect 162834 424046 162890 424102
rect 162958 424046 163014 424102
rect 163082 424046 163138 424102
rect 163206 424046 163262 424102
rect 162834 423922 162890 423978
rect 162958 423922 163014 423978
rect 163082 423922 163138 423978
rect 163206 423922 163262 423978
rect 162834 406294 162890 406350
rect 162958 406294 163014 406350
rect 163082 406294 163138 406350
rect 163206 406294 163262 406350
rect 162834 406170 162890 406226
rect 162958 406170 163014 406226
rect 163082 406170 163138 406226
rect 163206 406170 163262 406226
rect 162834 406046 162890 406102
rect 162958 406046 163014 406102
rect 163082 406046 163138 406102
rect 163206 406046 163262 406102
rect 162834 405922 162890 405978
rect 162958 405922 163014 405978
rect 163082 405922 163138 405978
rect 163206 405922 163262 405978
rect 162834 388294 162890 388350
rect 162958 388294 163014 388350
rect 163082 388294 163138 388350
rect 163206 388294 163262 388350
rect 162834 388170 162890 388226
rect 162958 388170 163014 388226
rect 163082 388170 163138 388226
rect 163206 388170 163262 388226
rect 162834 388046 162890 388102
rect 162958 388046 163014 388102
rect 163082 388046 163138 388102
rect 163206 388046 163262 388102
rect 162834 387922 162890 387978
rect 162958 387922 163014 387978
rect 163082 387922 163138 387978
rect 163206 387922 163262 387978
rect 162834 370294 162890 370350
rect 162958 370294 163014 370350
rect 163082 370294 163138 370350
rect 163206 370294 163262 370350
rect 162834 370170 162890 370226
rect 162958 370170 163014 370226
rect 163082 370170 163138 370226
rect 163206 370170 163262 370226
rect 162834 370046 162890 370102
rect 162958 370046 163014 370102
rect 163082 370046 163138 370102
rect 163206 370046 163262 370102
rect 162834 369922 162890 369978
rect 162958 369922 163014 369978
rect 163082 369922 163138 369978
rect 163206 369922 163262 369978
rect 132114 352294 132170 352350
rect 132238 352294 132294 352350
rect 132362 352294 132418 352350
rect 132486 352294 132542 352350
rect 132114 352170 132170 352226
rect 132238 352170 132294 352226
rect 132362 352170 132418 352226
rect 132486 352170 132542 352226
rect 132114 352046 132170 352102
rect 132238 352046 132294 352102
rect 132362 352046 132418 352102
rect 132486 352046 132542 352102
rect 132114 351922 132170 351978
rect 132238 351922 132294 351978
rect 132362 351922 132418 351978
rect 132486 351922 132542 351978
rect 149878 352294 149934 352350
rect 150002 352294 150058 352350
rect 149878 352170 149934 352226
rect 150002 352170 150058 352226
rect 149878 352046 149934 352102
rect 150002 352046 150058 352102
rect 149878 351922 149934 351978
rect 150002 351922 150058 351978
rect 134518 346294 134574 346350
rect 134642 346294 134698 346350
rect 134518 346170 134574 346226
rect 134642 346170 134698 346226
rect 134518 346046 134574 346102
rect 134642 346046 134698 346102
rect 134518 345922 134574 345978
rect 134642 345922 134698 345978
rect 165238 346294 165294 346350
rect 165362 346294 165418 346350
rect 165238 346170 165294 346226
rect 165362 346170 165418 346226
rect 165238 346046 165294 346102
rect 165362 346046 165418 346102
rect 165238 345922 165294 345978
rect 165362 345922 165418 345978
rect 132114 334294 132170 334350
rect 132238 334294 132294 334350
rect 132362 334294 132418 334350
rect 132486 334294 132542 334350
rect 132114 334170 132170 334226
rect 132238 334170 132294 334226
rect 132362 334170 132418 334226
rect 132486 334170 132542 334226
rect 132114 334046 132170 334102
rect 132238 334046 132294 334102
rect 132362 334046 132418 334102
rect 132486 334046 132542 334102
rect 132114 333922 132170 333978
rect 132238 333922 132294 333978
rect 132362 333922 132418 333978
rect 132486 333922 132542 333978
rect 149878 334294 149934 334350
rect 150002 334294 150058 334350
rect 149878 334170 149934 334226
rect 150002 334170 150058 334226
rect 149878 334046 149934 334102
rect 150002 334046 150058 334102
rect 149878 333922 149934 333978
rect 150002 333922 150058 333978
rect 134518 328294 134574 328350
rect 134642 328294 134698 328350
rect 134518 328170 134574 328226
rect 134642 328170 134698 328226
rect 134518 328046 134574 328102
rect 134642 328046 134698 328102
rect 134518 327922 134574 327978
rect 134642 327922 134698 327978
rect 165238 328294 165294 328350
rect 165362 328294 165418 328350
rect 165238 328170 165294 328226
rect 165362 328170 165418 328226
rect 165238 328046 165294 328102
rect 165362 328046 165418 328102
rect 165238 327922 165294 327978
rect 165362 327922 165418 327978
rect 132114 316294 132170 316350
rect 132238 316294 132294 316350
rect 132362 316294 132418 316350
rect 132486 316294 132542 316350
rect 132114 316170 132170 316226
rect 132238 316170 132294 316226
rect 132362 316170 132418 316226
rect 132486 316170 132542 316226
rect 132114 316046 132170 316102
rect 132238 316046 132294 316102
rect 132362 316046 132418 316102
rect 132486 316046 132542 316102
rect 132114 315922 132170 315978
rect 132238 315922 132294 315978
rect 132362 315922 132418 315978
rect 132486 315922 132542 315978
rect 132114 298294 132170 298350
rect 132238 298294 132294 298350
rect 132362 298294 132418 298350
rect 132486 298294 132542 298350
rect 132114 298170 132170 298226
rect 132238 298170 132294 298226
rect 132362 298170 132418 298226
rect 132486 298170 132542 298226
rect 132114 298046 132170 298102
rect 132238 298046 132294 298102
rect 132362 298046 132418 298102
rect 132486 298046 132542 298102
rect 132114 297922 132170 297978
rect 132238 297922 132294 297978
rect 132362 297922 132418 297978
rect 132486 297922 132542 297978
rect 159114 310294 159170 310350
rect 159238 310294 159294 310350
rect 159362 310294 159418 310350
rect 159486 310294 159542 310350
rect 159114 310170 159170 310226
rect 159238 310170 159294 310226
rect 159362 310170 159418 310226
rect 159486 310170 159542 310226
rect 159114 310046 159170 310102
rect 159238 310046 159294 310102
rect 159362 310046 159418 310102
rect 159486 310046 159542 310102
rect 159114 309922 159170 309978
rect 159238 309922 159294 309978
rect 159362 309922 159418 309978
rect 159486 309922 159542 309978
rect 159114 292294 159170 292350
rect 159238 292294 159294 292350
rect 159362 292294 159418 292350
rect 159486 292294 159542 292350
rect 159114 292170 159170 292226
rect 159238 292170 159294 292226
rect 159362 292170 159418 292226
rect 159486 292170 159542 292226
rect 159114 292046 159170 292102
rect 159238 292046 159294 292102
rect 159362 292046 159418 292102
rect 159486 292046 159542 292102
rect 159114 291922 159170 291978
rect 159238 291922 159294 291978
rect 159362 291922 159418 291978
rect 159486 291922 159542 291978
rect 132114 280294 132170 280350
rect 132238 280294 132294 280350
rect 132362 280294 132418 280350
rect 132486 280294 132542 280350
rect 132114 280170 132170 280226
rect 132238 280170 132294 280226
rect 132362 280170 132418 280226
rect 132486 280170 132542 280226
rect 132114 280046 132170 280102
rect 132238 280046 132294 280102
rect 132362 280046 132418 280102
rect 132486 280046 132542 280102
rect 132114 279922 132170 279978
rect 132238 279922 132294 279978
rect 132362 279922 132418 279978
rect 132486 279922 132542 279978
rect 132114 262294 132170 262350
rect 132238 262294 132294 262350
rect 132362 262294 132418 262350
rect 132486 262294 132542 262350
rect 132114 262170 132170 262226
rect 132238 262170 132294 262226
rect 132362 262170 132418 262226
rect 132486 262170 132542 262226
rect 132114 262046 132170 262102
rect 132238 262046 132294 262102
rect 132362 262046 132418 262102
rect 132486 262046 132542 262102
rect 132114 261922 132170 261978
rect 132238 261922 132294 261978
rect 132362 261922 132418 261978
rect 132486 261922 132542 261978
rect 132114 244294 132170 244350
rect 132238 244294 132294 244350
rect 132362 244294 132418 244350
rect 132486 244294 132542 244350
rect 132114 244170 132170 244226
rect 132238 244170 132294 244226
rect 132362 244170 132418 244226
rect 132486 244170 132542 244226
rect 132114 244046 132170 244102
rect 132238 244046 132294 244102
rect 132362 244046 132418 244102
rect 132486 244046 132542 244102
rect 132114 243922 132170 243978
rect 132238 243922 132294 243978
rect 132362 243922 132418 243978
rect 132486 243922 132542 243978
rect 132114 226294 132170 226350
rect 132238 226294 132294 226350
rect 132362 226294 132418 226350
rect 132486 226294 132542 226350
rect 132114 226170 132170 226226
rect 132238 226170 132294 226226
rect 132362 226170 132418 226226
rect 132486 226170 132542 226226
rect 132114 226046 132170 226102
rect 132238 226046 132294 226102
rect 132362 226046 132418 226102
rect 132486 226046 132542 226102
rect 132114 225922 132170 225978
rect 132238 225922 132294 225978
rect 132362 225922 132418 225978
rect 132486 225922 132542 225978
rect 162834 316294 162890 316350
rect 162958 316294 163014 316350
rect 163082 316294 163138 316350
rect 163206 316294 163262 316350
rect 162834 316170 162890 316226
rect 162958 316170 163014 316226
rect 163082 316170 163138 316226
rect 163206 316170 163262 316226
rect 162834 316046 162890 316102
rect 162958 316046 163014 316102
rect 163082 316046 163138 316102
rect 163206 316046 163262 316102
rect 162834 315922 162890 315978
rect 162958 315922 163014 315978
rect 163082 315922 163138 315978
rect 163206 315922 163262 315978
rect 172172 322622 172228 322678
rect 162834 298294 162890 298350
rect 162958 298294 163014 298350
rect 163082 298294 163138 298350
rect 163206 298294 163262 298350
rect 162834 298170 162890 298226
rect 162958 298170 163014 298226
rect 163082 298170 163138 298226
rect 163206 298170 163262 298226
rect 162834 298046 162890 298102
rect 162958 298046 163014 298102
rect 163082 298046 163138 298102
rect 163206 298046 163262 298102
rect 162834 297922 162890 297978
rect 162958 297922 163014 297978
rect 163082 297922 163138 297978
rect 163206 297922 163262 297978
rect 147078 280294 147134 280350
rect 147202 280294 147258 280350
rect 147078 280170 147134 280226
rect 147202 280170 147258 280226
rect 147078 280046 147134 280102
rect 147202 280046 147258 280102
rect 147078 279922 147134 279978
rect 147202 279922 147258 279978
rect 152902 280294 152958 280350
rect 153026 280294 153082 280350
rect 152902 280170 152958 280226
rect 153026 280170 153082 280226
rect 152902 280046 152958 280102
rect 153026 280046 153082 280102
rect 152902 279922 152958 279978
rect 153026 279922 153082 279978
rect 158726 280294 158782 280350
rect 158850 280294 158906 280350
rect 158726 280170 158782 280226
rect 158850 280170 158906 280226
rect 158726 280046 158782 280102
rect 158850 280046 158906 280102
rect 158726 279922 158782 279978
rect 158850 279922 158906 279978
rect 164550 280294 164606 280350
rect 164674 280294 164730 280350
rect 164550 280170 164606 280226
rect 164674 280170 164730 280226
rect 164550 280046 164606 280102
rect 164674 280046 164730 280102
rect 164550 279922 164606 279978
rect 164674 279922 164730 279978
rect 144166 274294 144222 274350
rect 144290 274294 144346 274350
rect 144166 274170 144222 274226
rect 144290 274170 144346 274226
rect 144166 274046 144222 274102
rect 144290 274046 144346 274102
rect 144166 273922 144222 273978
rect 144290 273922 144346 273978
rect 149990 274294 150046 274350
rect 150114 274294 150170 274350
rect 149990 274170 150046 274226
rect 150114 274170 150170 274226
rect 149990 274046 150046 274102
rect 150114 274046 150170 274102
rect 149990 273922 150046 273978
rect 150114 273922 150170 273978
rect 155814 274294 155870 274350
rect 155938 274294 155994 274350
rect 155814 274170 155870 274226
rect 155938 274170 155994 274226
rect 155814 274046 155870 274102
rect 155938 274046 155994 274102
rect 155814 273922 155870 273978
rect 155938 273922 155994 273978
rect 161638 274294 161694 274350
rect 161762 274294 161818 274350
rect 161638 274170 161694 274226
rect 161762 274170 161818 274226
rect 161638 274046 161694 274102
rect 161762 274046 161818 274102
rect 161638 273922 161694 273978
rect 161762 273922 161818 273978
rect 162834 262294 162890 262350
rect 162958 262294 163014 262350
rect 163082 262294 163138 262350
rect 163206 262294 163262 262350
rect 162834 262170 162890 262226
rect 162958 262170 163014 262226
rect 163082 262170 163138 262226
rect 163206 262170 163262 262226
rect 162834 262046 162890 262102
rect 162958 262046 163014 262102
rect 163082 262046 163138 262102
rect 163206 262046 163262 262102
rect 162834 261922 162890 261978
rect 162958 261922 163014 261978
rect 163082 261922 163138 261978
rect 163206 261922 163262 261978
rect 159114 256294 159170 256350
rect 159238 256294 159294 256350
rect 159362 256294 159418 256350
rect 159486 256294 159542 256350
rect 159114 256170 159170 256226
rect 159238 256170 159294 256226
rect 159362 256170 159418 256226
rect 159486 256170 159542 256226
rect 159114 256046 159170 256102
rect 159238 256046 159294 256102
rect 159362 256046 159418 256102
rect 159486 256046 159542 256102
rect 159114 255922 159170 255978
rect 159238 255922 159294 255978
rect 159362 255922 159418 255978
rect 159486 255922 159542 255978
rect 159114 238294 159170 238350
rect 159238 238294 159294 238350
rect 159362 238294 159418 238350
rect 159486 238294 159542 238350
rect 159114 238170 159170 238226
rect 159238 238170 159294 238226
rect 159362 238170 159418 238226
rect 159486 238170 159542 238226
rect 159114 238046 159170 238102
rect 159238 238046 159294 238102
rect 159362 238046 159418 238102
rect 159486 238046 159542 238102
rect 159114 237922 159170 237978
rect 159238 237922 159294 237978
rect 159362 237922 159418 237978
rect 159486 237922 159542 237978
rect 159114 220294 159170 220350
rect 159238 220294 159294 220350
rect 159362 220294 159418 220350
rect 159486 220294 159542 220350
rect 159114 220170 159170 220226
rect 159238 220170 159294 220226
rect 159362 220170 159418 220226
rect 159486 220170 159542 220226
rect 159114 220046 159170 220102
rect 159238 220046 159294 220102
rect 159362 220046 159418 220102
rect 159486 220046 159542 220102
rect 159114 219922 159170 219978
rect 159238 219922 159294 219978
rect 159362 219922 159418 219978
rect 159486 219922 159542 219978
rect 162834 244294 162890 244350
rect 162958 244294 163014 244350
rect 163082 244294 163138 244350
rect 163206 244294 163262 244350
rect 162834 244170 162890 244226
rect 162958 244170 163014 244226
rect 163082 244170 163138 244226
rect 163206 244170 163262 244226
rect 162834 244046 162890 244102
rect 162958 244046 163014 244102
rect 163082 244046 163138 244102
rect 163206 244046 163262 244102
rect 162834 243922 162890 243978
rect 162958 243922 163014 243978
rect 163082 243922 163138 243978
rect 163206 243922 163262 243978
rect 162834 226294 162890 226350
rect 162958 226294 163014 226350
rect 163082 226294 163138 226350
rect 163206 226294 163262 226350
rect 162834 226170 162890 226226
rect 162958 226170 163014 226226
rect 163082 226170 163138 226226
rect 163206 226170 163262 226226
rect 162834 226046 162890 226102
rect 162958 226046 163014 226102
rect 163082 226046 163138 226102
rect 163206 226046 163262 226102
rect 162834 225922 162890 225978
rect 162958 225922 163014 225978
rect 163082 225922 163138 225978
rect 163206 225922 163262 225978
rect 170492 281402 170548 281458
rect 178108 340082 178164 340138
rect 184492 378782 184548 378838
rect 189834 562294 189890 562350
rect 189958 562294 190014 562350
rect 190082 562294 190138 562350
rect 190206 562294 190262 562350
rect 189834 562170 189890 562226
rect 189958 562170 190014 562226
rect 190082 562170 190138 562226
rect 190206 562170 190262 562226
rect 189834 562046 189890 562102
rect 189958 562046 190014 562102
rect 190082 562046 190138 562102
rect 190206 562046 190262 562102
rect 189834 561922 189890 561978
rect 189958 561922 190014 561978
rect 190082 561922 190138 561978
rect 190206 561922 190262 561978
rect 189834 544294 189890 544350
rect 189958 544294 190014 544350
rect 190082 544294 190138 544350
rect 190206 544294 190262 544350
rect 189834 544170 189890 544226
rect 189958 544170 190014 544226
rect 190082 544170 190138 544226
rect 190206 544170 190262 544226
rect 189834 544046 189890 544102
rect 189958 544046 190014 544102
rect 190082 544046 190138 544102
rect 190206 544046 190262 544102
rect 189834 543922 189890 543978
rect 189958 543922 190014 543978
rect 190082 543922 190138 543978
rect 190206 543922 190262 543978
rect 186172 403982 186228 404038
rect 185948 402362 186004 402418
rect 185500 211022 185556 211078
rect 189834 526294 189890 526350
rect 189958 526294 190014 526350
rect 190082 526294 190138 526350
rect 190206 526294 190262 526350
rect 189834 526170 189890 526226
rect 189958 526170 190014 526226
rect 190082 526170 190138 526226
rect 190206 526170 190262 526226
rect 189834 526046 189890 526102
rect 189958 526046 190014 526102
rect 190082 526046 190138 526102
rect 190206 526046 190262 526102
rect 189834 525922 189890 525978
rect 189958 525922 190014 525978
rect 190082 525922 190138 525978
rect 190206 525922 190262 525978
rect 189834 508294 189890 508350
rect 189958 508294 190014 508350
rect 190082 508294 190138 508350
rect 190206 508294 190262 508350
rect 189834 508170 189890 508226
rect 189958 508170 190014 508226
rect 190082 508170 190138 508226
rect 190206 508170 190262 508226
rect 189834 508046 189890 508102
rect 189958 508046 190014 508102
rect 190082 508046 190138 508102
rect 190206 508046 190262 508102
rect 189834 507922 189890 507978
rect 189958 507922 190014 507978
rect 190082 507922 190138 507978
rect 190206 507922 190262 507978
rect 189834 490294 189890 490350
rect 189958 490294 190014 490350
rect 190082 490294 190138 490350
rect 190206 490294 190262 490350
rect 189834 490170 189890 490226
rect 189958 490170 190014 490226
rect 190082 490170 190138 490226
rect 190206 490170 190262 490226
rect 189834 490046 189890 490102
rect 189958 490046 190014 490102
rect 190082 490046 190138 490102
rect 190206 490046 190262 490102
rect 189834 489922 189890 489978
rect 189958 489922 190014 489978
rect 190082 489922 190138 489978
rect 190206 489922 190262 489978
rect 186396 268802 186452 268858
rect 187404 322622 187460 322678
rect 187292 288962 187348 289018
rect 187180 287162 187236 287218
rect 189834 472294 189890 472350
rect 189958 472294 190014 472350
rect 190082 472294 190138 472350
rect 190206 472294 190262 472350
rect 189834 472170 189890 472226
rect 189958 472170 190014 472226
rect 190082 472170 190138 472226
rect 190206 472170 190262 472226
rect 189834 472046 189890 472102
rect 189958 472046 190014 472102
rect 190082 472046 190138 472102
rect 190206 472046 190262 472102
rect 189834 471922 189890 471978
rect 189958 471922 190014 471978
rect 190082 471922 190138 471978
rect 190206 471922 190262 471978
rect 189834 454294 189890 454350
rect 189958 454294 190014 454350
rect 190082 454294 190138 454350
rect 190206 454294 190262 454350
rect 189834 454170 189890 454226
rect 189958 454170 190014 454226
rect 190082 454170 190138 454226
rect 190206 454170 190262 454226
rect 189834 454046 189890 454102
rect 189958 454046 190014 454102
rect 190082 454046 190138 454102
rect 190206 454046 190262 454102
rect 189834 453922 189890 453978
rect 189958 453922 190014 453978
rect 190082 453922 190138 453978
rect 190206 453922 190262 453978
rect 189834 436294 189890 436350
rect 189958 436294 190014 436350
rect 190082 436294 190138 436350
rect 190206 436294 190262 436350
rect 189834 436170 189890 436226
rect 189958 436170 190014 436226
rect 190082 436170 190138 436226
rect 190206 436170 190262 436226
rect 189834 436046 189890 436102
rect 189958 436046 190014 436102
rect 190082 436046 190138 436102
rect 190206 436046 190262 436102
rect 189834 435922 189890 435978
rect 189958 435922 190014 435978
rect 190082 435922 190138 435978
rect 190206 435922 190262 435978
rect 190652 421820 190708 421858
rect 190652 421802 190708 421820
rect 192332 421802 192388 421858
rect 189834 418294 189890 418350
rect 189958 418294 190014 418350
rect 190082 418294 190138 418350
rect 190206 418294 190262 418350
rect 189834 418170 189890 418226
rect 189958 418170 190014 418226
rect 190082 418170 190138 418226
rect 190206 418170 190262 418226
rect 189834 418046 189890 418102
rect 189958 418046 190014 418102
rect 190082 418046 190138 418102
rect 190206 418046 190262 418102
rect 189834 417922 189890 417978
rect 189958 417922 190014 417978
rect 190082 417922 190138 417978
rect 190206 417922 190262 417978
rect 189834 400294 189890 400350
rect 189958 400294 190014 400350
rect 190082 400294 190138 400350
rect 190206 400294 190262 400350
rect 189834 400170 189890 400226
rect 189958 400170 190014 400226
rect 190082 400170 190138 400226
rect 190206 400170 190262 400226
rect 189834 400046 189890 400102
rect 189958 400046 190014 400102
rect 190082 400046 190138 400102
rect 190206 400046 190262 400102
rect 189834 399922 189890 399978
rect 189958 399922 190014 399978
rect 190082 399922 190138 399978
rect 190206 399922 190262 399978
rect 189834 382294 189890 382350
rect 189958 382294 190014 382350
rect 190082 382294 190138 382350
rect 190206 382294 190262 382350
rect 189834 382170 189890 382226
rect 189958 382170 190014 382226
rect 190082 382170 190138 382226
rect 190206 382170 190262 382226
rect 189834 382046 189890 382102
rect 189958 382046 190014 382102
rect 190082 382046 190138 382102
rect 190206 382046 190262 382102
rect 189834 381922 189890 381978
rect 189958 381922 190014 381978
rect 190082 381922 190138 381978
rect 190206 381922 190262 381978
rect 220554 597156 220610 597212
rect 220678 597156 220734 597212
rect 220802 597156 220858 597212
rect 220926 597156 220982 597212
rect 220554 597032 220610 597088
rect 220678 597032 220734 597088
rect 220802 597032 220858 597088
rect 220926 597032 220982 597088
rect 220554 596908 220610 596964
rect 220678 596908 220734 596964
rect 220802 596908 220858 596964
rect 220926 596908 220982 596964
rect 220554 596784 220610 596840
rect 220678 596784 220734 596840
rect 220802 596784 220858 596840
rect 220926 596784 220982 596840
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 193554 406294 193610 406350
rect 193678 406294 193734 406350
rect 193802 406294 193858 406350
rect 193926 406294 193982 406350
rect 193554 406170 193610 406226
rect 193678 406170 193734 406226
rect 193802 406170 193858 406226
rect 193926 406170 193982 406226
rect 193554 406046 193610 406102
rect 193678 406046 193734 406102
rect 193802 406046 193858 406102
rect 193926 406046 193982 406102
rect 193554 405922 193610 405978
rect 193678 405922 193734 405978
rect 193802 405922 193858 405978
rect 193926 405922 193982 405978
rect 220554 580294 220610 580350
rect 220678 580294 220734 580350
rect 220802 580294 220858 580350
rect 220926 580294 220982 580350
rect 220554 580170 220610 580226
rect 220678 580170 220734 580226
rect 220802 580170 220858 580226
rect 220926 580170 220982 580226
rect 220554 580046 220610 580102
rect 220678 580046 220734 580102
rect 220802 580046 220858 580102
rect 220926 580046 220982 580102
rect 220554 579922 220610 579978
rect 220678 579922 220734 579978
rect 220802 579922 220858 579978
rect 220926 579922 220982 579978
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 251274 597156 251330 597212
rect 251398 597156 251454 597212
rect 251522 597156 251578 597212
rect 251646 597156 251702 597212
rect 251274 597032 251330 597088
rect 251398 597032 251454 597088
rect 251522 597032 251578 597088
rect 251646 597032 251702 597088
rect 251274 596908 251330 596964
rect 251398 596908 251454 596964
rect 251522 596908 251578 596964
rect 251646 596908 251702 596964
rect 251274 596784 251330 596840
rect 251398 596784 251454 596840
rect 251522 596784 251578 596840
rect 251646 596784 251702 596840
rect 251274 580294 251330 580350
rect 251398 580294 251454 580350
rect 251522 580294 251578 580350
rect 251646 580294 251702 580350
rect 251274 580170 251330 580226
rect 251398 580170 251454 580226
rect 251522 580170 251578 580226
rect 251646 580170 251702 580226
rect 251274 580046 251330 580102
rect 251398 580046 251454 580102
rect 251522 580046 251578 580102
rect 251646 580046 251702 580102
rect 251274 579922 251330 579978
rect 251398 579922 251454 579978
rect 251522 579922 251578 579978
rect 251646 579922 251702 579978
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 281994 597156 282050 597212
rect 282118 597156 282174 597212
rect 282242 597156 282298 597212
rect 282366 597156 282422 597212
rect 281994 597032 282050 597088
rect 282118 597032 282174 597088
rect 282242 597032 282298 597088
rect 282366 597032 282422 597088
rect 281994 596908 282050 596964
rect 282118 596908 282174 596964
rect 282242 596908 282298 596964
rect 282366 596908 282422 596964
rect 281994 596784 282050 596840
rect 282118 596784 282174 596840
rect 282242 596784 282298 596840
rect 282366 596784 282422 596840
rect 281994 580294 282050 580350
rect 282118 580294 282174 580350
rect 282242 580294 282298 580350
rect 282366 580294 282422 580350
rect 281994 580170 282050 580226
rect 282118 580170 282174 580226
rect 282242 580170 282298 580226
rect 282366 580170 282422 580226
rect 281994 580046 282050 580102
rect 282118 580046 282174 580102
rect 282242 580046 282298 580102
rect 282366 580046 282422 580102
rect 281994 579922 282050 579978
rect 282118 579922 282174 579978
rect 282242 579922 282298 579978
rect 282366 579922 282422 579978
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 312714 597156 312770 597212
rect 312838 597156 312894 597212
rect 312962 597156 313018 597212
rect 313086 597156 313142 597212
rect 312714 597032 312770 597088
rect 312838 597032 312894 597088
rect 312962 597032 313018 597088
rect 313086 597032 313142 597088
rect 312714 596908 312770 596964
rect 312838 596908 312894 596964
rect 312962 596908 313018 596964
rect 313086 596908 313142 596964
rect 312714 596784 312770 596840
rect 312838 596784 312894 596840
rect 312962 596784 313018 596840
rect 313086 596784 313142 596840
rect 312714 580294 312770 580350
rect 312838 580294 312894 580350
rect 312962 580294 313018 580350
rect 313086 580294 313142 580350
rect 312714 580170 312770 580226
rect 312838 580170 312894 580226
rect 312962 580170 313018 580226
rect 313086 580170 313142 580226
rect 312714 580046 312770 580102
rect 312838 580046 312894 580102
rect 312962 580046 313018 580102
rect 313086 580046 313142 580102
rect 312714 579922 312770 579978
rect 312838 579922 312894 579978
rect 312962 579922 313018 579978
rect 313086 579922 313142 579978
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 343434 597156 343490 597212
rect 343558 597156 343614 597212
rect 343682 597156 343738 597212
rect 343806 597156 343862 597212
rect 343434 597032 343490 597088
rect 343558 597032 343614 597088
rect 343682 597032 343738 597088
rect 343806 597032 343862 597088
rect 343434 596908 343490 596964
rect 343558 596908 343614 596964
rect 343682 596908 343738 596964
rect 343806 596908 343862 596964
rect 343434 596784 343490 596840
rect 343558 596784 343614 596840
rect 343682 596784 343738 596840
rect 343806 596784 343862 596840
rect 343434 580294 343490 580350
rect 343558 580294 343614 580350
rect 343682 580294 343738 580350
rect 343806 580294 343862 580350
rect 343434 580170 343490 580226
rect 343558 580170 343614 580226
rect 343682 580170 343738 580226
rect 343806 580170 343862 580226
rect 343434 580046 343490 580102
rect 343558 580046 343614 580102
rect 343682 580046 343738 580102
rect 343806 580046 343862 580102
rect 343434 579922 343490 579978
rect 343558 579922 343614 579978
rect 343682 579922 343738 579978
rect 343806 579922 343862 579978
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 374154 597156 374210 597212
rect 374278 597156 374334 597212
rect 374402 597156 374458 597212
rect 374526 597156 374582 597212
rect 374154 597032 374210 597088
rect 374278 597032 374334 597088
rect 374402 597032 374458 597088
rect 374526 597032 374582 597088
rect 374154 596908 374210 596964
rect 374278 596908 374334 596964
rect 374402 596908 374458 596964
rect 374526 596908 374582 596964
rect 374154 596784 374210 596840
rect 374278 596784 374334 596840
rect 374402 596784 374458 596840
rect 374526 596784 374582 596840
rect 374154 580294 374210 580350
rect 374278 580294 374334 580350
rect 374402 580294 374458 580350
rect 374526 580294 374582 580350
rect 374154 580170 374210 580226
rect 374278 580170 374334 580226
rect 374402 580170 374458 580226
rect 374526 580170 374582 580226
rect 374154 580046 374210 580102
rect 374278 580046 374334 580102
rect 374402 580046 374458 580102
rect 374526 580046 374582 580102
rect 374154 579922 374210 579978
rect 374278 579922 374334 579978
rect 374402 579922 374458 579978
rect 374526 579922 374582 579978
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 404874 597156 404930 597212
rect 404998 597156 405054 597212
rect 405122 597156 405178 597212
rect 405246 597156 405302 597212
rect 404874 597032 404930 597088
rect 404998 597032 405054 597088
rect 405122 597032 405178 597088
rect 405246 597032 405302 597088
rect 404874 596908 404930 596964
rect 404998 596908 405054 596964
rect 405122 596908 405178 596964
rect 405246 596908 405302 596964
rect 404874 596784 404930 596840
rect 404998 596784 405054 596840
rect 405122 596784 405178 596840
rect 405246 596784 405302 596840
rect 404874 580294 404930 580350
rect 404998 580294 405054 580350
rect 405122 580294 405178 580350
rect 405246 580294 405302 580350
rect 404874 580170 404930 580226
rect 404998 580170 405054 580226
rect 405122 580170 405178 580226
rect 405246 580170 405302 580226
rect 404874 580046 404930 580102
rect 404998 580046 405054 580102
rect 405122 580046 405178 580102
rect 405246 580046 405302 580102
rect 404874 579922 404930 579978
rect 404998 579922 405054 579978
rect 405122 579922 405178 579978
rect 405246 579922 405302 579978
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 435594 597156 435650 597212
rect 435718 597156 435774 597212
rect 435842 597156 435898 597212
rect 435966 597156 436022 597212
rect 435594 597032 435650 597088
rect 435718 597032 435774 597088
rect 435842 597032 435898 597088
rect 435966 597032 436022 597088
rect 435594 596908 435650 596964
rect 435718 596908 435774 596964
rect 435842 596908 435898 596964
rect 435966 596908 436022 596964
rect 435594 596784 435650 596840
rect 435718 596784 435774 596840
rect 435842 596784 435898 596840
rect 435966 596784 436022 596840
rect 435594 580294 435650 580350
rect 435718 580294 435774 580350
rect 435842 580294 435898 580350
rect 435966 580294 436022 580350
rect 435594 580170 435650 580226
rect 435718 580170 435774 580226
rect 435842 580170 435898 580226
rect 435966 580170 436022 580226
rect 435594 580046 435650 580102
rect 435718 580046 435774 580102
rect 435842 580046 435898 580102
rect 435966 580046 436022 580102
rect 435594 579922 435650 579978
rect 435718 579922 435774 579978
rect 435842 579922 435898 579978
rect 435966 579922 436022 579978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 466314 597156 466370 597212
rect 466438 597156 466494 597212
rect 466562 597156 466618 597212
rect 466686 597156 466742 597212
rect 466314 597032 466370 597088
rect 466438 597032 466494 597088
rect 466562 597032 466618 597088
rect 466686 597032 466742 597088
rect 466314 596908 466370 596964
rect 466438 596908 466494 596964
rect 466562 596908 466618 596964
rect 466686 596908 466742 596964
rect 466314 596784 466370 596840
rect 466438 596784 466494 596840
rect 466562 596784 466618 596840
rect 466686 596784 466742 596840
rect 466314 580294 466370 580350
rect 466438 580294 466494 580350
rect 466562 580294 466618 580350
rect 466686 580294 466742 580350
rect 466314 580170 466370 580226
rect 466438 580170 466494 580226
rect 466562 580170 466618 580226
rect 466686 580170 466742 580226
rect 466314 580046 466370 580102
rect 466438 580046 466494 580102
rect 466562 580046 466618 580102
rect 466686 580046 466742 580102
rect 466314 579922 466370 579978
rect 466438 579922 466494 579978
rect 466562 579922 466618 579978
rect 466686 579922 466742 579978
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 497034 597156 497090 597212
rect 497158 597156 497214 597212
rect 497282 597156 497338 597212
rect 497406 597156 497462 597212
rect 497034 597032 497090 597088
rect 497158 597032 497214 597088
rect 497282 597032 497338 597088
rect 497406 597032 497462 597088
rect 497034 596908 497090 596964
rect 497158 596908 497214 596964
rect 497282 596908 497338 596964
rect 497406 596908 497462 596964
rect 497034 596784 497090 596840
rect 497158 596784 497214 596840
rect 497282 596784 497338 596840
rect 497406 596784 497462 596840
rect 497034 580294 497090 580350
rect 497158 580294 497214 580350
rect 497282 580294 497338 580350
rect 497406 580294 497462 580350
rect 497034 580170 497090 580226
rect 497158 580170 497214 580226
rect 497282 580170 497338 580226
rect 497406 580170 497462 580226
rect 497034 580046 497090 580102
rect 497158 580046 497214 580102
rect 497282 580046 497338 580102
rect 497406 580046 497462 580102
rect 497034 579922 497090 579978
rect 497158 579922 497214 579978
rect 497282 579922 497338 579978
rect 497406 579922 497462 579978
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 527754 597156 527810 597212
rect 527878 597156 527934 597212
rect 528002 597156 528058 597212
rect 528126 597156 528182 597212
rect 527754 597032 527810 597088
rect 527878 597032 527934 597088
rect 528002 597032 528058 597088
rect 528126 597032 528182 597088
rect 527754 596908 527810 596964
rect 527878 596908 527934 596964
rect 528002 596908 528058 596964
rect 528126 596908 528182 596964
rect 527754 596784 527810 596840
rect 527878 596784 527934 596840
rect 528002 596784 528058 596840
rect 528126 596784 528182 596840
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 194518 562294 194574 562350
rect 194642 562294 194698 562350
rect 194518 562170 194574 562226
rect 194642 562170 194698 562226
rect 194518 562046 194574 562102
rect 194642 562046 194698 562102
rect 194518 561922 194574 561978
rect 194642 561922 194698 561978
rect 225238 562294 225294 562350
rect 225362 562294 225418 562350
rect 225238 562170 225294 562226
rect 225362 562170 225418 562226
rect 225238 562046 225294 562102
rect 225362 562046 225418 562102
rect 225238 561922 225294 561978
rect 225362 561922 225418 561978
rect 255958 562294 256014 562350
rect 256082 562294 256138 562350
rect 255958 562170 256014 562226
rect 256082 562170 256138 562226
rect 255958 562046 256014 562102
rect 256082 562046 256138 562102
rect 255958 561922 256014 561978
rect 256082 561922 256138 561978
rect 286678 562294 286734 562350
rect 286802 562294 286858 562350
rect 286678 562170 286734 562226
rect 286802 562170 286858 562226
rect 286678 562046 286734 562102
rect 286802 562046 286858 562102
rect 286678 561922 286734 561978
rect 286802 561922 286858 561978
rect 317398 562294 317454 562350
rect 317522 562294 317578 562350
rect 317398 562170 317454 562226
rect 317522 562170 317578 562226
rect 317398 562046 317454 562102
rect 317522 562046 317578 562102
rect 317398 561922 317454 561978
rect 317522 561922 317578 561978
rect 348118 562294 348174 562350
rect 348242 562294 348298 562350
rect 348118 562170 348174 562226
rect 348242 562170 348298 562226
rect 348118 562046 348174 562102
rect 348242 562046 348298 562102
rect 348118 561922 348174 561978
rect 348242 561922 348298 561978
rect 378838 562294 378894 562350
rect 378962 562294 379018 562350
rect 378838 562170 378894 562226
rect 378962 562170 379018 562226
rect 378838 562046 378894 562102
rect 378962 562046 379018 562102
rect 378838 561922 378894 561978
rect 378962 561922 379018 561978
rect 409558 562294 409614 562350
rect 409682 562294 409738 562350
rect 409558 562170 409614 562226
rect 409682 562170 409738 562226
rect 409558 562046 409614 562102
rect 409682 562046 409738 562102
rect 409558 561922 409614 561978
rect 409682 561922 409738 561978
rect 440278 562294 440334 562350
rect 440402 562294 440458 562350
rect 440278 562170 440334 562226
rect 440402 562170 440458 562226
rect 440278 562046 440334 562102
rect 440402 562046 440458 562102
rect 440278 561922 440334 561978
rect 440402 561922 440458 561978
rect 470998 562294 471054 562350
rect 471122 562294 471178 562350
rect 470998 562170 471054 562226
rect 471122 562170 471178 562226
rect 470998 562046 471054 562102
rect 471122 562046 471178 562102
rect 470998 561922 471054 561978
rect 471122 561922 471178 561978
rect 501718 562294 501774 562350
rect 501842 562294 501898 562350
rect 501718 562170 501774 562226
rect 501842 562170 501898 562226
rect 501718 562046 501774 562102
rect 501842 562046 501898 562102
rect 501718 561922 501774 561978
rect 501842 561922 501898 561978
rect 209878 550294 209934 550350
rect 210002 550294 210058 550350
rect 209878 550170 209934 550226
rect 210002 550170 210058 550226
rect 209878 550046 209934 550102
rect 210002 550046 210058 550102
rect 209878 549922 209934 549978
rect 210002 549922 210058 549978
rect 240598 550294 240654 550350
rect 240722 550294 240778 550350
rect 240598 550170 240654 550226
rect 240722 550170 240778 550226
rect 240598 550046 240654 550102
rect 240722 550046 240778 550102
rect 240598 549922 240654 549978
rect 240722 549922 240778 549978
rect 271318 550294 271374 550350
rect 271442 550294 271498 550350
rect 271318 550170 271374 550226
rect 271442 550170 271498 550226
rect 271318 550046 271374 550102
rect 271442 550046 271498 550102
rect 271318 549922 271374 549978
rect 271442 549922 271498 549978
rect 302038 550294 302094 550350
rect 302162 550294 302218 550350
rect 302038 550170 302094 550226
rect 302162 550170 302218 550226
rect 302038 550046 302094 550102
rect 302162 550046 302218 550102
rect 302038 549922 302094 549978
rect 302162 549922 302218 549978
rect 332758 550294 332814 550350
rect 332882 550294 332938 550350
rect 332758 550170 332814 550226
rect 332882 550170 332938 550226
rect 332758 550046 332814 550102
rect 332882 550046 332938 550102
rect 332758 549922 332814 549978
rect 332882 549922 332938 549978
rect 363478 550294 363534 550350
rect 363602 550294 363658 550350
rect 363478 550170 363534 550226
rect 363602 550170 363658 550226
rect 363478 550046 363534 550102
rect 363602 550046 363658 550102
rect 363478 549922 363534 549978
rect 363602 549922 363658 549978
rect 394198 550294 394254 550350
rect 394322 550294 394378 550350
rect 394198 550170 394254 550226
rect 394322 550170 394378 550226
rect 394198 550046 394254 550102
rect 394322 550046 394378 550102
rect 394198 549922 394254 549978
rect 394322 549922 394378 549978
rect 424918 550294 424974 550350
rect 425042 550294 425098 550350
rect 424918 550170 424974 550226
rect 425042 550170 425098 550226
rect 424918 550046 424974 550102
rect 425042 550046 425098 550102
rect 424918 549922 424974 549978
rect 425042 549922 425098 549978
rect 455638 550294 455694 550350
rect 455762 550294 455818 550350
rect 455638 550170 455694 550226
rect 455762 550170 455818 550226
rect 455638 550046 455694 550102
rect 455762 550046 455818 550102
rect 455638 549922 455694 549978
rect 455762 549922 455818 549978
rect 486358 550294 486414 550350
rect 486482 550294 486538 550350
rect 486358 550170 486414 550226
rect 486482 550170 486538 550226
rect 486358 550046 486414 550102
rect 486482 550046 486538 550102
rect 486358 549922 486414 549978
rect 486482 549922 486538 549978
rect 194518 544294 194574 544350
rect 194642 544294 194698 544350
rect 194518 544170 194574 544226
rect 194642 544170 194698 544226
rect 194518 544046 194574 544102
rect 194642 544046 194698 544102
rect 194518 543922 194574 543978
rect 194642 543922 194698 543978
rect 225238 544294 225294 544350
rect 225362 544294 225418 544350
rect 225238 544170 225294 544226
rect 225362 544170 225418 544226
rect 225238 544046 225294 544102
rect 225362 544046 225418 544102
rect 225238 543922 225294 543978
rect 225362 543922 225418 543978
rect 255958 544294 256014 544350
rect 256082 544294 256138 544350
rect 255958 544170 256014 544226
rect 256082 544170 256138 544226
rect 255958 544046 256014 544102
rect 256082 544046 256138 544102
rect 255958 543922 256014 543978
rect 256082 543922 256138 543978
rect 286678 544294 286734 544350
rect 286802 544294 286858 544350
rect 286678 544170 286734 544226
rect 286802 544170 286858 544226
rect 286678 544046 286734 544102
rect 286802 544046 286858 544102
rect 286678 543922 286734 543978
rect 286802 543922 286858 543978
rect 317398 544294 317454 544350
rect 317522 544294 317578 544350
rect 317398 544170 317454 544226
rect 317522 544170 317578 544226
rect 317398 544046 317454 544102
rect 317522 544046 317578 544102
rect 317398 543922 317454 543978
rect 317522 543922 317578 543978
rect 348118 544294 348174 544350
rect 348242 544294 348298 544350
rect 348118 544170 348174 544226
rect 348242 544170 348298 544226
rect 348118 544046 348174 544102
rect 348242 544046 348298 544102
rect 348118 543922 348174 543978
rect 348242 543922 348298 543978
rect 378838 544294 378894 544350
rect 378962 544294 379018 544350
rect 378838 544170 378894 544226
rect 378962 544170 379018 544226
rect 378838 544046 378894 544102
rect 378962 544046 379018 544102
rect 378838 543922 378894 543978
rect 378962 543922 379018 543978
rect 409558 544294 409614 544350
rect 409682 544294 409738 544350
rect 409558 544170 409614 544226
rect 409682 544170 409738 544226
rect 409558 544046 409614 544102
rect 409682 544046 409738 544102
rect 409558 543922 409614 543978
rect 409682 543922 409738 543978
rect 440278 544294 440334 544350
rect 440402 544294 440458 544350
rect 440278 544170 440334 544226
rect 440402 544170 440458 544226
rect 440278 544046 440334 544102
rect 440402 544046 440458 544102
rect 440278 543922 440334 543978
rect 440402 543922 440458 543978
rect 470998 544294 471054 544350
rect 471122 544294 471178 544350
rect 470998 544170 471054 544226
rect 471122 544170 471178 544226
rect 470998 544046 471054 544102
rect 471122 544046 471178 544102
rect 470998 543922 471054 543978
rect 471122 543922 471178 543978
rect 501718 544294 501774 544350
rect 501842 544294 501898 544350
rect 501718 544170 501774 544226
rect 501842 544170 501898 544226
rect 501718 544046 501774 544102
rect 501842 544046 501898 544102
rect 501718 543922 501774 543978
rect 501842 543922 501898 543978
rect 209878 532294 209934 532350
rect 210002 532294 210058 532350
rect 209878 532170 209934 532226
rect 210002 532170 210058 532226
rect 209878 532046 209934 532102
rect 210002 532046 210058 532102
rect 209878 531922 209934 531978
rect 210002 531922 210058 531978
rect 240598 532294 240654 532350
rect 240722 532294 240778 532350
rect 240598 532170 240654 532226
rect 240722 532170 240778 532226
rect 240598 532046 240654 532102
rect 240722 532046 240778 532102
rect 240598 531922 240654 531978
rect 240722 531922 240778 531978
rect 271318 532294 271374 532350
rect 271442 532294 271498 532350
rect 271318 532170 271374 532226
rect 271442 532170 271498 532226
rect 271318 532046 271374 532102
rect 271442 532046 271498 532102
rect 271318 531922 271374 531978
rect 271442 531922 271498 531978
rect 302038 532294 302094 532350
rect 302162 532294 302218 532350
rect 302038 532170 302094 532226
rect 302162 532170 302218 532226
rect 302038 532046 302094 532102
rect 302162 532046 302218 532102
rect 302038 531922 302094 531978
rect 302162 531922 302218 531978
rect 332758 532294 332814 532350
rect 332882 532294 332938 532350
rect 332758 532170 332814 532226
rect 332882 532170 332938 532226
rect 332758 532046 332814 532102
rect 332882 532046 332938 532102
rect 332758 531922 332814 531978
rect 332882 531922 332938 531978
rect 363478 532294 363534 532350
rect 363602 532294 363658 532350
rect 363478 532170 363534 532226
rect 363602 532170 363658 532226
rect 363478 532046 363534 532102
rect 363602 532046 363658 532102
rect 363478 531922 363534 531978
rect 363602 531922 363658 531978
rect 394198 532294 394254 532350
rect 394322 532294 394378 532350
rect 394198 532170 394254 532226
rect 394322 532170 394378 532226
rect 394198 532046 394254 532102
rect 394322 532046 394378 532102
rect 394198 531922 394254 531978
rect 394322 531922 394378 531978
rect 424918 532294 424974 532350
rect 425042 532294 425098 532350
rect 424918 532170 424974 532226
rect 425042 532170 425098 532226
rect 424918 532046 424974 532102
rect 425042 532046 425098 532102
rect 424918 531922 424974 531978
rect 425042 531922 425098 531978
rect 455638 532294 455694 532350
rect 455762 532294 455818 532350
rect 455638 532170 455694 532226
rect 455762 532170 455818 532226
rect 455638 532046 455694 532102
rect 455762 532046 455818 532102
rect 455638 531922 455694 531978
rect 455762 531922 455818 531978
rect 486358 532294 486414 532350
rect 486482 532294 486538 532350
rect 486358 532170 486414 532226
rect 486482 532170 486538 532226
rect 486358 532046 486414 532102
rect 486482 532046 486538 532102
rect 486358 531922 486414 531978
rect 486482 531922 486538 531978
rect 194518 526294 194574 526350
rect 194642 526294 194698 526350
rect 194518 526170 194574 526226
rect 194642 526170 194698 526226
rect 194518 526046 194574 526102
rect 194642 526046 194698 526102
rect 194518 525922 194574 525978
rect 194642 525922 194698 525978
rect 225238 526294 225294 526350
rect 225362 526294 225418 526350
rect 225238 526170 225294 526226
rect 225362 526170 225418 526226
rect 225238 526046 225294 526102
rect 225362 526046 225418 526102
rect 225238 525922 225294 525978
rect 225362 525922 225418 525978
rect 255958 526294 256014 526350
rect 256082 526294 256138 526350
rect 255958 526170 256014 526226
rect 256082 526170 256138 526226
rect 255958 526046 256014 526102
rect 256082 526046 256138 526102
rect 255958 525922 256014 525978
rect 256082 525922 256138 525978
rect 286678 526294 286734 526350
rect 286802 526294 286858 526350
rect 286678 526170 286734 526226
rect 286802 526170 286858 526226
rect 286678 526046 286734 526102
rect 286802 526046 286858 526102
rect 286678 525922 286734 525978
rect 286802 525922 286858 525978
rect 317398 526294 317454 526350
rect 317522 526294 317578 526350
rect 317398 526170 317454 526226
rect 317522 526170 317578 526226
rect 317398 526046 317454 526102
rect 317522 526046 317578 526102
rect 317398 525922 317454 525978
rect 317522 525922 317578 525978
rect 348118 526294 348174 526350
rect 348242 526294 348298 526350
rect 348118 526170 348174 526226
rect 348242 526170 348298 526226
rect 348118 526046 348174 526102
rect 348242 526046 348298 526102
rect 348118 525922 348174 525978
rect 348242 525922 348298 525978
rect 378838 526294 378894 526350
rect 378962 526294 379018 526350
rect 378838 526170 378894 526226
rect 378962 526170 379018 526226
rect 378838 526046 378894 526102
rect 378962 526046 379018 526102
rect 378838 525922 378894 525978
rect 378962 525922 379018 525978
rect 409558 526294 409614 526350
rect 409682 526294 409738 526350
rect 409558 526170 409614 526226
rect 409682 526170 409738 526226
rect 409558 526046 409614 526102
rect 409682 526046 409738 526102
rect 409558 525922 409614 525978
rect 409682 525922 409738 525978
rect 440278 526294 440334 526350
rect 440402 526294 440458 526350
rect 440278 526170 440334 526226
rect 440402 526170 440458 526226
rect 440278 526046 440334 526102
rect 440402 526046 440458 526102
rect 440278 525922 440334 525978
rect 440402 525922 440458 525978
rect 470998 526294 471054 526350
rect 471122 526294 471178 526350
rect 470998 526170 471054 526226
rect 471122 526170 471178 526226
rect 470998 526046 471054 526102
rect 471122 526046 471178 526102
rect 470998 525922 471054 525978
rect 471122 525922 471178 525978
rect 501718 526294 501774 526350
rect 501842 526294 501898 526350
rect 501718 526170 501774 526226
rect 501842 526170 501898 526226
rect 501718 526046 501774 526102
rect 501842 526046 501898 526102
rect 501718 525922 501774 525978
rect 501842 525922 501898 525978
rect 209878 514294 209934 514350
rect 210002 514294 210058 514350
rect 209878 514170 209934 514226
rect 210002 514170 210058 514226
rect 209878 514046 209934 514102
rect 210002 514046 210058 514102
rect 209878 513922 209934 513978
rect 210002 513922 210058 513978
rect 240598 514294 240654 514350
rect 240722 514294 240778 514350
rect 240598 514170 240654 514226
rect 240722 514170 240778 514226
rect 240598 514046 240654 514102
rect 240722 514046 240778 514102
rect 240598 513922 240654 513978
rect 240722 513922 240778 513978
rect 271318 514294 271374 514350
rect 271442 514294 271498 514350
rect 271318 514170 271374 514226
rect 271442 514170 271498 514226
rect 271318 514046 271374 514102
rect 271442 514046 271498 514102
rect 271318 513922 271374 513978
rect 271442 513922 271498 513978
rect 302038 514294 302094 514350
rect 302162 514294 302218 514350
rect 302038 514170 302094 514226
rect 302162 514170 302218 514226
rect 302038 514046 302094 514102
rect 302162 514046 302218 514102
rect 302038 513922 302094 513978
rect 302162 513922 302218 513978
rect 332758 514294 332814 514350
rect 332882 514294 332938 514350
rect 332758 514170 332814 514226
rect 332882 514170 332938 514226
rect 332758 514046 332814 514102
rect 332882 514046 332938 514102
rect 332758 513922 332814 513978
rect 332882 513922 332938 513978
rect 363478 514294 363534 514350
rect 363602 514294 363658 514350
rect 363478 514170 363534 514226
rect 363602 514170 363658 514226
rect 363478 514046 363534 514102
rect 363602 514046 363658 514102
rect 363478 513922 363534 513978
rect 363602 513922 363658 513978
rect 394198 514294 394254 514350
rect 394322 514294 394378 514350
rect 394198 514170 394254 514226
rect 394322 514170 394378 514226
rect 394198 514046 394254 514102
rect 394322 514046 394378 514102
rect 394198 513922 394254 513978
rect 394322 513922 394378 513978
rect 424918 514294 424974 514350
rect 425042 514294 425098 514350
rect 424918 514170 424974 514226
rect 425042 514170 425098 514226
rect 424918 514046 424974 514102
rect 425042 514046 425098 514102
rect 424918 513922 424974 513978
rect 425042 513922 425098 513978
rect 455638 514294 455694 514350
rect 455762 514294 455818 514350
rect 455638 514170 455694 514226
rect 455762 514170 455818 514226
rect 455638 514046 455694 514102
rect 455762 514046 455818 514102
rect 455638 513922 455694 513978
rect 455762 513922 455818 513978
rect 486358 514294 486414 514350
rect 486482 514294 486538 514350
rect 486358 514170 486414 514226
rect 486482 514170 486538 514226
rect 486358 514046 486414 514102
rect 486482 514046 486538 514102
rect 486358 513922 486414 513978
rect 486482 513922 486538 513978
rect 194518 508294 194574 508350
rect 194642 508294 194698 508350
rect 194518 508170 194574 508226
rect 194642 508170 194698 508226
rect 194518 508046 194574 508102
rect 194642 508046 194698 508102
rect 194518 507922 194574 507978
rect 194642 507922 194698 507978
rect 225238 508294 225294 508350
rect 225362 508294 225418 508350
rect 225238 508170 225294 508226
rect 225362 508170 225418 508226
rect 225238 508046 225294 508102
rect 225362 508046 225418 508102
rect 225238 507922 225294 507978
rect 225362 507922 225418 507978
rect 255958 508294 256014 508350
rect 256082 508294 256138 508350
rect 255958 508170 256014 508226
rect 256082 508170 256138 508226
rect 255958 508046 256014 508102
rect 256082 508046 256138 508102
rect 255958 507922 256014 507978
rect 256082 507922 256138 507978
rect 286678 508294 286734 508350
rect 286802 508294 286858 508350
rect 286678 508170 286734 508226
rect 286802 508170 286858 508226
rect 286678 508046 286734 508102
rect 286802 508046 286858 508102
rect 286678 507922 286734 507978
rect 286802 507922 286858 507978
rect 317398 508294 317454 508350
rect 317522 508294 317578 508350
rect 317398 508170 317454 508226
rect 317522 508170 317578 508226
rect 317398 508046 317454 508102
rect 317522 508046 317578 508102
rect 317398 507922 317454 507978
rect 317522 507922 317578 507978
rect 348118 508294 348174 508350
rect 348242 508294 348298 508350
rect 348118 508170 348174 508226
rect 348242 508170 348298 508226
rect 348118 508046 348174 508102
rect 348242 508046 348298 508102
rect 348118 507922 348174 507978
rect 348242 507922 348298 507978
rect 378838 508294 378894 508350
rect 378962 508294 379018 508350
rect 378838 508170 378894 508226
rect 378962 508170 379018 508226
rect 378838 508046 378894 508102
rect 378962 508046 379018 508102
rect 378838 507922 378894 507978
rect 378962 507922 379018 507978
rect 409558 508294 409614 508350
rect 409682 508294 409738 508350
rect 409558 508170 409614 508226
rect 409682 508170 409738 508226
rect 409558 508046 409614 508102
rect 409682 508046 409738 508102
rect 409558 507922 409614 507978
rect 409682 507922 409738 507978
rect 440278 508294 440334 508350
rect 440402 508294 440458 508350
rect 440278 508170 440334 508226
rect 440402 508170 440458 508226
rect 440278 508046 440334 508102
rect 440402 508046 440458 508102
rect 440278 507922 440334 507978
rect 440402 507922 440458 507978
rect 470998 508294 471054 508350
rect 471122 508294 471178 508350
rect 470998 508170 471054 508226
rect 471122 508170 471178 508226
rect 470998 508046 471054 508102
rect 471122 508046 471178 508102
rect 470998 507922 471054 507978
rect 471122 507922 471178 507978
rect 501718 508294 501774 508350
rect 501842 508294 501898 508350
rect 501718 508170 501774 508226
rect 501842 508170 501898 508226
rect 501718 508046 501774 508102
rect 501842 508046 501898 508102
rect 501718 507922 501774 507978
rect 501842 507922 501898 507978
rect 209878 496294 209934 496350
rect 210002 496294 210058 496350
rect 209878 496170 209934 496226
rect 210002 496170 210058 496226
rect 209878 496046 209934 496102
rect 210002 496046 210058 496102
rect 209878 495922 209934 495978
rect 210002 495922 210058 495978
rect 240598 496294 240654 496350
rect 240722 496294 240778 496350
rect 240598 496170 240654 496226
rect 240722 496170 240778 496226
rect 240598 496046 240654 496102
rect 240722 496046 240778 496102
rect 240598 495922 240654 495978
rect 240722 495922 240778 495978
rect 271318 496294 271374 496350
rect 271442 496294 271498 496350
rect 271318 496170 271374 496226
rect 271442 496170 271498 496226
rect 271318 496046 271374 496102
rect 271442 496046 271498 496102
rect 271318 495922 271374 495978
rect 271442 495922 271498 495978
rect 302038 496294 302094 496350
rect 302162 496294 302218 496350
rect 302038 496170 302094 496226
rect 302162 496170 302218 496226
rect 302038 496046 302094 496102
rect 302162 496046 302218 496102
rect 302038 495922 302094 495978
rect 302162 495922 302218 495978
rect 332758 496294 332814 496350
rect 332882 496294 332938 496350
rect 332758 496170 332814 496226
rect 332882 496170 332938 496226
rect 332758 496046 332814 496102
rect 332882 496046 332938 496102
rect 332758 495922 332814 495978
rect 332882 495922 332938 495978
rect 363478 496294 363534 496350
rect 363602 496294 363658 496350
rect 363478 496170 363534 496226
rect 363602 496170 363658 496226
rect 363478 496046 363534 496102
rect 363602 496046 363658 496102
rect 363478 495922 363534 495978
rect 363602 495922 363658 495978
rect 394198 496294 394254 496350
rect 394322 496294 394378 496350
rect 394198 496170 394254 496226
rect 394322 496170 394378 496226
rect 394198 496046 394254 496102
rect 394322 496046 394378 496102
rect 394198 495922 394254 495978
rect 394322 495922 394378 495978
rect 424918 496294 424974 496350
rect 425042 496294 425098 496350
rect 424918 496170 424974 496226
rect 425042 496170 425098 496226
rect 424918 496046 424974 496102
rect 425042 496046 425098 496102
rect 424918 495922 424974 495978
rect 425042 495922 425098 495978
rect 455638 496294 455694 496350
rect 455762 496294 455818 496350
rect 455638 496170 455694 496226
rect 455762 496170 455818 496226
rect 455638 496046 455694 496102
rect 455762 496046 455818 496102
rect 455638 495922 455694 495978
rect 455762 495922 455818 495978
rect 486358 496294 486414 496350
rect 486482 496294 486538 496350
rect 486358 496170 486414 496226
rect 486482 496170 486538 496226
rect 486358 496046 486414 496102
rect 486482 496046 486538 496102
rect 486358 495922 486414 495978
rect 486482 495922 486538 495978
rect 194518 490294 194574 490350
rect 194642 490294 194698 490350
rect 194518 490170 194574 490226
rect 194642 490170 194698 490226
rect 194518 490046 194574 490102
rect 194642 490046 194698 490102
rect 194518 489922 194574 489978
rect 194642 489922 194698 489978
rect 225238 490294 225294 490350
rect 225362 490294 225418 490350
rect 225238 490170 225294 490226
rect 225362 490170 225418 490226
rect 225238 490046 225294 490102
rect 225362 490046 225418 490102
rect 225238 489922 225294 489978
rect 225362 489922 225418 489978
rect 255958 490294 256014 490350
rect 256082 490294 256138 490350
rect 255958 490170 256014 490226
rect 256082 490170 256138 490226
rect 255958 490046 256014 490102
rect 256082 490046 256138 490102
rect 255958 489922 256014 489978
rect 256082 489922 256138 489978
rect 286678 490294 286734 490350
rect 286802 490294 286858 490350
rect 286678 490170 286734 490226
rect 286802 490170 286858 490226
rect 286678 490046 286734 490102
rect 286802 490046 286858 490102
rect 286678 489922 286734 489978
rect 286802 489922 286858 489978
rect 317398 490294 317454 490350
rect 317522 490294 317578 490350
rect 317398 490170 317454 490226
rect 317522 490170 317578 490226
rect 317398 490046 317454 490102
rect 317522 490046 317578 490102
rect 317398 489922 317454 489978
rect 317522 489922 317578 489978
rect 348118 490294 348174 490350
rect 348242 490294 348298 490350
rect 348118 490170 348174 490226
rect 348242 490170 348298 490226
rect 348118 490046 348174 490102
rect 348242 490046 348298 490102
rect 348118 489922 348174 489978
rect 348242 489922 348298 489978
rect 378838 490294 378894 490350
rect 378962 490294 379018 490350
rect 378838 490170 378894 490226
rect 378962 490170 379018 490226
rect 378838 490046 378894 490102
rect 378962 490046 379018 490102
rect 378838 489922 378894 489978
rect 378962 489922 379018 489978
rect 409558 490294 409614 490350
rect 409682 490294 409738 490350
rect 409558 490170 409614 490226
rect 409682 490170 409738 490226
rect 409558 490046 409614 490102
rect 409682 490046 409738 490102
rect 409558 489922 409614 489978
rect 409682 489922 409738 489978
rect 440278 490294 440334 490350
rect 440402 490294 440458 490350
rect 440278 490170 440334 490226
rect 440402 490170 440458 490226
rect 440278 490046 440334 490102
rect 440402 490046 440458 490102
rect 440278 489922 440334 489978
rect 440402 489922 440458 489978
rect 470998 490294 471054 490350
rect 471122 490294 471178 490350
rect 470998 490170 471054 490226
rect 471122 490170 471178 490226
rect 470998 490046 471054 490102
rect 471122 490046 471178 490102
rect 470998 489922 471054 489978
rect 471122 489922 471178 489978
rect 501718 490294 501774 490350
rect 501842 490294 501898 490350
rect 501718 490170 501774 490226
rect 501842 490170 501898 490226
rect 501718 490046 501774 490102
rect 501842 490046 501898 490102
rect 501718 489922 501774 489978
rect 501842 489922 501898 489978
rect 209878 478294 209934 478350
rect 210002 478294 210058 478350
rect 209878 478170 209934 478226
rect 210002 478170 210058 478226
rect 209878 478046 209934 478102
rect 210002 478046 210058 478102
rect 209878 477922 209934 477978
rect 210002 477922 210058 477978
rect 240598 478294 240654 478350
rect 240722 478294 240778 478350
rect 240598 478170 240654 478226
rect 240722 478170 240778 478226
rect 240598 478046 240654 478102
rect 240722 478046 240778 478102
rect 240598 477922 240654 477978
rect 240722 477922 240778 477978
rect 271318 478294 271374 478350
rect 271442 478294 271498 478350
rect 271318 478170 271374 478226
rect 271442 478170 271498 478226
rect 271318 478046 271374 478102
rect 271442 478046 271498 478102
rect 271318 477922 271374 477978
rect 271442 477922 271498 477978
rect 302038 478294 302094 478350
rect 302162 478294 302218 478350
rect 302038 478170 302094 478226
rect 302162 478170 302218 478226
rect 302038 478046 302094 478102
rect 302162 478046 302218 478102
rect 302038 477922 302094 477978
rect 302162 477922 302218 477978
rect 332758 478294 332814 478350
rect 332882 478294 332938 478350
rect 332758 478170 332814 478226
rect 332882 478170 332938 478226
rect 332758 478046 332814 478102
rect 332882 478046 332938 478102
rect 332758 477922 332814 477978
rect 332882 477922 332938 477978
rect 363478 478294 363534 478350
rect 363602 478294 363658 478350
rect 363478 478170 363534 478226
rect 363602 478170 363658 478226
rect 363478 478046 363534 478102
rect 363602 478046 363658 478102
rect 363478 477922 363534 477978
rect 363602 477922 363658 477978
rect 394198 478294 394254 478350
rect 394322 478294 394378 478350
rect 394198 478170 394254 478226
rect 394322 478170 394378 478226
rect 394198 478046 394254 478102
rect 394322 478046 394378 478102
rect 394198 477922 394254 477978
rect 394322 477922 394378 477978
rect 424918 478294 424974 478350
rect 425042 478294 425098 478350
rect 424918 478170 424974 478226
rect 425042 478170 425098 478226
rect 424918 478046 424974 478102
rect 425042 478046 425098 478102
rect 424918 477922 424974 477978
rect 425042 477922 425098 477978
rect 455638 478294 455694 478350
rect 455762 478294 455818 478350
rect 455638 478170 455694 478226
rect 455762 478170 455818 478226
rect 455638 478046 455694 478102
rect 455762 478046 455818 478102
rect 455638 477922 455694 477978
rect 455762 477922 455818 477978
rect 486358 478294 486414 478350
rect 486482 478294 486538 478350
rect 486358 478170 486414 478226
rect 486482 478170 486538 478226
rect 486358 478046 486414 478102
rect 486482 478046 486538 478102
rect 486358 477922 486414 477978
rect 486482 477922 486538 477978
rect 194518 472294 194574 472350
rect 194642 472294 194698 472350
rect 194518 472170 194574 472226
rect 194642 472170 194698 472226
rect 194518 472046 194574 472102
rect 194642 472046 194698 472102
rect 194518 471922 194574 471978
rect 194642 471922 194698 471978
rect 225238 472294 225294 472350
rect 225362 472294 225418 472350
rect 225238 472170 225294 472226
rect 225362 472170 225418 472226
rect 225238 472046 225294 472102
rect 225362 472046 225418 472102
rect 225238 471922 225294 471978
rect 225362 471922 225418 471978
rect 255958 472294 256014 472350
rect 256082 472294 256138 472350
rect 255958 472170 256014 472226
rect 256082 472170 256138 472226
rect 255958 472046 256014 472102
rect 256082 472046 256138 472102
rect 255958 471922 256014 471978
rect 256082 471922 256138 471978
rect 286678 472294 286734 472350
rect 286802 472294 286858 472350
rect 286678 472170 286734 472226
rect 286802 472170 286858 472226
rect 286678 472046 286734 472102
rect 286802 472046 286858 472102
rect 286678 471922 286734 471978
rect 286802 471922 286858 471978
rect 317398 472294 317454 472350
rect 317522 472294 317578 472350
rect 317398 472170 317454 472226
rect 317522 472170 317578 472226
rect 317398 472046 317454 472102
rect 317522 472046 317578 472102
rect 317398 471922 317454 471978
rect 317522 471922 317578 471978
rect 348118 472294 348174 472350
rect 348242 472294 348298 472350
rect 348118 472170 348174 472226
rect 348242 472170 348298 472226
rect 348118 472046 348174 472102
rect 348242 472046 348298 472102
rect 348118 471922 348174 471978
rect 348242 471922 348298 471978
rect 378838 472294 378894 472350
rect 378962 472294 379018 472350
rect 378838 472170 378894 472226
rect 378962 472170 379018 472226
rect 378838 472046 378894 472102
rect 378962 472046 379018 472102
rect 378838 471922 378894 471978
rect 378962 471922 379018 471978
rect 409558 472294 409614 472350
rect 409682 472294 409738 472350
rect 409558 472170 409614 472226
rect 409682 472170 409738 472226
rect 409558 472046 409614 472102
rect 409682 472046 409738 472102
rect 409558 471922 409614 471978
rect 409682 471922 409738 471978
rect 440278 472294 440334 472350
rect 440402 472294 440458 472350
rect 440278 472170 440334 472226
rect 440402 472170 440458 472226
rect 440278 472046 440334 472102
rect 440402 472046 440458 472102
rect 440278 471922 440334 471978
rect 440402 471922 440458 471978
rect 470998 472294 471054 472350
rect 471122 472294 471178 472350
rect 470998 472170 471054 472226
rect 471122 472170 471178 472226
rect 470998 472046 471054 472102
rect 471122 472046 471178 472102
rect 470998 471922 471054 471978
rect 471122 471922 471178 471978
rect 501718 472294 501774 472350
rect 501842 472294 501898 472350
rect 501718 472170 501774 472226
rect 501842 472170 501898 472226
rect 501718 472046 501774 472102
rect 501842 472046 501898 472102
rect 501718 471922 501774 471978
rect 501842 471922 501898 471978
rect 209878 460294 209934 460350
rect 210002 460294 210058 460350
rect 209878 460170 209934 460226
rect 210002 460170 210058 460226
rect 209878 460046 209934 460102
rect 210002 460046 210058 460102
rect 209878 459922 209934 459978
rect 210002 459922 210058 459978
rect 240598 460294 240654 460350
rect 240722 460294 240778 460350
rect 240598 460170 240654 460226
rect 240722 460170 240778 460226
rect 240598 460046 240654 460102
rect 240722 460046 240778 460102
rect 240598 459922 240654 459978
rect 240722 459922 240778 459978
rect 271318 460294 271374 460350
rect 271442 460294 271498 460350
rect 271318 460170 271374 460226
rect 271442 460170 271498 460226
rect 271318 460046 271374 460102
rect 271442 460046 271498 460102
rect 271318 459922 271374 459978
rect 271442 459922 271498 459978
rect 302038 460294 302094 460350
rect 302162 460294 302218 460350
rect 302038 460170 302094 460226
rect 302162 460170 302218 460226
rect 302038 460046 302094 460102
rect 302162 460046 302218 460102
rect 302038 459922 302094 459978
rect 302162 459922 302218 459978
rect 332758 460294 332814 460350
rect 332882 460294 332938 460350
rect 332758 460170 332814 460226
rect 332882 460170 332938 460226
rect 332758 460046 332814 460102
rect 332882 460046 332938 460102
rect 332758 459922 332814 459978
rect 332882 459922 332938 459978
rect 363478 460294 363534 460350
rect 363602 460294 363658 460350
rect 363478 460170 363534 460226
rect 363602 460170 363658 460226
rect 363478 460046 363534 460102
rect 363602 460046 363658 460102
rect 363478 459922 363534 459978
rect 363602 459922 363658 459978
rect 394198 460294 394254 460350
rect 394322 460294 394378 460350
rect 394198 460170 394254 460226
rect 394322 460170 394378 460226
rect 394198 460046 394254 460102
rect 394322 460046 394378 460102
rect 394198 459922 394254 459978
rect 394322 459922 394378 459978
rect 424918 460294 424974 460350
rect 425042 460294 425098 460350
rect 424918 460170 424974 460226
rect 425042 460170 425098 460226
rect 424918 460046 424974 460102
rect 425042 460046 425098 460102
rect 424918 459922 424974 459978
rect 425042 459922 425098 459978
rect 455638 460294 455694 460350
rect 455762 460294 455818 460350
rect 455638 460170 455694 460226
rect 455762 460170 455818 460226
rect 455638 460046 455694 460102
rect 455762 460046 455818 460102
rect 455638 459922 455694 459978
rect 455762 459922 455818 459978
rect 486358 460294 486414 460350
rect 486482 460294 486538 460350
rect 486358 460170 486414 460226
rect 486482 460170 486538 460226
rect 486358 460046 486414 460102
rect 486482 460046 486538 460102
rect 486358 459922 486414 459978
rect 486482 459922 486538 459978
rect 194518 454294 194574 454350
rect 194642 454294 194698 454350
rect 194518 454170 194574 454226
rect 194642 454170 194698 454226
rect 194518 454046 194574 454102
rect 194642 454046 194698 454102
rect 194518 453922 194574 453978
rect 194642 453922 194698 453978
rect 225238 454294 225294 454350
rect 225362 454294 225418 454350
rect 225238 454170 225294 454226
rect 225362 454170 225418 454226
rect 225238 454046 225294 454102
rect 225362 454046 225418 454102
rect 225238 453922 225294 453978
rect 225362 453922 225418 453978
rect 255958 454294 256014 454350
rect 256082 454294 256138 454350
rect 255958 454170 256014 454226
rect 256082 454170 256138 454226
rect 255958 454046 256014 454102
rect 256082 454046 256138 454102
rect 255958 453922 256014 453978
rect 256082 453922 256138 453978
rect 286678 454294 286734 454350
rect 286802 454294 286858 454350
rect 286678 454170 286734 454226
rect 286802 454170 286858 454226
rect 286678 454046 286734 454102
rect 286802 454046 286858 454102
rect 286678 453922 286734 453978
rect 286802 453922 286858 453978
rect 317398 454294 317454 454350
rect 317522 454294 317578 454350
rect 317398 454170 317454 454226
rect 317522 454170 317578 454226
rect 317398 454046 317454 454102
rect 317522 454046 317578 454102
rect 317398 453922 317454 453978
rect 317522 453922 317578 453978
rect 348118 454294 348174 454350
rect 348242 454294 348298 454350
rect 348118 454170 348174 454226
rect 348242 454170 348298 454226
rect 348118 454046 348174 454102
rect 348242 454046 348298 454102
rect 348118 453922 348174 453978
rect 348242 453922 348298 453978
rect 378838 454294 378894 454350
rect 378962 454294 379018 454350
rect 378838 454170 378894 454226
rect 378962 454170 379018 454226
rect 378838 454046 378894 454102
rect 378962 454046 379018 454102
rect 378838 453922 378894 453978
rect 378962 453922 379018 453978
rect 409558 454294 409614 454350
rect 409682 454294 409738 454350
rect 409558 454170 409614 454226
rect 409682 454170 409738 454226
rect 409558 454046 409614 454102
rect 409682 454046 409738 454102
rect 409558 453922 409614 453978
rect 409682 453922 409738 453978
rect 440278 454294 440334 454350
rect 440402 454294 440458 454350
rect 440278 454170 440334 454226
rect 440402 454170 440458 454226
rect 440278 454046 440334 454102
rect 440402 454046 440458 454102
rect 440278 453922 440334 453978
rect 440402 453922 440458 453978
rect 470998 454294 471054 454350
rect 471122 454294 471178 454350
rect 470998 454170 471054 454226
rect 471122 454170 471178 454226
rect 470998 454046 471054 454102
rect 471122 454046 471178 454102
rect 470998 453922 471054 453978
rect 471122 453922 471178 453978
rect 501718 454294 501774 454350
rect 501842 454294 501898 454350
rect 501718 454170 501774 454226
rect 501842 454170 501898 454226
rect 501718 454046 501774 454102
rect 501842 454046 501898 454102
rect 501718 453922 501774 453978
rect 501842 453922 501898 453978
rect 209878 442294 209934 442350
rect 210002 442294 210058 442350
rect 209878 442170 209934 442226
rect 210002 442170 210058 442226
rect 209878 442046 209934 442102
rect 210002 442046 210058 442102
rect 209878 441922 209934 441978
rect 210002 441922 210058 441978
rect 240598 442294 240654 442350
rect 240722 442294 240778 442350
rect 240598 442170 240654 442226
rect 240722 442170 240778 442226
rect 240598 442046 240654 442102
rect 240722 442046 240778 442102
rect 240598 441922 240654 441978
rect 240722 441922 240778 441978
rect 271318 442294 271374 442350
rect 271442 442294 271498 442350
rect 271318 442170 271374 442226
rect 271442 442170 271498 442226
rect 271318 442046 271374 442102
rect 271442 442046 271498 442102
rect 271318 441922 271374 441978
rect 271442 441922 271498 441978
rect 302038 442294 302094 442350
rect 302162 442294 302218 442350
rect 302038 442170 302094 442226
rect 302162 442170 302218 442226
rect 302038 442046 302094 442102
rect 302162 442046 302218 442102
rect 302038 441922 302094 441978
rect 302162 441922 302218 441978
rect 332758 442294 332814 442350
rect 332882 442294 332938 442350
rect 332758 442170 332814 442226
rect 332882 442170 332938 442226
rect 332758 442046 332814 442102
rect 332882 442046 332938 442102
rect 332758 441922 332814 441978
rect 332882 441922 332938 441978
rect 363478 442294 363534 442350
rect 363602 442294 363658 442350
rect 363478 442170 363534 442226
rect 363602 442170 363658 442226
rect 363478 442046 363534 442102
rect 363602 442046 363658 442102
rect 363478 441922 363534 441978
rect 363602 441922 363658 441978
rect 394198 442294 394254 442350
rect 394322 442294 394378 442350
rect 394198 442170 394254 442226
rect 394322 442170 394378 442226
rect 394198 442046 394254 442102
rect 394322 442046 394378 442102
rect 394198 441922 394254 441978
rect 394322 441922 394378 441978
rect 424918 442294 424974 442350
rect 425042 442294 425098 442350
rect 424918 442170 424974 442226
rect 425042 442170 425098 442226
rect 424918 442046 424974 442102
rect 425042 442046 425098 442102
rect 424918 441922 424974 441978
rect 425042 441922 425098 441978
rect 455638 442294 455694 442350
rect 455762 442294 455818 442350
rect 455638 442170 455694 442226
rect 455762 442170 455818 442226
rect 455638 442046 455694 442102
rect 455762 442046 455818 442102
rect 455638 441922 455694 441978
rect 455762 441922 455818 441978
rect 486358 442294 486414 442350
rect 486482 442294 486538 442350
rect 486358 442170 486414 442226
rect 486482 442170 486538 442226
rect 486358 442046 486414 442102
rect 486482 442046 486538 442102
rect 486358 441922 486414 441978
rect 486482 441922 486538 441978
rect 194518 436294 194574 436350
rect 194642 436294 194698 436350
rect 194518 436170 194574 436226
rect 194642 436170 194698 436226
rect 194518 436046 194574 436102
rect 194642 436046 194698 436102
rect 194518 435922 194574 435978
rect 194642 435922 194698 435978
rect 225238 436294 225294 436350
rect 225362 436294 225418 436350
rect 225238 436170 225294 436226
rect 225362 436170 225418 436226
rect 225238 436046 225294 436102
rect 225362 436046 225418 436102
rect 225238 435922 225294 435978
rect 225362 435922 225418 435978
rect 255958 436294 256014 436350
rect 256082 436294 256138 436350
rect 255958 436170 256014 436226
rect 256082 436170 256138 436226
rect 255958 436046 256014 436102
rect 256082 436046 256138 436102
rect 255958 435922 256014 435978
rect 256082 435922 256138 435978
rect 286678 436294 286734 436350
rect 286802 436294 286858 436350
rect 286678 436170 286734 436226
rect 286802 436170 286858 436226
rect 286678 436046 286734 436102
rect 286802 436046 286858 436102
rect 286678 435922 286734 435978
rect 286802 435922 286858 435978
rect 317398 436294 317454 436350
rect 317522 436294 317578 436350
rect 317398 436170 317454 436226
rect 317522 436170 317578 436226
rect 317398 436046 317454 436102
rect 317522 436046 317578 436102
rect 317398 435922 317454 435978
rect 317522 435922 317578 435978
rect 348118 436294 348174 436350
rect 348242 436294 348298 436350
rect 348118 436170 348174 436226
rect 348242 436170 348298 436226
rect 348118 436046 348174 436102
rect 348242 436046 348298 436102
rect 348118 435922 348174 435978
rect 348242 435922 348298 435978
rect 378838 436294 378894 436350
rect 378962 436294 379018 436350
rect 378838 436170 378894 436226
rect 378962 436170 379018 436226
rect 378838 436046 378894 436102
rect 378962 436046 379018 436102
rect 378838 435922 378894 435978
rect 378962 435922 379018 435978
rect 409558 436294 409614 436350
rect 409682 436294 409738 436350
rect 409558 436170 409614 436226
rect 409682 436170 409738 436226
rect 409558 436046 409614 436102
rect 409682 436046 409738 436102
rect 409558 435922 409614 435978
rect 409682 435922 409738 435978
rect 440278 436294 440334 436350
rect 440402 436294 440458 436350
rect 440278 436170 440334 436226
rect 440402 436170 440458 436226
rect 440278 436046 440334 436102
rect 440402 436046 440458 436102
rect 440278 435922 440334 435978
rect 440402 435922 440458 435978
rect 470998 436294 471054 436350
rect 471122 436294 471178 436350
rect 470998 436170 471054 436226
rect 471122 436170 471178 436226
rect 470998 436046 471054 436102
rect 471122 436046 471178 436102
rect 470998 435922 471054 435978
rect 471122 435922 471178 435978
rect 501718 436294 501774 436350
rect 501842 436294 501898 436350
rect 501718 436170 501774 436226
rect 501842 436170 501898 436226
rect 501718 436046 501774 436102
rect 501842 436046 501898 436102
rect 501718 435922 501774 435978
rect 501842 435922 501898 435978
rect 209878 424294 209934 424350
rect 210002 424294 210058 424350
rect 209878 424170 209934 424226
rect 210002 424170 210058 424226
rect 209878 424046 209934 424102
rect 210002 424046 210058 424102
rect 209878 423922 209934 423978
rect 210002 423922 210058 423978
rect 240598 424294 240654 424350
rect 240722 424294 240778 424350
rect 240598 424170 240654 424226
rect 240722 424170 240778 424226
rect 240598 424046 240654 424102
rect 240722 424046 240778 424102
rect 240598 423922 240654 423978
rect 240722 423922 240778 423978
rect 271318 424294 271374 424350
rect 271442 424294 271498 424350
rect 271318 424170 271374 424226
rect 271442 424170 271498 424226
rect 271318 424046 271374 424102
rect 271442 424046 271498 424102
rect 271318 423922 271374 423978
rect 271442 423922 271498 423978
rect 302038 424294 302094 424350
rect 302162 424294 302218 424350
rect 302038 424170 302094 424226
rect 302162 424170 302218 424226
rect 302038 424046 302094 424102
rect 302162 424046 302218 424102
rect 302038 423922 302094 423978
rect 302162 423922 302218 423978
rect 332758 424294 332814 424350
rect 332882 424294 332938 424350
rect 332758 424170 332814 424226
rect 332882 424170 332938 424226
rect 332758 424046 332814 424102
rect 332882 424046 332938 424102
rect 332758 423922 332814 423978
rect 332882 423922 332938 423978
rect 363478 424294 363534 424350
rect 363602 424294 363658 424350
rect 363478 424170 363534 424226
rect 363602 424170 363658 424226
rect 363478 424046 363534 424102
rect 363602 424046 363658 424102
rect 363478 423922 363534 423978
rect 363602 423922 363658 423978
rect 394198 424294 394254 424350
rect 394322 424294 394378 424350
rect 394198 424170 394254 424226
rect 394322 424170 394378 424226
rect 394198 424046 394254 424102
rect 394322 424046 394378 424102
rect 394198 423922 394254 423978
rect 394322 423922 394378 423978
rect 424918 424294 424974 424350
rect 425042 424294 425098 424350
rect 424918 424170 424974 424226
rect 425042 424170 425098 424226
rect 424918 424046 424974 424102
rect 425042 424046 425098 424102
rect 424918 423922 424974 423978
rect 425042 423922 425098 423978
rect 455638 424294 455694 424350
rect 455762 424294 455818 424350
rect 455638 424170 455694 424226
rect 455762 424170 455818 424226
rect 455638 424046 455694 424102
rect 455762 424046 455818 424102
rect 455638 423922 455694 423978
rect 455762 423922 455818 423978
rect 486358 424294 486414 424350
rect 486482 424294 486538 424350
rect 486358 424170 486414 424226
rect 486482 424170 486538 424226
rect 486358 424046 486414 424102
rect 486482 424046 486538 424102
rect 486358 423922 486414 423978
rect 486482 423922 486538 423978
rect 194518 418294 194574 418350
rect 194642 418294 194698 418350
rect 194518 418170 194574 418226
rect 194642 418170 194698 418226
rect 194518 418046 194574 418102
rect 194642 418046 194698 418102
rect 194518 417922 194574 417978
rect 194642 417922 194698 417978
rect 225238 418294 225294 418350
rect 225362 418294 225418 418350
rect 225238 418170 225294 418226
rect 225362 418170 225418 418226
rect 225238 418046 225294 418102
rect 225362 418046 225418 418102
rect 225238 417922 225294 417978
rect 225362 417922 225418 417978
rect 255958 418294 256014 418350
rect 256082 418294 256138 418350
rect 255958 418170 256014 418226
rect 256082 418170 256138 418226
rect 255958 418046 256014 418102
rect 256082 418046 256138 418102
rect 255958 417922 256014 417978
rect 256082 417922 256138 417978
rect 286678 418294 286734 418350
rect 286802 418294 286858 418350
rect 286678 418170 286734 418226
rect 286802 418170 286858 418226
rect 286678 418046 286734 418102
rect 286802 418046 286858 418102
rect 286678 417922 286734 417978
rect 286802 417922 286858 417978
rect 317398 418294 317454 418350
rect 317522 418294 317578 418350
rect 317398 418170 317454 418226
rect 317522 418170 317578 418226
rect 317398 418046 317454 418102
rect 317522 418046 317578 418102
rect 317398 417922 317454 417978
rect 317522 417922 317578 417978
rect 348118 418294 348174 418350
rect 348242 418294 348298 418350
rect 348118 418170 348174 418226
rect 348242 418170 348298 418226
rect 348118 418046 348174 418102
rect 348242 418046 348298 418102
rect 348118 417922 348174 417978
rect 348242 417922 348298 417978
rect 378838 418294 378894 418350
rect 378962 418294 379018 418350
rect 378838 418170 378894 418226
rect 378962 418170 379018 418226
rect 378838 418046 378894 418102
rect 378962 418046 379018 418102
rect 378838 417922 378894 417978
rect 378962 417922 379018 417978
rect 409558 418294 409614 418350
rect 409682 418294 409738 418350
rect 409558 418170 409614 418226
rect 409682 418170 409738 418226
rect 409558 418046 409614 418102
rect 409682 418046 409738 418102
rect 409558 417922 409614 417978
rect 409682 417922 409738 417978
rect 440278 418294 440334 418350
rect 440402 418294 440458 418350
rect 440278 418170 440334 418226
rect 440402 418170 440458 418226
rect 440278 418046 440334 418102
rect 440402 418046 440458 418102
rect 440278 417922 440334 417978
rect 440402 417922 440458 417978
rect 470998 418294 471054 418350
rect 471122 418294 471178 418350
rect 470998 418170 471054 418226
rect 471122 418170 471178 418226
rect 470998 418046 471054 418102
rect 471122 418046 471178 418102
rect 470998 417922 471054 417978
rect 471122 417922 471178 417978
rect 501718 418294 501774 418350
rect 501842 418294 501898 418350
rect 501718 418170 501774 418226
rect 501842 418170 501898 418226
rect 501718 418046 501774 418102
rect 501842 418046 501898 418102
rect 501718 417922 501774 417978
rect 501842 417922 501898 417978
rect 357196 411002 357252 411058
rect 334236 410822 334292 410878
rect 324156 410642 324212 410698
rect 209916 404522 209972 404578
rect 208236 404342 208292 404398
rect 206556 404162 206612 404218
rect 193554 388294 193610 388350
rect 193678 388294 193734 388350
rect 193802 388294 193858 388350
rect 193926 388294 193982 388350
rect 193554 388170 193610 388226
rect 193678 388170 193734 388226
rect 193802 388170 193858 388226
rect 193926 388170 193982 388226
rect 193554 388046 193610 388102
rect 193678 388046 193734 388102
rect 193802 388046 193858 388102
rect 193926 388046 193982 388102
rect 193554 387922 193610 387978
rect 193678 387922 193734 387978
rect 193802 387922 193858 387978
rect 193926 387922 193982 387978
rect 189834 364294 189890 364350
rect 189958 364294 190014 364350
rect 190082 364294 190138 364350
rect 190206 364294 190262 364350
rect 189834 364170 189890 364226
rect 189958 364170 190014 364226
rect 190082 364170 190138 364226
rect 190206 364170 190262 364226
rect 189834 364046 189890 364102
rect 189958 364046 190014 364102
rect 190082 364046 190138 364102
rect 190206 364046 190262 364102
rect 189834 363922 189890 363978
rect 189958 363922 190014 363978
rect 190082 363922 190138 363978
rect 190206 363922 190262 363978
rect 189834 346294 189890 346350
rect 189958 346294 190014 346350
rect 190082 346294 190138 346350
rect 190206 346294 190262 346350
rect 189834 346170 189890 346226
rect 189958 346170 190014 346226
rect 190082 346170 190138 346226
rect 190206 346170 190262 346226
rect 189834 346046 189890 346102
rect 189958 346046 190014 346102
rect 190082 346046 190138 346102
rect 190206 346046 190262 346102
rect 189834 345922 189890 345978
rect 189958 345922 190014 345978
rect 190082 345922 190138 345978
rect 190206 345922 190262 345978
rect 189834 328294 189890 328350
rect 189958 328294 190014 328350
rect 190082 328294 190138 328350
rect 190206 328294 190262 328350
rect 189834 328170 189890 328226
rect 189958 328170 190014 328226
rect 190082 328170 190138 328226
rect 190206 328170 190262 328226
rect 189834 328046 189890 328102
rect 189958 328046 190014 328102
rect 190082 328046 190138 328102
rect 190206 328046 190262 328102
rect 189834 327922 189890 327978
rect 189958 327922 190014 327978
rect 190082 327922 190138 327978
rect 190206 327922 190262 327978
rect 196476 402002 196532 402058
rect 198156 401822 198212 401878
rect 198044 393182 198100 393238
rect 197484 391742 197540 391798
rect 193554 370294 193610 370350
rect 193678 370294 193734 370350
rect 193802 370294 193858 370350
rect 193926 370294 193982 370350
rect 193554 370170 193610 370226
rect 193678 370170 193734 370226
rect 193802 370170 193858 370226
rect 193926 370170 193982 370226
rect 193554 370046 193610 370102
rect 193678 370046 193734 370102
rect 193802 370046 193858 370102
rect 193926 370046 193982 370102
rect 193554 369922 193610 369978
rect 193678 369922 193734 369978
rect 193802 369922 193858 369978
rect 193926 369922 193982 369978
rect 194518 364294 194574 364350
rect 194642 364294 194698 364350
rect 194518 364170 194574 364226
rect 194642 364170 194698 364226
rect 194518 364046 194574 364102
rect 194642 364046 194698 364102
rect 194518 363922 194574 363978
rect 194642 363922 194698 363978
rect 193554 352294 193610 352350
rect 193678 352294 193734 352350
rect 193802 352294 193858 352350
rect 193926 352294 193982 352350
rect 193554 352170 193610 352226
rect 193678 352170 193734 352226
rect 193802 352170 193858 352226
rect 193926 352170 193982 352226
rect 193554 352046 193610 352102
rect 193678 352046 193734 352102
rect 193802 352046 193858 352102
rect 193926 352046 193982 352102
rect 193554 351922 193610 351978
rect 193678 351922 193734 351978
rect 193802 351922 193858 351978
rect 193926 351922 193982 351978
rect 194518 346294 194574 346350
rect 194642 346294 194698 346350
rect 194518 346170 194574 346226
rect 194642 346170 194698 346226
rect 194518 346046 194574 346102
rect 194642 346046 194698 346102
rect 194518 345922 194574 345978
rect 194642 345922 194698 345978
rect 193554 334294 193610 334350
rect 193678 334294 193734 334350
rect 193802 334294 193858 334350
rect 193926 334294 193982 334350
rect 193554 334170 193610 334226
rect 193678 334170 193734 334226
rect 193802 334170 193858 334226
rect 193926 334170 193982 334226
rect 193554 334046 193610 334102
rect 193678 334046 193734 334102
rect 193802 334046 193858 334102
rect 193926 334046 193982 334102
rect 193554 333922 193610 333978
rect 193678 333922 193734 333978
rect 193802 333922 193858 333978
rect 193926 333922 193982 333978
rect 190652 323372 190708 323398
rect 190652 323342 190708 323372
rect 192332 323342 192388 323398
rect 189834 310294 189890 310350
rect 189958 310294 190014 310350
rect 190082 310294 190138 310350
rect 190206 310294 190262 310350
rect 189834 310170 189890 310226
rect 189958 310170 190014 310226
rect 190082 310170 190138 310226
rect 190206 310170 190262 310226
rect 189834 310046 189890 310102
rect 189958 310046 190014 310102
rect 190082 310046 190138 310102
rect 190206 310046 190262 310102
rect 189834 309922 189890 309978
rect 189958 309922 190014 309978
rect 190082 309922 190138 309978
rect 190206 309922 190262 309978
rect 189834 292294 189890 292350
rect 189958 292294 190014 292350
rect 190082 292294 190138 292350
rect 190206 292294 190262 292350
rect 189834 292170 189890 292226
rect 189958 292170 190014 292226
rect 190082 292170 190138 292226
rect 190206 292170 190262 292226
rect 189834 292046 189890 292102
rect 189958 292046 190014 292102
rect 190082 292046 190138 292102
rect 190206 292046 190262 292102
rect 189834 291922 189890 291978
rect 189958 291922 190014 291978
rect 190082 291922 190138 291978
rect 190206 291922 190262 291978
rect 188076 285722 188132 285778
rect 187852 281402 187908 281458
rect 189834 274294 189890 274350
rect 189958 274294 190014 274350
rect 190082 274294 190138 274350
rect 190206 274294 190262 274350
rect 189834 274170 189890 274226
rect 189958 274170 190014 274226
rect 190082 274170 190138 274226
rect 190206 274170 190262 274226
rect 189834 274046 189890 274102
rect 189958 274046 190014 274102
rect 190082 274046 190138 274102
rect 190206 274046 190262 274102
rect 189834 273922 189890 273978
rect 189958 273922 190014 273978
rect 190082 273922 190138 273978
rect 190206 273922 190262 273978
rect 189834 256294 189890 256350
rect 189958 256294 190014 256350
rect 190082 256294 190138 256350
rect 190206 256294 190262 256350
rect 189834 256170 189890 256226
rect 189958 256170 190014 256226
rect 190082 256170 190138 256226
rect 190206 256170 190262 256226
rect 189834 256046 189890 256102
rect 189958 256046 190014 256102
rect 190082 256046 190138 256102
rect 190206 256046 190262 256102
rect 189834 255922 189890 255978
rect 189958 255922 190014 255978
rect 190082 255922 190138 255978
rect 190206 255922 190262 255978
rect 187852 214082 187908 214138
rect 189834 238294 189890 238350
rect 189958 238294 190014 238350
rect 190082 238294 190138 238350
rect 190206 238294 190262 238350
rect 189834 238170 189890 238226
rect 189958 238170 190014 238226
rect 190082 238170 190138 238226
rect 190206 238170 190262 238226
rect 189834 238046 189890 238102
rect 189958 238046 190014 238102
rect 190082 238046 190138 238102
rect 190206 238046 190262 238102
rect 189834 237922 189890 237978
rect 189958 237922 190014 237978
rect 190082 237922 190138 237978
rect 190206 237922 190262 237978
rect 189834 220294 189890 220350
rect 189958 220294 190014 220350
rect 190082 220294 190138 220350
rect 190206 220294 190262 220350
rect 189834 220170 189890 220226
rect 189958 220170 190014 220226
rect 190082 220170 190138 220226
rect 190206 220170 190262 220226
rect 189834 220046 189890 220102
rect 189958 220046 190014 220102
rect 190082 220046 190138 220102
rect 190206 220046 190262 220102
rect 189834 219922 189890 219978
rect 189958 219922 190014 219978
rect 190082 219922 190138 219978
rect 190206 219922 190262 219978
rect 190652 249722 190708 249778
rect 190652 248642 190708 248698
rect 190652 247212 190708 247258
rect 190652 247202 190708 247212
rect 190876 243062 190932 243118
rect 190652 241982 190708 242038
rect 190652 234962 190708 235018
rect 192332 214442 192388 214498
rect 194518 328294 194574 328350
rect 194642 328294 194698 328350
rect 194518 328170 194574 328226
rect 194642 328170 194698 328226
rect 194518 328046 194574 328102
rect 194642 328046 194698 328102
rect 194518 327922 194574 327978
rect 194642 327922 194698 327978
rect 193554 316294 193610 316350
rect 193678 316294 193734 316350
rect 193802 316294 193858 316350
rect 193926 316294 193982 316350
rect 193554 316170 193610 316226
rect 193678 316170 193734 316226
rect 193802 316170 193858 316226
rect 193926 316170 193982 316226
rect 193554 316046 193610 316102
rect 193678 316046 193734 316102
rect 193802 316046 193858 316102
rect 193926 316046 193982 316102
rect 193554 315922 193610 315978
rect 193678 315922 193734 315978
rect 193802 315922 193858 315978
rect 193926 315922 193982 315978
rect 194518 310294 194574 310350
rect 194642 310294 194698 310350
rect 194518 310170 194574 310226
rect 194642 310170 194698 310226
rect 194518 310046 194574 310102
rect 194642 310046 194698 310102
rect 194518 309922 194574 309978
rect 194642 309922 194698 309978
rect 193554 298294 193610 298350
rect 193678 298294 193734 298350
rect 193802 298294 193858 298350
rect 193926 298294 193982 298350
rect 193554 298170 193610 298226
rect 193678 298170 193734 298226
rect 193802 298170 193858 298226
rect 193926 298170 193982 298226
rect 193554 298046 193610 298102
rect 193678 298046 193734 298102
rect 193802 298046 193858 298102
rect 193926 298046 193982 298102
rect 193554 297922 193610 297978
rect 193678 297922 193734 297978
rect 193802 297922 193858 297978
rect 193926 297922 193982 297978
rect 194518 292294 194574 292350
rect 194642 292294 194698 292350
rect 194518 292170 194574 292226
rect 194642 292170 194698 292226
rect 194518 292046 194574 292102
rect 194642 292046 194698 292102
rect 194518 291922 194574 291978
rect 194642 291922 194698 291978
rect 193554 280294 193610 280350
rect 193678 280294 193734 280350
rect 193802 280294 193858 280350
rect 193926 280294 193982 280350
rect 193554 280170 193610 280226
rect 193678 280170 193734 280226
rect 193802 280170 193858 280226
rect 193926 280170 193982 280226
rect 193554 280046 193610 280102
rect 193678 280046 193734 280102
rect 193802 280046 193858 280102
rect 193926 280046 193982 280102
rect 193554 279922 193610 279978
rect 193678 279922 193734 279978
rect 193802 279922 193858 279978
rect 193926 279922 193982 279978
rect 194518 274294 194574 274350
rect 194642 274294 194698 274350
rect 194518 274170 194574 274226
rect 194642 274170 194698 274226
rect 194518 274046 194574 274102
rect 194642 274046 194698 274102
rect 194518 273922 194574 273978
rect 194642 273922 194698 273978
rect 193554 262294 193610 262350
rect 193678 262294 193734 262350
rect 193802 262294 193858 262350
rect 193926 262294 193982 262350
rect 193554 262170 193610 262226
rect 193678 262170 193734 262226
rect 193802 262170 193858 262226
rect 193926 262170 193982 262226
rect 193554 262046 193610 262102
rect 193678 262046 193734 262102
rect 193802 262046 193858 262102
rect 193926 262046 193982 262102
rect 193554 261922 193610 261978
rect 193678 261922 193734 261978
rect 193802 261922 193858 261978
rect 193926 261922 193982 261978
rect 194518 256294 194574 256350
rect 194642 256294 194698 256350
rect 194518 256170 194574 256226
rect 194642 256170 194698 256226
rect 194518 256046 194574 256102
rect 194642 256046 194698 256102
rect 194518 255922 194574 255978
rect 194642 255922 194698 255978
rect 193554 244294 193610 244350
rect 193678 244294 193734 244350
rect 193802 244294 193858 244350
rect 193926 244294 193982 244350
rect 193554 244170 193610 244226
rect 193678 244170 193734 244226
rect 193802 244170 193858 244226
rect 193926 244170 193982 244226
rect 193554 244046 193610 244102
rect 193678 244046 193734 244102
rect 193802 244046 193858 244102
rect 193926 244046 193982 244102
rect 193554 243922 193610 243978
rect 193678 243922 193734 243978
rect 193802 243922 193858 243978
rect 193926 243922 193982 243978
rect 193554 226294 193610 226350
rect 193678 226294 193734 226350
rect 193802 226294 193858 226350
rect 193926 226294 193982 226350
rect 193554 226170 193610 226226
rect 193678 226170 193734 226226
rect 193802 226170 193858 226226
rect 193926 226170 193982 226226
rect 193554 226046 193610 226102
rect 193678 226046 193734 226102
rect 193802 226046 193858 226102
rect 193926 226046 193982 226102
rect 193554 225922 193610 225978
rect 193678 225922 193734 225978
rect 193802 225922 193858 225978
rect 193926 225922 193982 225978
rect 194236 248642 194292 248698
rect 199836 401642 199892 401698
rect 199724 393542 199780 393598
rect 199388 373742 199444 373798
rect 197596 340082 197652 340138
rect 199276 368702 199332 368758
rect 197484 287162 197540 287218
rect 197596 288962 197652 289018
rect 197484 281402 197540 281458
rect 197708 285722 197764 285778
rect 198044 268802 198100 268858
rect 197820 249722 197876 249778
rect 196476 211382 196532 211438
rect 197932 247202 197988 247258
rect 197932 214262 197988 214318
rect 201516 393362 201572 393418
rect 201404 391922 201460 391978
rect 204876 392102 204932 392158
rect 220554 400294 220610 400350
rect 220678 400294 220734 400350
rect 220802 400294 220858 400350
rect 220926 400294 220982 400350
rect 220554 400170 220610 400226
rect 220678 400170 220734 400226
rect 220802 400170 220858 400226
rect 220926 400170 220982 400226
rect 220554 400046 220610 400102
rect 220678 400046 220734 400102
rect 220802 400046 220858 400102
rect 220926 400046 220982 400102
rect 220554 399922 220610 399978
rect 220678 399922 220734 399978
rect 220802 399922 220858 399978
rect 220926 399922 220982 399978
rect 215068 391382 215124 391438
rect 216636 391412 216692 391438
rect 216636 391382 216692 391412
rect 220554 382294 220610 382350
rect 220678 382294 220734 382350
rect 220802 382294 220858 382350
rect 220926 382294 220982 382350
rect 220554 382170 220610 382226
rect 220678 382170 220734 382226
rect 220802 382170 220858 382226
rect 220926 382170 220982 382226
rect 220554 382046 220610 382102
rect 220678 382046 220734 382102
rect 220802 382046 220858 382102
rect 220926 382046 220982 382102
rect 220554 381922 220610 381978
rect 220678 381922 220734 381978
rect 220802 381922 220858 381978
rect 220926 381922 220982 381978
rect 209878 370294 209934 370350
rect 210002 370294 210058 370350
rect 209878 370170 209934 370226
rect 210002 370170 210058 370226
rect 209878 370046 209934 370102
rect 210002 370046 210058 370102
rect 209878 369922 209934 369978
rect 210002 369922 210058 369978
rect 243516 407582 243572 407638
rect 248892 406862 248948 406918
rect 224274 406294 224330 406350
rect 224398 406294 224454 406350
rect 224522 406294 224578 406350
rect 224646 406294 224702 406350
rect 224274 406170 224330 406226
rect 224398 406170 224454 406226
rect 224522 406170 224578 406226
rect 224646 406170 224702 406226
rect 224274 406046 224330 406102
rect 224398 406046 224454 406102
rect 224522 406046 224578 406102
rect 224646 406046 224702 406102
rect 224274 405922 224330 405978
rect 224398 405922 224454 405978
rect 224522 405922 224578 405978
rect 224646 405922 224702 405978
rect 227612 406682 227668 406738
rect 251274 400294 251330 400350
rect 251398 400294 251454 400350
rect 251522 400294 251578 400350
rect 251646 400294 251702 400350
rect 251274 400170 251330 400226
rect 251398 400170 251454 400226
rect 251522 400170 251578 400226
rect 251646 400170 251702 400226
rect 251274 400046 251330 400102
rect 251398 400046 251454 400102
rect 251522 400046 251578 400102
rect 251646 400046 251702 400102
rect 251274 399922 251330 399978
rect 251398 399922 251454 399978
rect 251522 399922 251578 399978
rect 251646 399922 251702 399978
rect 231644 395162 231700 395218
rect 224274 388294 224330 388350
rect 224398 388294 224454 388350
rect 224522 388294 224578 388350
rect 224646 388294 224702 388350
rect 224274 388170 224330 388226
rect 224398 388170 224454 388226
rect 224522 388170 224578 388226
rect 224646 388170 224702 388226
rect 224274 388046 224330 388102
rect 224398 388046 224454 388102
rect 224522 388046 224578 388102
rect 224646 388046 224702 388102
rect 224274 387922 224330 387978
rect 224398 387922 224454 387978
rect 224522 387922 224578 387978
rect 224646 387922 224702 387978
rect 230076 393722 230132 393778
rect 231756 394982 231812 395038
rect 251274 382294 251330 382350
rect 251398 382294 251454 382350
rect 251522 382294 251578 382350
rect 251646 382294 251702 382350
rect 251274 382170 251330 382226
rect 251398 382170 251454 382226
rect 251522 382170 251578 382226
rect 251646 382170 251702 382226
rect 251274 382046 251330 382102
rect 251398 382046 251454 382102
rect 251522 382046 251578 382102
rect 251646 382046 251702 382102
rect 251274 381922 251330 381978
rect 251398 381922 251454 381978
rect 251522 381922 251578 381978
rect 251646 381922 251702 381978
rect 236124 379708 236180 379738
rect 236124 379682 236180 379708
rect 224274 370294 224330 370350
rect 224398 370294 224454 370350
rect 224522 370294 224578 370350
rect 224646 370294 224702 370350
rect 224274 370170 224330 370226
rect 224398 370170 224454 370226
rect 224522 370170 224578 370226
rect 224646 370170 224702 370226
rect 224274 370046 224330 370102
rect 224398 370046 224454 370102
rect 224522 370046 224578 370102
rect 224646 370046 224702 370102
rect 224274 369922 224330 369978
rect 224398 369922 224454 369978
rect 224522 369922 224578 369978
rect 224646 369922 224702 369978
rect 237020 373742 237076 373798
rect 235228 368702 235284 368758
rect 240598 370294 240654 370350
rect 240722 370294 240778 370350
rect 240598 370170 240654 370226
rect 240722 370170 240778 370226
rect 240598 370046 240654 370102
rect 240722 370046 240778 370102
rect 240598 369922 240654 369978
rect 240722 369922 240778 369978
rect 238476 368702 238532 368758
rect 277116 407402 277172 407458
rect 254994 406294 255050 406350
rect 255118 406294 255174 406350
rect 255242 406294 255298 406350
rect 255366 406294 255422 406350
rect 254994 406170 255050 406226
rect 255118 406170 255174 406226
rect 255242 406170 255298 406226
rect 255366 406170 255422 406226
rect 254994 406046 255050 406102
rect 255118 406046 255174 406102
rect 255242 406046 255298 406102
rect 255366 406046 255422 406102
rect 254994 405922 255050 405978
rect 255118 405922 255174 405978
rect 255242 405922 255298 405978
rect 255366 405922 255422 405978
rect 254994 388294 255050 388350
rect 255118 388294 255174 388350
rect 255242 388294 255298 388350
rect 255366 388294 255422 388350
rect 254994 388170 255050 388226
rect 255118 388170 255174 388226
rect 255242 388170 255298 388226
rect 255366 388170 255422 388226
rect 254994 388046 255050 388102
rect 255118 388046 255174 388102
rect 255242 388046 255298 388102
rect 255366 388046 255422 388102
rect 254994 387922 255050 387978
rect 255118 387922 255174 387978
rect 255242 387922 255298 387978
rect 255366 387922 255422 387978
rect 254994 370294 255050 370350
rect 255118 370294 255174 370350
rect 255242 370294 255298 370350
rect 255366 370294 255422 370350
rect 254994 370170 255050 370226
rect 255118 370170 255174 370226
rect 255242 370170 255298 370226
rect 255366 370170 255422 370226
rect 254994 370046 255050 370102
rect 255118 370046 255174 370102
rect 255242 370046 255298 370102
rect 255366 370046 255422 370102
rect 254994 369922 255050 369978
rect 255118 369922 255174 369978
rect 255242 369922 255298 369978
rect 255366 369922 255422 369978
rect 266252 368882 266308 368938
rect 281372 373742 281428 373798
rect 281994 400294 282050 400350
rect 282118 400294 282174 400350
rect 282242 400294 282298 400350
rect 282366 400294 282422 400350
rect 281994 400170 282050 400226
rect 282118 400170 282174 400226
rect 282242 400170 282298 400226
rect 282366 400170 282422 400226
rect 281994 400046 282050 400102
rect 282118 400046 282174 400102
rect 282242 400046 282298 400102
rect 282366 400046 282422 400102
rect 281994 399922 282050 399978
rect 282118 399922 282174 399978
rect 282242 399922 282298 399978
rect 282366 399922 282422 399978
rect 281994 382294 282050 382350
rect 282118 382294 282174 382350
rect 282242 382294 282298 382350
rect 282366 382294 282422 382350
rect 281994 382170 282050 382226
rect 282118 382170 282174 382226
rect 282242 382170 282298 382226
rect 282366 382170 282422 382226
rect 281994 382046 282050 382102
rect 282118 382046 282174 382102
rect 282242 382046 282298 382102
rect 282366 382046 282422 382102
rect 281994 381922 282050 381978
rect 282118 381922 282174 381978
rect 282242 381922 282298 381978
rect 282366 381922 282422 381978
rect 276332 373022 276388 373078
rect 271318 370294 271374 370350
rect 271442 370294 271498 370350
rect 271318 370170 271374 370226
rect 271442 370170 271498 370226
rect 271318 370046 271374 370102
rect 271442 370046 271498 370102
rect 271318 369922 271374 369978
rect 271442 369922 271498 369978
rect 285714 406294 285770 406350
rect 285838 406294 285894 406350
rect 285962 406294 286018 406350
rect 286086 406294 286142 406350
rect 285714 406170 285770 406226
rect 285838 406170 285894 406226
rect 285962 406170 286018 406226
rect 286086 406170 286142 406226
rect 285714 406046 285770 406102
rect 285838 406046 285894 406102
rect 285962 406046 286018 406102
rect 286086 406046 286142 406102
rect 285714 405922 285770 405978
rect 285838 405922 285894 405978
rect 285962 405922 286018 405978
rect 286086 405922 286142 405978
rect 285714 388294 285770 388350
rect 285838 388294 285894 388350
rect 285962 388294 286018 388350
rect 286086 388294 286142 388350
rect 285714 388170 285770 388226
rect 285838 388170 285894 388226
rect 285962 388170 286018 388226
rect 286086 388170 286142 388226
rect 285714 388046 285770 388102
rect 285838 388046 285894 388102
rect 285962 388046 286018 388102
rect 286086 388046 286142 388102
rect 285714 387922 285770 387978
rect 285838 387922 285894 387978
rect 285962 387922 286018 387978
rect 286086 387922 286142 387978
rect 312714 400294 312770 400350
rect 312838 400294 312894 400350
rect 312962 400294 313018 400350
rect 313086 400294 313142 400350
rect 312714 400170 312770 400226
rect 312838 400170 312894 400226
rect 312962 400170 313018 400226
rect 313086 400170 313142 400226
rect 312714 400046 312770 400102
rect 312838 400046 312894 400102
rect 312962 400046 313018 400102
rect 313086 400046 313142 400102
rect 312714 399922 312770 399978
rect 312838 399922 312894 399978
rect 312962 399922 313018 399978
rect 313086 399922 313142 399978
rect 307356 399122 307412 399178
rect 305676 398942 305732 398998
rect 312714 382294 312770 382350
rect 312838 382294 312894 382350
rect 312962 382294 313018 382350
rect 313086 382294 313142 382350
rect 312714 382170 312770 382226
rect 312838 382170 312894 382226
rect 312962 382170 313018 382226
rect 313086 382170 313142 382226
rect 286412 372122 286468 372178
rect 312714 382046 312770 382102
rect 312838 382046 312894 382102
rect 312962 382046 313018 382102
rect 313086 382046 313142 382102
rect 312714 381922 312770 381978
rect 312838 381922 312894 381978
rect 312962 381922 313018 381978
rect 313086 381922 313142 381978
rect 285714 370294 285770 370350
rect 285838 370294 285894 370350
rect 285962 370294 286018 370350
rect 286086 370294 286142 370350
rect 285714 370170 285770 370226
rect 285838 370170 285894 370226
rect 285962 370170 286018 370226
rect 286086 370170 286142 370226
rect 285714 370046 285770 370102
rect 285838 370046 285894 370102
rect 285962 370046 286018 370102
rect 286086 370046 286142 370102
rect 285714 369922 285770 369978
rect 285838 369922 285894 369978
rect 285962 369922 286018 369978
rect 286086 369922 286142 369978
rect 302038 370294 302094 370350
rect 302162 370294 302218 370350
rect 302038 370170 302094 370226
rect 302162 370170 302218 370226
rect 302038 370046 302094 370102
rect 302162 370046 302218 370102
rect 302038 369922 302094 369978
rect 302162 369922 302218 369978
rect 316434 406294 316490 406350
rect 316558 406294 316614 406350
rect 316682 406294 316738 406350
rect 316806 406294 316862 406350
rect 316434 406170 316490 406226
rect 316558 406170 316614 406226
rect 316682 406170 316738 406226
rect 316806 406170 316862 406226
rect 316434 406046 316490 406102
rect 316558 406046 316614 406102
rect 316682 406046 316738 406102
rect 316806 406046 316862 406102
rect 316434 405922 316490 405978
rect 316558 405922 316614 405978
rect 316682 405922 316738 405978
rect 316806 405922 316862 405978
rect 316434 388294 316490 388350
rect 316558 388294 316614 388350
rect 316682 388294 316738 388350
rect 316806 388294 316862 388350
rect 316434 388170 316490 388226
rect 316558 388170 316614 388226
rect 316682 388170 316738 388226
rect 316806 388170 316862 388226
rect 316434 388046 316490 388102
rect 316558 388046 316614 388102
rect 316682 388046 316738 388102
rect 316806 388046 316862 388102
rect 316434 387922 316490 387978
rect 316558 387922 316614 387978
rect 316682 387922 316738 387978
rect 316806 387922 316862 387978
rect 319116 400562 319172 400618
rect 320796 399302 320852 399358
rect 329196 409202 329252 409258
rect 323372 376262 323428 376318
rect 316434 370294 316490 370350
rect 316558 370294 316614 370350
rect 316682 370294 316738 370350
rect 316806 370294 316862 370350
rect 316434 370170 316490 370226
rect 316558 370170 316614 370226
rect 316682 370170 316738 370226
rect 316806 370170 316862 370226
rect 316434 370046 316490 370102
rect 316558 370046 316614 370102
rect 316682 370046 316738 370102
rect 316806 370046 316862 370102
rect 316434 369922 316490 369978
rect 316558 369922 316614 369978
rect 316682 369922 316738 369978
rect 316806 369922 316862 369978
rect 330876 405602 330932 405658
rect 332758 370294 332814 370350
rect 332882 370294 332938 370350
rect 332758 370170 332814 370226
rect 332882 370170 332938 370226
rect 332758 370046 332814 370102
rect 332882 370046 332938 370102
rect 332758 369922 332814 369978
rect 332882 369922 332938 369978
rect 329084 369062 329140 369118
rect 276332 367082 276388 367138
rect 270508 365822 270564 365878
rect 272076 366542 272132 366598
rect 272076 365822 272132 365878
rect 225238 364294 225294 364350
rect 225362 364294 225418 364350
rect 225238 364170 225294 364226
rect 225362 364170 225418 364226
rect 225238 364046 225294 364102
rect 225362 364046 225418 364102
rect 225238 363922 225294 363978
rect 225362 363922 225418 363978
rect 255958 364294 256014 364350
rect 256082 364294 256138 364350
rect 255958 364170 256014 364226
rect 256082 364170 256138 364226
rect 255958 364046 256014 364102
rect 256082 364046 256138 364102
rect 255958 363922 256014 363978
rect 256082 363922 256138 363978
rect 286678 364294 286734 364350
rect 286802 364294 286858 364350
rect 286678 364170 286734 364226
rect 286802 364170 286858 364226
rect 286678 364046 286734 364102
rect 286802 364046 286858 364102
rect 286678 363922 286734 363978
rect 286802 363922 286858 363978
rect 317398 364294 317454 364350
rect 317522 364294 317578 364350
rect 317398 364170 317454 364226
rect 317522 364170 317578 364226
rect 317398 364046 317454 364102
rect 317522 364046 317578 364102
rect 317398 363922 317454 363978
rect 317522 363922 317578 363978
rect 335916 356102 335972 356158
rect 336028 368702 336084 368758
rect 209878 352294 209934 352350
rect 210002 352294 210058 352350
rect 209878 352170 209934 352226
rect 210002 352170 210058 352226
rect 209878 352046 209934 352102
rect 210002 352046 210058 352102
rect 209878 351922 209934 351978
rect 210002 351922 210058 351978
rect 240598 352294 240654 352350
rect 240722 352294 240778 352350
rect 240598 352170 240654 352226
rect 240722 352170 240778 352226
rect 240598 352046 240654 352102
rect 240722 352046 240778 352102
rect 240598 351922 240654 351978
rect 240722 351922 240778 351978
rect 271318 352294 271374 352350
rect 271442 352294 271498 352350
rect 271318 352170 271374 352226
rect 271442 352170 271498 352226
rect 271318 352046 271374 352102
rect 271442 352046 271498 352102
rect 271318 351922 271374 351978
rect 271442 351922 271498 351978
rect 302038 352294 302094 352350
rect 302162 352294 302218 352350
rect 302038 352170 302094 352226
rect 302162 352170 302218 352226
rect 302038 352046 302094 352102
rect 302162 352046 302218 352102
rect 302038 351922 302094 351978
rect 302162 351922 302218 351978
rect 332758 352294 332814 352350
rect 332882 352294 332938 352350
rect 332758 352170 332814 352226
rect 332882 352170 332938 352226
rect 332758 352046 332814 352102
rect 332882 352046 332938 352102
rect 332758 351922 332814 351978
rect 332882 351922 332938 351978
rect 225238 346294 225294 346350
rect 225362 346294 225418 346350
rect 225238 346170 225294 346226
rect 225362 346170 225418 346226
rect 225238 346046 225294 346102
rect 225362 346046 225418 346102
rect 225238 345922 225294 345978
rect 225362 345922 225418 345978
rect 255958 346294 256014 346350
rect 256082 346294 256138 346350
rect 255958 346170 256014 346226
rect 256082 346170 256138 346226
rect 255958 346046 256014 346102
rect 256082 346046 256138 346102
rect 255958 345922 256014 345978
rect 256082 345922 256138 345978
rect 286678 346294 286734 346350
rect 286802 346294 286858 346350
rect 286678 346170 286734 346226
rect 286802 346170 286858 346226
rect 286678 346046 286734 346102
rect 286802 346046 286858 346102
rect 286678 345922 286734 345978
rect 286802 345922 286858 345978
rect 317398 346294 317454 346350
rect 317522 346294 317578 346350
rect 317398 346170 317454 346226
rect 317522 346170 317578 346226
rect 317398 346046 317454 346102
rect 317522 346046 317578 346102
rect 317398 345922 317454 345978
rect 317522 345922 317578 345978
rect 209878 334294 209934 334350
rect 210002 334294 210058 334350
rect 209878 334170 209934 334226
rect 210002 334170 210058 334226
rect 209878 334046 209934 334102
rect 210002 334046 210058 334102
rect 209878 333922 209934 333978
rect 210002 333922 210058 333978
rect 240598 334294 240654 334350
rect 240722 334294 240778 334350
rect 240598 334170 240654 334226
rect 240722 334170 240778 334226
rect 240598 334046 240654 334102
rect 240722 334046 240778 334102
rect 240598 333922 240654 333978
rect 240722 333922 240778 333978
rect 271318 334294 271374 334350
rect 271442 334294 271498 334350
rect 271318 334170 271374 334226
rect 271442 334170 271498 334226
rect 271318 334046 271374 334102
rect 271442 334046 271498 334102
rect 271318 333922 271374 333978
rect 271442 333922 271498 333978
rect 302038 334294 302094 334350
rect 302162 334294 302218 334350
rect 302038 334170 302094 334226
rect 302162 334170 302218 334226
rect 302038 334046 302094 334102
rect 302162 334046 302218 334102
rect 302038 333922 302094 333978
rect 302162 333922 302218 333978
rect 332758 334294 332814 334350
rect 332882 334294 332938 334350
rect 332758 334170 332814 334226
rect 332882 334170 332938 334226
rect 332758 334046 332814 334102
rect 332882 334046 332938 334102
rect 332758 333922 332814 333978
rect 332882 333922 332938 333978
rect 225238 328294 225294 328350
rect 225362 328294 225418 328350
rect 225238 328170 225294 328226
rect 225362 328170 225418 328226
rect 225238 328046 225294 328102
rect 225362 328046 225418 328102
rect 225238 327922 225294 327978
rect 225362 327922 225418 327978
rect 255958 328294 256014 328350
rect 256082 328294 256138 328350
rect 255958 328170 256014 328226
rect 256082 328170 256138 328226
rect 255958 328046 256014 328102
rect 256082 328046 256138 328102
rect 255958 327922 256014 327978
rect 256082 327922 256138 327978
rect 286678 328294 286734 328350
rect 286802 328294 286858 328350
rect 286678 328170 286734 328226
rect 286802 328170 286858 328226
rect 286678 328046 286734 328102
rect 286802 328046 286858 328102
rect 286678 327922 286734 327978
rect 286802 327922 286858 327978
rect 317398 328294 317454 328350
rect 317522 328294 317578 328350
rect 317398 328170 317454 328226
rect 317522 328170 317578 328226
rect 317398 328046 317454 328102
rect 317522 328046 317578 328102
rect 317398 327922 317454 327978
rect 317522 327922 317578 327978
rect 209878 316294 209934 316350
rect 210002 316294 210058 316350
rect 209878 316170 209934 316226
rect 210002 316170 210058 316226
rect 209878 316046 209934 316102
rect 210002 316046 210058 316102
rect 209878 315922 209934 315978
rect 210002 315922 210058 315978
rect 240598 316294 240654 316350
rect 240722 316294 240778 316350
rect 240598 316170 240654 316226
rect 240722 316170 240778 316226
rect 240598 316046 240654 316102
rect 240722 316046 240778 316102
rect 240598 315922 240654 315978
rect 240722 315922 240778 315978
rect 271318 316294 271374 316350
rect 271442 316294 271498 316350
rect 271318 316170 271374 316226
rect 271442 316170 271498 316226
rect 271318 316046 271374 316102
rect 271442 316046 271498 316102
rect 271318 315922 271374 315978
rect 271442 315922 271498 315978
rect 302038 316294 302094 316350
rect 302162 316294 302218 316350
rect 302038 316170 302094 316226
rect 302162 316170 302218 316226
rect 302038 316046 302094 316102
rect 302162 316046 302218 316102
rect 302038 315922 302094 315978
rect 302162 315922 302218 315978
rect 332758 316294 332814 316350
rect 332882 316294 332938 316350
rect 332758 316170 332814 316226
rect 332882 316170 332938 316226
rect 332758 316046 332814 316102
rect 332882 316046 332938 316102
rect 332758 315922 332814 315978
rect 332882 315922 332938 315978
rect 225238 310294 225294 310350
rect 225362 310294 225418 310350
rect 225238 310170 225294 310226
rect 225362 310170 225418 310226
rect 225238 310046 225294 310102
rect 225362 310046 225418 310102
rect 225238 309922 225294 309978
rect 225362 309922 225418 309978
rect 255958 310294 256014 310350
rect 256082 310294 256138 310350
rect 255958 310170 256014 310226
rect 256082 310170 256138 310226
rect 255958 310046 256014 310102
rect 256082 310046 256138 310102
rect 255958 309922 256014 309978
rect 256082 309922 256138 309978
rect 286678 310294 286734 310350
rect 286802 310294 286858 310350
rect 286678 310170 286734 310226
rect 286802 310170 286858 310226
rect 286678 310046 286734 310102
rect 286802 310046 286858 310102
rect 286678 309922 286734 309978
rect 286802 309922 286858 309978
rect 317398 310294 317454 310350
rect 317522 310294 317578 310350
rect 317398 310170 317454 310226
rect 317522 310170 317578 310226
rect 317398 310046 317454 310102
rect 317522 310046 317578 310102
rect 317398 309922 317454 309978
rect 317522 309922 317578 309978
rect 209878 298294 209934 298350
rect 210002 298294 210058 298350
rect 209878 298170 209934 298226
rect 210002 298170 210058 298226
rect 209878 298046 209934 298102
rect 210002 298046 210058 298102
rect 209878 297922 209934 297978
rect 210002 297922 210058 297978
rect 240598 298294 240654 298350
rect 240722 298294 240778 298350
rect 240598 298170 240654 298226
rect 240722 298170 240778 298226
rect 240598 298046 240654 298102
rect 240722 298046 240778 298102
rect 240598 297922 240654 297978
rect 240722 297922 240778 297978
rect 271318 298294 271374 298350
rect 271442 298294 271498 298350
rect 271318 298170 271374 298226
rect 271442 298170 271498 298226
rect 271318 298046 271374 298102
rect 271442 298046 271498 298102
rect 271318 297922 271374 297978
rect 271442 297922 271498 297978
rect 302038 298294 302094 298350
rect 302162 298294 302218 298350
rect 302038 298170 302094 298226
rect 302162 298170 302218 298226
rect 302038 298046 302094 298102
rect 302162 298046 302218 298102
rect 302038 297922 302094 297978
rect 302162 297922 302218 297978
rect 332758 298294 332814 298350
rect 332882 298294 332938 298350
rect 332758 298170 332814 298226
rect 332882 298170 332938 298226
rect 332758 298046 332814 298102
rect 332882 298046 332938 298102
rect 332758 297922 332814 297978
rect 332882 297922 332938 297978
rect 225238 292294 225294 292350
rect 225362 292294 225418 292350
rect 225238 292170 225294 292226
rect 225362 292170 225418 292226
rect 225238 292046 225294 292102
rect 225362 292046 225418 292102
rect 225238 291922 225294 291978
rect 225362 291922 225418 291978
rect 255958 292294 256014 292350
rect 256082 292294 256138 292350
rect 255958 292170 256014 292226
rect 256082 292170 256138 292226
rect 255958 292046 256014 292102
rect 256082 292046 256138 292102
rect 255958 291922 256014 291978
rect 256082 291922 256138 291978
rect 286678 292294 286734 292350
rect 286802 292294 286858 292350
rect 286678 292170 286734 292226
rect 286802 292170 286858 292226
rect 286678 292046 286734 292102
rect 286802 292046 286858 292102
rect 286678 291922 286734 291978
rect 286802 291922 286858 291978
rect 317398 292294 317454 292350
rect 317522 292294 317578 292350
rect 317398 292170 317454 292226
rect 317522 292170 317578 292226
rect 317398 292046 317454 292102
rect 317522 292046 317578 292102
rect 317398 291922 317454 291978
rect 317522 291922 317578 291978
rect 209878 280294 209934 280350
rect 210002 280294 210058 280350
rect 209878 280170 209934 280226
rect 210002 280170 210058 280226
rect 209878 280046 209934 280102
rect 210002 280046 210058 280102
rect 209878 279922 209934 279978
rect 210002 279922 210058 279978
rect 240598 280294 240654 280350
rect 240722 280294 240778 280350
rect 240598 280170 240654 280226
rect 240722 280170 240778 280226
rect 240598 280046 240654 280102
rect 240722 280046 240778 280102
rect 240598 279922 240654 279978
rect 240722 279922 240778 279978
rect 271318 280294 271374 280350
rect 271442 280294 271498 280350
rect 271318 280170 271374 280226
rect 271442 280170 271498 280226
rect 271318 280046 271374 280102
rect 271442 280046 271498 280102
rect 271318 279922 271374 279978
rect 271442 279922 271498 279978
rect 302038 280294 302094 280350
rect 302162 280294 302218 280350
rect 302038 280170 302094 280226
rect 302162 280170 302218 280226
rect 302038 280046 302094 280102
rect 302162 280046 302218 280102
rect 302038 279922 302094 279978
rect 302162 279922 302218 279978
rect 332758 280294 332814 280350
rect 332882 280294 332938 280350
rect 332758 280170 332814 280226
rect 332882 280170 332938 280226
rect 332758 280046 332814 280102
rect 332882 280046 332938 280102
rect 332758 279922 332814 279978
rect 332882 279922 332938 279978
rect 225238 274294 225294 274350
rect 225362 274294 225418 274350
rect 225238 274170 225294 274226
rect 225362 274170 225418 274226
rect 225238 274046 225294 274102
rect 225362 274046 225418 274102
rect 225238 273922 225294 273978
rect 225362 273922 225418 273978
rect 255958 274294 256014 274350
rect 256082 274294 256138 274350
rect 255958 274170 256014 274226
rect 256082 274170 256138 274226
rect 255958 274046 256014 274102
rect 256082 274046 256138 274102
rect 255958 273922 256014 273978
rect 256082 273922 256138 273978
rect 286678 274294 286734 274350
rect 286802 274294 286858 274350
rect 286678 274170 286734 274226
rect 286802 274170 286858 274226
rect 286678 274046 286734 274102
rect 286802 274046 286858 274102
rect 286678 273922 286734 273978
rect 286802 273922 286858 273978
rect 317398 274294 317454 274350
rect 317522 274294 317578 274350
rect 317398 274170 317454 274226
rect 317522 274170 317578 274226
rect 317398 274046 317454 274102
rect 317522 274046 317578 274102
rect 317398 273922 317454 273978
rect 317522 273922 317578 273978
rect 209878 262294 209934 262350
rect 210002 262294 210058 262350
rect 209878 262170 209934 262226
rect 210002 262170 210058 262226
rect 209878 262046 209934 262102
rect 210002 262046 210058 262102
rect 209878 261922 209934 261978
rect 210002 261922 210058 261978
rect 240598 262294 240654 262350
rect 240722 262294 240778 262350
rect 240598 262170 240654 262226
rect 240722 262170 240778 262226
rect 240598 262046 240654 262102
rect 240722 262046 240778 262102
rect 240598 261922 240654 261978
rect 240722 261922 240778 261978
rect 271318 262294 271374 262350
rect 271442 262294 271498 262350
rect 271318 262170 271374 262226
rect 271442 262170 271498 262226
rect 271318 262046 271374 262102
rect 271442 262046 271498 262102
rect 271318 261922 271374 261978
rect 271442 261922 271498 261978
rect 302038 262294 302094 262350
rect 302162 262294 302218 262350
rect 302038 262170 302094 262226
rect 302162 262170 302218 262226
rect 302038 262046 302094 262102
rect 302162 262046 302218 262102
rect 302038 261922 302094 261978
rect 302162 261922 302218 261978
rect 332758 262294 332814 262350
rect 332882 262294 332938 262350
rect 332758 262170 332814 262226
rect 332882 262170 332938 262226
rect 332758 262046 332814 262102
rect 332882 262046 332938 262102
rect 332758 261922 332814 261978
rect 332882 261922 332938 261978
rect 225238 256294 225294 256350
rect 225362 256294 225418 256350
rect 225238 256170 225294 256226
rect 225362 256170 225418 256226
rect 225238 256046 225294 256102
rect 225362 256046 225418 256102
rect 225238 255922 225294 255978
rect 225362 255922 225418 255978
rect 255958 256294 256014 256350
rect 256082 256294 256138 256350
rect 255958 256170 256014 256226
rect 256082 256170 256138 256226
rect 255958 256046 256014 256102
rect 256082 256046 256138 256102
rect 255958 255922 256014 255978
rect 256082 255922 256138 255978
rect 286678 256294 286734 256350
rect 286802 256294 286858 256350
rect 286678 256170 286734 256226
rect 286802 256170 286858 256226
rect 286678 256046 286734 256102
rect 286802 256046 286858 256102
rect 286678 255922 286734 255978
rect 286802 255922 286858 255978
rect 317398 256294 317454 256350
rect 317522 256294 317578 256350
rect 317398 256170 317454 256226
rect 317522 256170 317578 256226
rect 317398 256046 317454 256102
rect 317522 256046 317578 256102
rect 317398 255922 317454 255978
rect 317522 255922 317578 255978
rect 335804 253502 335860 253558
rect 209878 244294 209934 244350
rect 210002 244294 210058 244350
rect 209878 244170 209934 244226
rect 210002 244170 210058 244226
rect 209878 244046 209934 244102
rect 210002 244046 210058 244102
rect 209878 243922 209934 243978
rect 210002 243922 210058 243978
rect 240598 244294 240654 244350
rect 240722 244294 240778 244350
rect 240598 244170 240654 244226
rect 240722 244170 240778 244226
rect 240598 244046 240654 244102
rect 240722 244046 240778 244102
rect 240598 243922 240654 243978
rect 240722 243922 240778 243978
rect 271318 244294 271374 244350
rect 271442 244294 271498 244350
rect 271318 244170 271374 244226
rect 271442 244170 271498 244226
rect 271318 244046 271374 244102
rect 271442 244046 271498 244102
rect 271318 243922 271374 243978
rect 271442 243922 271498 243978
rect 302038 244294 302094 244350
rect 302162 244294 302218 244350
rect 302038 244170 302094 244226
rect 302162 244170 302218 244226
rect 302038 244046 302094 244102
rect 302162 244046 302218 244102
rect 302038 243922 302094 243978
rect 302162 243922 302218 243978
rect 332758 244294 332814 244350
rect 332882 244294 332938 244350
rect 332758 244170 332814 244226
rect 332882 244170 332938 244226
rect 332758 244046 332814 244102
rect 332882 244046 332938 244102
rect 332758 243922 332814 243978
rect 332882 243922 332938 243978
rect 323260 242702 323316 242758
rect 278012 241982 278068 242038
rect 220554 238294 220610 238350
rect 220678 238294 220734 238350
rect 220802 238294 220858 238350
rect 220926 238294 220982 238350
rect 220554 238170 220610 238226
rect 220678 238170 220734 238226
rect 220802 238170 220858 238226
rect 220926 238170 220982 238226
rect 220554 238046 220610 238102
rect 220678 238046 220734 238102
rect 220802 238046 220858 238102
rect 220926 238046 220982 238102
rect 220554 237922 220610 237978
rect 220678 237922 220734 237978
rect 220802 237922 220858 237978
rect 220926 237922 220982 237978
rect 219996 231362 220052 231418
rect 218316 231182 218372 231238
rect 233212 234422 233268 234478
rect 242620 237122 242676 237178
rect 251274 238294 251330 238350
rect 251398 238294 251454 238350
rect 251522 238294 251578 238350
rect 251646 238294 251702 238350
rect 251274 238170 251330 238226
rect 251398 238170 251454 238226
rect 251522 238170 251578 238226
rect 251646 238170 251702 238226
rect 251274 238046 251330 238102
rect 251398 238046 251454 238102
rect 251522 238046 251578 238102
rect 251646 238046 251702 238102
rect 251274 237922 251330 237978
rect 251398 237922 251454 237978
rect 251522 237922 251578 237978
rect 251646 237922 251702 237978
rect 235900 234422 235956 234478
rect 241948 236942 242004 236998
rect 228508 231002 228564 231058
rect 236796 227762 236852 227818
rect 220554 220294 220610 220350
rect 220678 220294 220734 220350
rect 220802 220294 220858 220350
rect 220926 220294 220982 220350
rect 220554 220170 220610 220226
rect 220678 220170 220734 220226
rect 220802 220170 220858 220226
rect 220926 220170 220982 220226
rect 220554 220046 220610 220102
rect 220678 220046 220734 220102
rect 220802 220046 220858 220102
rect 220926 220046 220982 220102
rect 220554 219922 220610 219978
rect 220678 219922 220734 219978
rect 220802 219922 220858 219978
rect 220926 219922 220982 219978
rect 199276 211202 199332 211258
rect 197820 210842 197876 210898
rect 251274 220294 251330 220350
rect 251398 220294 251454 220350
rect 251522 220294 251578 220350
rect 251646 220294 251702 220350
rect 251274 220170 251330 220226
rect 251398 220170 251454 220226
rect 251522 220170 251578 220226
rect 251646 220170 251702 220226
rect 251274 220046 251330 220102
rect 251398 220046 251454 220102
rect 251522 220046 251578 220102
rect 251646 220046 251702 220102
rect 251274 219922 251330 219978
rect 251398 219922 251454 219978
rect 251522 219922 251578 219978
rect 251646 219922 251702 219978
rect 75238 202294 75294 202350
rect 75362 202294 75418 202350
rect 75238 202170 75294 202226
rect 75362 202170 75418 202226
rect 75238 202046 75294 202102
rect 75362 202046 75418 202102
rect 75238 201922 75294 201978
rect 75362 201922 75418 201978
rect 105958 202294 106014 202350
rect 106082 202294 106138 202350
rect 105958 202170 106014 202226
rect 106082 202170 106138 202226
rect 105958 202046 106014 202102
rect 106082 202046 106138 202102
rect 105958 201922 106014 201978
rect 106082 201922 106138 201978
rect 136678 202294 136734 202350
rect 136802 202294 136858 202350
rect 136678 202170 136734 202226
rect 136802 202170 136858 202226
rect 136678 202046 136734 202102
rect 136802 202046 136858 202102
rect 136678 201922 136734 201978
rect 136802 201922 136858 201978
rect 167398 202294 167454 202350
rect 167522 202294 167578 202350
rect 167398 202170 167454 202226
rect 167522 202170 167578 202226
rect 167398 202046 167454 202102
rect 167522 202046 167578 202102
rect 167398 201922 167454 201978
rect 167522 201922 167578 201978
rect 198118 202294 198174 202350
rect 198242 202294 198298 202350
rect 198118 202170 198174 202226
rect 198242 202170 198298 202226
rect 198118 202046 198174 202102
rect 198242 202046 198298 202102
rect 198118 201922 198174 201978
rect 198242 201922 198298 201978
rect 228838 202294 228894 202350
rect 228962 202294 229018 202350
rect 228838 202170 228894 202226
rect 228962 202170 229018 202226
rect 228838 202046 228894 202102
rect 228962 202046 229018 202102
rect 228838 201922 228894 201978
rect 228962 201922 229018 201978
rect 259558 202294 259614 202350
rect 259682 202294 259738 202350
rect 259558 202170 259614 202226
rect 259682 202170 259738 202226
rect 259558 202046 259614 202102
rect 259682 202046 259738 202102
rect 259558 201922 259614 201978
rect 259682 201922 259738 201978
rect 59878 190294 59934 190350
rect 60002 190294 60058 190350
rect 59878 190170 59934 190226
rect 60002 190170 60058 190226
rect 59878 190046 59934 190102
rect 60002 190046 60058 190102
rect 59878 189922 59934 189978
rect 60002 189922 60058 189978
rect 90598 190294 90654 190350
rect 90722 190294 90778 190350
rect 90598 190170 90654 190226
rect 90722 190170 90778 190226
rect 90598 190046 90654 190102
rect 90722 190046 90778 190102
rect 90598 189922 90654 189978
rect 90722 189922 90778 189978
rect 121318 190294 121374 190350
rect 121442 190294 121498 190350
rect 121318 190170 121374 190226
rect 121442 190170 121498 190226
rect 121318 190046 121374 190102
rect 121442 190046 121498 190102
rect 121318 189922 121374 189978
rect 121442 189922 121498 189978
rect 152038 190294 152094 190350
rect 152162 190294 152218 190350
rect 152038 190170 152094 190226
rect 152162 190170 152218 190226
rect 152038 190046 152094 190102
rect 152162 190046 152218 190102
rect 152038 189922 152094 189978
rect 152162 189922 152218 189978
rect 182758 190294 182814 190350
rect 182882 190294 182938 190350
rect 182758 190170 182814 190226
rect 182882 190170 182938 190226
rect 182758 190046 182814 190102
rect 182882 190046 182938 190102
rect 182758 189922 182814 189978
rect 182882 189922 182938 189978
rect 213478 190294 213534 190350
rect 213602 190294 213658 190350
rect 213478 190170 213534 190226
rect 213602 190170 213658 190226
rect 213478 190046 213534 190102
rect 213602 190046 213658 190102
rect 213478 189922 213534 189978
rect 213602 189922 213658 189978
rect 244198 190294 244254 190350
rect 244322 190294 244378 190350
rect 244198 190170 244254 190226
rect 244322 190170 244378 190226
rect 244198 190046 244254 190102
rect 244322 190046 244378 190102
rect 244198 189922 244254 189978
rect 244322 189922 244378 189978
rect 75238 184294 75294 184350
rect 75362 184294 75418 184350
rect 75238 184170 75294 184226
rect 75362 184170 75418 184226
rect 75238 184046 75294 184102
rect 75362 184046 75418 184102
rect 75238 183922 75294 183978
rect 75362 183922 75418 183978
rect 105958 184294 106014 184350
rect 106082 184294 106138 184350
rect 105958 184170 106014 184226
rect 106082 184170 106138 184226
rect 105958 184046 106014 184102
rect 106082 184046 106138 184102
rect 105958 183922 106014 183978
rect 106082 183922 106138 183978
rect 136678 184294 136734 184350
rect 136802 184294 136858 184350
rect 136678 184170 136734 184226
rect 136802 184170 136858 184226
rect 136678 184046 136734 184102
rect 136802 184046 136858 184102
rect 136678 183922 136734 183978
rect 136802 183922 136858 183978
rect 167398 184294 167454 184350
rect 167522 184294 167578 184350
rect 167398 184170 167454 184226
rect 167522 184170 167578 184226
rect 167398 184046 167454 184102
rect 167522 184046 167578 184102
rect 167398 183922 167454 183978
rect 167522 183922 167578 183978
rect 198118 184294 198174 184350
rect 198242 184294 198298 184350
rect 198118 184170 198174 184226
rect 198242 184170 198298 184226
rect 198118 184046 198174 184102
rect 198242 184046 198298 184102
rect 198118 183922 198174 183978
rect 198242 183922 198298 183978
rect 228838 184294 228894 184350
rect 228962 184294 229018 184350
rect 228838 184170 228894 184226
rect 228962 184170 229018 184226
rect 228838 184046 228894 184102
rect 228962 184046 229018 184102
rect 228838 183922 228894 183978
rect 228962 183922 229018 183978
rect 259558 184294 259614 184350
rect 259682 184294 259738 184350
rect 259558 184170 259614 184226
rect 259682 184170 259738 184226
rect 259558 184046 259614 184102
rect 259682 184046 259738 184102
rect 259558 183922 259614 183978
rect 259682 183922 259738 183978
rect 59878 172294 59934 172350
rect 60002 172294 60058 172350
rect 59878 172170 59934 172226
rect 60002 172170 60058 172226
rect 59878 172046 59934 172102
rect 60002 172046 60058 172102
rect 59878 171922 59934 171978
rect 60002 171922 60058 171978
rect 90598 172294 90654 172350
rect 90722 172294 90778 172350
rect 90598 172170 90654 172226
rect 90722 172170 90778 172226
rect 90598 172046 90654 172102
rect 90722 172046 90778 172102
rect 90598 171922 90654 171978
rect 90722 171922 90778 171978
rect 121318 172294 121374 172350
rect 121442 172294 121498 172350
rect 121318 172170 121374 172226
rect 121442 172170 121498 172226
rect 121318 172046 121374 172102
rect 121442 172046 121498 172102
rect 121318 171922 121374 171978
rect 121442 171922 121498 171978
rect 152038 172294 152094 172350
rect 152162 172294 152218 172350
rect 152038 172170 152094 172226
rect 152162 172170 152218 172226
rect 152038 172046 152094 172102
rect 152162 172046 152218 172102
rect 152038 171922 152094 171978
rect 152162 171922 152218 171978
rect 182758 172294 182814 172350
rect 182882 172294 182938 172350
rect 182758 172170 182814 172226
rect 182882 172170 182938 172226
rect 182758 172046 182814 172102
rect 182882 172046 182938 172102
rect 182758 171922 182814 171978
rect 182882 171922 182938 171978
rect 213478 172294 213534 172350
rect 213602 172294 213658 172350
rect 213478 172170 213534 172226
rect 213602 172170 213658 172226
rect 213478 172046 213534 172102
rect 213602 172046 213658 172102
rect 213478 171922 213534 171978
rect 213602 171922 213658 171978
rect 244198 172294 244254 172350
rect 244322 172294 244378 172350
rect 244198 172170 244254 172226
rect 244322 172170 244378 172226
rect 244198 172046 244254 172102
rect 244322 172046 244378 172102
rect 244198 171922 244254 171978
rect 244322 171922 244378 171978
rect 75238 166294 75294 166350
rect 75362 166294 75418 166350
rect 75238 166170 75294 166226
rect 75362 166170 75418 166226
rect 75238 166046 75294 166102
rect 75362 166046 75418 166102
rect 75238 165922 75294 165978
rect 75362 165922 75418 165978
rect 105958 166294 106014 166350
rect 106082 166294 106138 166350
rect 105958 166170 106014 166226
rect 106082 166170 106138 166226
rect 105958 166046 106014 166102
rect 106082 166046 106138 166102
rect 105958 165922 106014 165978
rect 106082 165922 106138 165978
rect 136678 166294 136734 166350
rect 136802 166294 136858 166350
rect 136678 166170 136734 166226
rect 136802 166170 136858 166226
rect 136678 166046 136734 166102
rect 136802 166046 136858 166102
rect 136678 165922 136734 165978
rect 136802 165922 136858 165978
rect 167398 166294 167454 166350
rect 167522 166294 167578 166350
rect 167398 166170 167454 166226
rect 167522 166170 167578 166226
rect 167398 166046 167454 166102
rect 167522 166046 167578 166102
rect 167398 165922 167454 165978
rect 167522 165922 167578 165978
rect 198118 166294 198174 166350
rect 198242 166294 198298 166350
rect 198118 166170 198174 166226
rect 198242 166170 198298 166226
rect 198118 166046 198174 166102
rect 198242 166046 198298 166102
rect 198118 165922 198174 165978
rect 198242 165922 198298 165978
rect 228838 166294 228894 166350
rect 228962 166294 229018 166350
rect 228838 166170 228894 166226
rect 228962 166170 229018 166226
rect 228838 166046 228894 166102
rect 228962 166046 229018 166102
rect 228838 165922 228894 165978
rect 228962 165922 229018 165978
rect 259558 166294 259614 166350
rect 259682 166294 259738 166350
rect 259558 166170 259614 166226
rect 259682 166170 259738 166226
rect 259558 166046 259614 166102
rect 259682 166046 259738 166102
rect 259558 165922 259614 165978
rect 259682 165922 259738 165978
rect 59878 154294 59934 154350
rect 60002 154294 60058 154350
rect 59878 154170 59934 154226
rect 60002 154170 60058 154226
rect 59878 154046 59934 154102
rect 60002 154046 60058 154102
rect 59878 153922 59934 153978
rect 60002 153922 60058 153978
rect 90598 154294 90654 154350
rect 90722 154294 90778 154350
rect 90598 154170 90654 154226
rect 90722 154170 90778 154226
rect 90598 154046 90654 154102
rect 90722 154046 90778 154102
rect 90598 153922 90654 153978
rect 90722 153922 90778 153978
rect 121318 154294 121374 154350
rect 121442 154294 121498 154350
rect 121318 154170 121374 154226
rect 121442 154170 121498 154226
rect 121318 154046 121374 154102
rect 121442 154046 121498 154102
rect 121318 153922 121374 153978
rect 121442 153922 121498 153978
rect 152038 154294 152094 154350
rect 152162 154294 152218 154350
rect 152038 154170 152094 154226
rect 152162 154170 152218 154226
rect 152038 154046 152094 154102
rect 152162 154046 152218 154102
rect 152038 153922 152094 153978
rect 152162 153922 152218 153978
rect 182758 154294 182814 154350
rect 182882 154294 182938 154350
rect 182758 154170 182814 154226
rect 182882 154170 182938 154226
rect 182758 154046 182814 154102
rect 182882 154046 182938 154102
rect 182758 153922 182814 153978
rect 182882 153922 182938 153978
rect 213478 154294 213534 154350
rect 213602 154294 213658 154350
rect 213478 154170 213534 154226
rect 213602 154170 213658 154226
rect 213478 154046 213534 154102
rect 213602 154046 213658 154102
rect 213478 153922 213534 153978
rect 213602 153922 213658 153978
rect 244198 154294 244254 154350
rect 244322 154294 244378 154350
rect 244198 154170 244254 154226
rect 244322 154170 244378 154226
rect 244198 154046 244254 154102
rect 244322 154046 244378 154102
rect 244198 153922 244254 153978
rect 244322 153922 244378 153978
rect 75238 148294 75294 148350
rect 75362 148294 75418 148350
rect 75238 148170 75294 148226
rect 75362 148170 75418 148226
rect 75238 148046 75294 148102
rect 75362 148046 75418 148102
rect 75238 147922 75294 147978
rect 75362 147922 75418 147978
rect 105958 148294 106014 148350
rect 106082 148294 106138 148350
rect 105958 148170 106014 148226
rect 106082 148170 106138 148226
rect 105958 148046 106014 148102
rect 106082 148046 106138 148102
rect 105958 147922 106014 147978
rect 106082 147922 106138 147978
rect 136678 148294 136734 148350
rect 136802 148294 136858 148350
rect 136678 148170 136734 148226
rect 136802 148170 136858 148226
rect 136678 148046 136734 148102
rect 136802 148046 136858 148102
rect 136678 147922 136734 147978
rect 136802 147922 136858 147978
rect 167398 148294 167454 148350
rect 167522 148294 167578 148350
rect 167398 148170 167454 148226
rect 167522 148170 167578 148226
rect 167398 148046 167454 148102
rect 167522 148046 167578 148102
rect 167398 147922 167454 147978
rect 167522 147922 167578 147978
rect 198118 148294 198174 148350
rect 198242 148294 198298 148350
rect 198118 148170 198174 148226
rect 198242 148170 198298 148226
rect 198118 148046 198174 148102
rect 198242 148046 198298 148102
rect 198118 147922 198174 147978
rect 198242 147922 198298 147978
rect 228838 148294 228894 148350
rect 228962 148294 229018 148350
rect 228838 148170 228894 148226
rect 228962 148170 229018 148226
rect 228838 148046 228894 148102
rect 228962 148046 229018 148102
rect 228838 147922 228894 147978
rect 228962 147922 229018 147978
rect 259558 148294 259614 148350
rect 259682 148294 259738 148350
rect 259558 148170 259614 148226
rect 259682 148170 259738 148226
rect 259558 148046 259614 148102
rect 259682 148046 259738 148102
rect 259558 147922 259614 147978
rect 259682 147922 259738 147978
rect 59878 136294 59934 136350
rect 60002 136294 60058 136350
rect 59878 136170 59934 136226
rect 60002 136170 60058 136226
rect 59878 136046 59934 136102
rect 60002 136046 60058 136102
rect 59878 135922 59934 135978
rect 60002 135922 60058 135978
rect 90598 136294 90654 136350
rect 90722 136294 90778 136350
rect 90598 136170 90654 136226
rect 90722 136170 90778 136226
rect 90598 136046 90654 136102
rect 90722 136046 90778 136102
rect 90598 135922 90654 135978
rect 90722 135922 90778 135978
rect 121318 136294 121374 136350
rect 121442 136294 121498 136350
rect 121318 136170 121374 136226
rect 121442 136170 121498 136226
rect 121318 136046 121374 136102
rect 121442 136046 121498 136102
rect 121318 135922 121374 135978
rect 121442 135922 121498 135978
rect 152038 136294 152094 136350
rect 152162 136294 152218 136350
rect 152038 136170 152094 136226
rect 152162 136170 152218 136226
rect 152038 136046 152094 136102
rect 152162 136046 152218 136102
rect 152038 135922 152094 135978
rect 152162 135922 152218 135978
rect 182758 136294 182814 136350
rect 182882 136294 182938 136350
rect 182758 136170 182814 136226
rect 182882 136170 182938 136226
rect 182758 136046 182814 136102
rect 182882 136046 182938 136102
rect 182758 135922 182814 135978
rect 182882 135922 182938 135978
rect 213478 136294 213534 136350
rect 213602 136294 213658 136350
rect 213478 136170 213534 136226
rect 213602 136170 213658 136226
rect 213478 136046 213534 136102
rect 213602 136046 213658 136102
rect 213478 135922 213534 135978
rect 213602 135922 213658 135978
rect 244198 136294 244254 136350
rect 244322 136294 244378 136350
rect 244198 136170 244254 136226
rect 244322 136170 244378 136226
rect 244198 136046 244254 136102
rect 244322 136046 244378 136102
rect 244198 135922 244254 135978
rect 244322 135922 244378 135978
rect 75238 130294 75294 130350
rect 75362 130294 75418 130350
rect 75238 130170 75294 130226
rect 75362 130170 75418 130226
rect 75238 130046 75294 130102
rect 75362 130046 75418 130102
rect 75238 129922 75294 129978
rect 75362 129922 75418 129978
rect 105958 130294 106014 130350
rect 106082 130294 106138 130350
rect 105958 130170 106014 130226
rect 106082 130170 106138 130226
rect 105958 130046 106014 130102
rect 106082 130046 106138 130102
rect 105958 129922 106014 129978
rect 106082 129922 106138 129978
rect 136678 130294 136734 130350
rect 136802 130294 136858 130350
rect 136678 130170 136734 130226
rect 136802 130170 136858 130226
rect 136678 130046 136734 130102
rect 136802 130046 136858 130102
rect 136678 129922 136734 129978
rect 136802 129922 136858 129978
rect 167398 130294 167454 130350
rect 167522 130294 167578 130350
rect 167398 130170 167454 130226
rect 167522 130170 167578 130226
rect 167398 130046 167454 130102
rect 167522 130046 167578 130102
rect 167398 129922 167454 129978
rect 167522 129922 167578 129978
rect 198118 130294 198174 130350
rect 198242 130294 198298 130350
rect 198118 130170 198174 130226
rect 198242 130170 198298 130226
rect 198118 130046 198174 130102
rect 198242 130046 198298 130102
rect 198118 129922 198174 129978
rect 198242 129922 198298 129978
rect 228838 130294 228894 130350
rect 228962 130294 229018 130350
rect 228838 130170 228894 130226
rect 228962 130170 229018 130226
rect 228838 130046 228894 130102
rect 228962 130046 229018 130102
rect 228838 129922 228894 129978
rect 228962 129922 229018 129978
rect 259558 130294 259614 130350
rect 259682 130294 259738 130350
rect 259558 130170 259614 130226
rect 259682 130170 259738 130226
rect 259558 130046 259614 130102
rect 259682 130046 259738 130102
rect 259558 129922 259614 129978
rect 259682 129922 259738 129978
rect 59878 118294 59934 118350
rect 60002 118294 60058 118350
rect 59878 118170 59934 118226
rect 60002 118170 60058 118226
rect 59878 118046 59934 118102
rect 60002 118046 60058 118102
rect 59878 117922 59934 117978
rect 60002 117922 60058 117978
rect 90598 118294 90654 118350
rect 90722 118294 90778 118350
rect 90598 118170 90654 118226
rect 90722 118170 90778 118226
rect 90598 118046 90654 118102
rect 90722 118046 90778 118102
rect 90598 117922 90654 117978
rect 90722 117922 90778 117978
rect 121318 118294 121374 118350
rect 121442 118294 121498 118350
rect 121318 118170 121374 118226
rect 121442 118170 121498 118226
rect 121318 118046 121374 118102
rect 121442 118046 121498 118102
rect 121318 117922 121374 117978
rect 121442 117922 121498 117978
rect 152038 118294 152094 118350
rect 152162 118294 152218 118350
rect 152038 118170 152094 118226
rect 152162 118170 152218 118226
rect 152038 118046 152094 118102
rect 152162 118046 152218 118102
rect 152038 117922 152094 117978
rect 152162 117922 152218 117978
rect 182758 118294 182814 118350
rect 182882 118294 182938 118350
rect 182758 118170 182814 118226
rect 182882 118170 182938 118226
rect 182758 118046 182814 118102
rect 182882 118046 182938 118102
rect 182758 117922 182814 117978
rect 182882 117922 182938 117978
rect 213478 118294 213534 118350
rect 213602 118294 213658 118350
rect 213478 118170 213534 118226
rect 213602 118170 213658 118226
rect 213478 118046 213534 118102
rect 213602 118046 213658 118102
rect 213478 117922 213534 117978
rect 213602 117922 213658 117978
rect 244198 118294 244254 118350
rect 244322 118294 244378 118350
rect 244198 118170 244254 118226
rect 244322 118170 244378 118226
rect 244198 118046 244254 118102
rect 244322 118046 244378 118102
rect 244198 117922 244254 117978
rect 244322 117922 244378 117978
rect 75238 112294 75294 112350
rect 75362 112294 75418 112350
rect 75238 112170 75294 112226
rect 75362 112170 75418 112226
rect 75238 112046 75294 112102
rect 75362 112046 75418 112102
rect 75238 111922 75294 111978
rect 75362 111922 75418 111978
rect 105958 112294 106014 112350
rect 106082 112294 106138 112350
rect 105958 112170 106014 112226
rect 106082 112170 106138 112226
rect 105958 112046 106014 112102
rect 106082 112046 106138 112102
rect 105958 111922 106014 111978
rect 106082 111922 106138 111978
rect 136678 112294 136734 112350
rect 136802 112294 136858 112350
rect 136678 112170 136734 112226
rect 136802 112170 136858 112226
rect 136678 112046 136734 112102
rect 136802 112046 136858 112102
rect 136678 111922 136734 111978
rect 136802 111922 136858 111978
rect 167398 112294 167454 112350
rect 167522 112294 167578 112350
rect 167398 112170 167454 112226
rect 167522 112170 167578 112226
rect 167398 112046 167454 112102
rect 167522 112046 167578 112102
rect 167398 111922 167454 111978
rect 167522 111922 167578 111978
rect 198118 112294 198174 112350
rect 198242 112294 198298 112350
rect 198118 112170 198174 112226
rect 198242 112170 198298 112226
rect 198118 112046 198174 112102
rect 198242 112046 198298 112102
rect 198118 111922 198174 111978
rect 198242 111922 198298 111978
rect 228838 112294 228894 112350
rect 228962 112294 229018 112350
rect 228838 112170 228894 112226
rect 228962 112170 229018 112226
rect 228838 112046 228894 112102
rect 228962 112046 229018 112102
rect 228838 111922 228894 111978
rect 228962 111922 229018 111978
rect 259558 112294 259614 112350
rect 259682 112294 259738 112350
rect 259558 112170 259614 112226
rect 259682 112170 259738 112226
rect 259558 112046 259614 112102
rect 259682 112046 259738 112102
rect 259558 111922 259614 111978
rect 259682 111922 259738 111978
rect 59878 100294 59934 100350
rect 60002 100294 60058 100350
rect 59878 100170 59934 100226
rect 60002 100170 60058 100226
rect 59878 100046 59934 100102
rect 60002 100046 60058 100102
rect 59878 99922 59934 99978
rect 60002 99922 60058 99978
rect 90598 100294 90654 100350
rect 90722 100294 90778 100350
rect 90598 100170 90654 100226
rect 90722 100170 90778 100226
rect 90598 100046 90654 100102
rect 90722 100046 90778 100102
rect 90598 99922 90654 99978
rect 90722 99922 90778 99978
rect 121318 100294 121374 100350
rect 121442 100294 121498 100350
rect 121318 100170 121374 100226
rect 121442 100170 121498 100226
rect 121318 100046 121374 100102
rect 121442 100046 121498 100102
rect 121318 99922 121374 99978
rect 121442 99922 121498 99978
rect 152038 100294 152094 100350
rect 152162 100294 152218 100350
rect 152038 100170 152094 100226
rect 152162 100170 152218 100226
rect 152038 100046 152094 100102
rect 152162 100046 152218 100102
rect 152038 99922 152094 99978
rect 152162 99922 152218 99978
rect 182758 100294 182814 100350
rect 182882 100294 182938 100350
rect 182758 100170 182814 100226
rect 182882 100170 182938 100226
rect 182758 100046 182814 100102
rect 182882 100046 182938 100102
rect 182758 99922 182814 99978
rect 182882 99922 182938 99978
rect 213478 100294 213534 100350
rect 213602 100294 213658 100350
rect 213478 100170 213534 100226
rect 213602 100170 213658 100226
rect 213478 100046 213534 100102
rect 213602 100046 213658 100102
rect 213478 99922 213534 99978
rect 213602 99922 213658 99978
rect 244198 100294 244254 100350
rect 244322 100294 244378 100350
rect 244198 100170 244254 100226
rect 244322 100170 244378 100226
rect 244198 100046 244254 100102
rect 244322 100046 244378 100102
rect 244198 99922 244254 99978
rect 244322 99922 244378 99978
rect 75238 94294 75294 94350
rect 75362 94294 75418 94350
rect 75238 94170 75294 94226
rect 75362 94170 75418 94226
rect 75238 94046 75294 94102
rect 75362 94046 75418 94102
rect 75238 93922 75294 93978
rect 75362 93922 75418 93978
rect 105958 94294 106014 94350
rect 106082 94294 106138 94350
rect 105958 94170 106014 94226
rect 106082 94170 106138 94226
rect 105958 94046 106014 94102
rect 106082 94046 106138 94102
rect 105958 93922 106014 93978
rect 106082 93922 106138 93978
rect 136678 94294 136734 94350
rect 136802 94294 136858 94350
rect 136678 94170 136734 94226
rect 136802 94170 136858 94226
rect 136678 94046 136734 94102
rect 136802 94046 136858 94102
rect 136678 93922 136734 93978
rect 136802 93922 136858 93978
rect 167398 94294 167454 94350
rect 167522 94294 167578 94350
rect 167398 94170 167454 94226
rect 167522 94170 167578 94226
rect 167398 94046 167454 94102
rect 167522 94046 167578 94102
rect 167398 93922 167454 93978
rect 167522 93922 167578 93978
rect 198118 94294 198174 94350
rect 198242 94294 198298 94350
rect 198118 94170 198174 94226
rect 198242 94170 198298 94226
rect 198118 94046 198174 94102
rect 198242 94046 198298 94102
rect 198118 93922 198174 93978
rect 198242 93922 198298 93978
rect 228838 94294 228894 94350
rect 228962 94294 229018 94350
rect 228838 94170 228894 94226
rect 228962 94170 229018 94226
rect 228838 94046 228894 94102
rect 228962 94046 229018 94102
rect 228838 93922 228894 93978
rect 228962 93922 229018 93978
rect 259558 94294 259614 94350
rect 259682 94294 259738 94350
rect 259558 94170 259614 94226
rect 259682 94170 259738 94226
rect 259558 94046 259614 94102
rect 259682 94046 259738 94102
rect 259558 93922 259614 93978
rect 259682 93922 259738 93978
rect 59878 82294 59934 82350
rect 60002 82294 60058 82350
rect 59878 82170 59934 82226
rect 60002 82170 60058 82226
rect 59878 82046 59934 82102
rect 60002 82046 60058 82102
rect 59878 81922 59934 81978
rect 60002 81922 60058 81978
rect 90598 82294 90654 82350
rect 90722 82294 90778 82350
rect 90598 82170 90654 82226
rect 90722 82170 90778 82226
rect 90598 82046 90654 82102
rect 90722 82046 90778 82102
rect 90598 81922 90654 81978
rect 90722 81922 90778 81978
rect 121318 82294 121374 82350
rect 121442 82294 121498 82350
rect 121318 82170 121374 82226
rect 121442 82170 121498 82226
rect 121318 82046 121374 82102
rect 121442 82046 121498 82102
rect 121318 81922 121374 81978
rect 121442 81922 121498 81978
rect 152038 82294 152094 82350
rect 152162 82294 152218 82350
rect 152038 82170 152094 82226
rect 152162 82170 152218 82226
rect 152038 82046 152094 82102
rect 152162 82046 152218 82102
rect 152038 81922 152094 81978
rect 152162 81922 152218 81978
rect 182758 82294 182814 82350
rect 182882 82294 182938 82350
rect 182758 82170 182814 82226
rect 182882 82170 182938 82226
rect 182758 82046 182814 82102
rect 182882 82046 182938 82102
rect 182758 81922 182814 81978
rect 182882 81922 182938 81978
rect 213478 82294 213534 82350
rect 213602 82294 213658 82350
rect 213478 82170 213534 82226
rect 213602 82170 213658 82226
rect 213478 82046 213534 82102
rect 213602 82046 213658 82102
rect 213478 81922 213534 81978
rect 213602 81922 213658 81978
rect 244198 82294 244254 82350
rect 244322 82294 244378 82350
rect 244198 82170 244254 82226
rect 244322 82170 244378 82226
rect 244198 82046 244254 82102
rect 244322 82046 244378 82102
rect 244198 81922 244254 81978
rect 244322 81922 244378 81978
rect 75238 76294 75294 76350
rect 75362 76294 75418 76350
rect 75238 76170 75294 76226
rect 75362 76170 75418 76226
rect 75238 76046 75294 76102
rect 75362 76046 75418 76102
rect 75238 75922 75294 75978
rect 75362 75922 75418 75978
rect 105958 76294 106014 76350
rect 106082 76294 106138 76350
rect 105958 76170 106014 76226
rect 106082 76170 106138 76226
rect 105958 76046 106014 76102
rect 106082 76046 106138 76102
rect 105958 75922 106014 75978
rect 106082 75922 106138 75978
rect 136678 76294 136734 76350
rect 136802 76294 136858 76350
rect 136678 76170 136734 76226
rect 136802 76170 136858 76226
rect 136678 76046 136734 76102
rect 136802 76046 136858 76102
rect 136678 75922 136734 75978
rect 136802 75922 136858 75978
rect 167398 76294 167454 76350
rect 167522 76294 167578 76350
rect 167398 76170 167454 76226
rect 167522 76170 167578 76226
rect 167398 76046 167454 76102
rect 167522 76046 167578 76102
rect 167398 75922 167454 75978
rect 167522 75922 167578 75978
rect 198118 76294 198174 76350
rect 198242 76294 198298 76350
rect 198118 76170 198174 76226
rect 198242 76170 198298 76226
rect 198118 76046 198174 76102
rect 198242 76046 198298 76102
rect 198118 75922 198174 75978
rect 198242 75922 198298 75978
rect 228838 76294 228894 76350
rect 228962 76294 229018 76350
rect 228838 76170 228894 76226
rect 228962 76170 229018 76226
rect 228838 76046 228894 76102
rect 228962 76046 229018 76102
rect 228838 75922 228894 75978
rect 228962 75922 229018 75978
rect 259558 76294 259614 76350
rect 259682 76294 259738 76350
rect 259558 76170 259614 76226
rect 259682 76170 259738 76226
rect 259558 76046 259614 76102
rect 259682 76046 259738 76102
rect 259558 75922 259614 75978
rect 259682 75922 259738 75978
rect 59878 64294 59934 64350
rect 60002 64294 60058 64350
rect 59878 64170 59934 64226
rect 60002 64170 60058 64226
rect 59878 64046 59934 64102
rect 60002 64046 60058 64102
rect 59878 63922 59934 63978
rect 60002 63922 60058 63978
rect 90598 64294 90654 64350
rect 90722 64294 90778 64350
rect 90598 64170 90654 64226
rect 90722 64170 90778 64226
rect 90598 64046 90654 64102
rect 90722 64046 90778 64102
rect 90598 63922 90654 63978
rect 90722 63922 90778 63978
rect 121318 64294 121374 64350
rect 121442 64294 121498 64350
rect 121318 64170 121374 64226
rect 121442 64170 121498 64226
rect 121318 64046 121374 64102
rect 121442 64046 121498 64102
rect 121318 63922 121374 63978
rect 121442 63922 121498 63978
rect 152038 64294 152094 64350
rect 152162 64294 152218 64350
rect 152038 64170 152094 64226
rect 152162 64170 152218 64226
rect 152038 64046 152094 64102
rect 152162 64046 152218 64102
rect 152038 63922 152094 63978
rect 152162 63922 152218 63978
rect 182758 64294 182814 64350
rect 182882 64294 182938 64350
rect 182758 64170 182814 64226
rect 182882 64170 182938 64226
rect 182758 64046 182814 64102
rect 182882 64046 182938 64102
rect 182758 63922 182814 63978
rect 182882 63922 182938 63978
rect 213478 64294 213534 64350
rect 213602 64294 213658 64350
rect 213478 64170 213534 64226
rect 213602 64170 213658 64226
rect 213478 64046 213534 64102
rect 213602 64046 213658 64102
rect 213478 63922 213534 63978
rect 213602 63922 213658 63978
rect 244198 64294 244254 64350
rect 244322 64294 244378 64350
rect 244198 64170 244254 64226
rect 244322 64170 244378 64226
rect 244198 64046 244254 64102
rect 244322 64046 244378 64102
rect 244198 63922 244254 63978
rect 244322 63922 244378 63978
rect 75238 58294 75294 58350
rect 75362 58294 75418 58350
rect 75238 58170 75294 58226
rect 75362 58170 75418 58226
rect 75238 58046 75294 58102
rect 75362 58046 75418 58102
rect 75238 57922 75294 57978
rect 75362 57922 75418 57978
rect 105958 58294 106014 58350
rect 106082 58294 106138 58350
rect 105958 58170 106014 58226
rect 106082 58170 106138 58226
rect 105958 58046 106014 58102
rect 106082 58046 106138 58102
rect 105958 57922 106014 57978
rect 106082 57922 106138 57978
rect 136678 58294 136734 58350
rect 136802 58294 136858 58350
rect 136678 58170 136734 58226
rect 136802 58170 136858 58226
rect 136678 58046 136734 58102
rect 136802 58046 136858 58102
rect 136678 57922 136734 57978
rect 136802 57922 136858 57978
rect 167398 58294 167454 58350
rect 167522 58294 167578 58350
rect 167398 58170 167454 58226
rect 167522 58170 167578 58226
rect 167398 58046 167454 58102
rect 167522 58046 167578 58102
rect 167398 57922 167454 57978
rect 167522 57922 167578 57978
rect 198118 58294 198174 58350
rect 198242 58294 198298 58350
rect 198118 58170 198174 58226
rect 198242 58170 198298 58226
rect 198118 58046 198174 58102
rect 198242 58046 198298 58102
rect 198118 57922 198174 57978
rect 198242 57922 198298 57978
rect 228838 58294 228894 58350
rect 228962 58294 229018 58350
rect 228838 58170 228894 58226
rect 228962 58170 229018 58226
rect 228838 58046 228894 58102
rect 228962 58046 229018 58102
rect 228838 57922 228894 57978
rect 228962 57922 229018 57978
rect 259558 58294 259614 58350
rect 259682 58294 259738 58350
rect 259558 58170 259614 58226
rect 259682 58170 259738 58226
rect 259558 58046 259614 58102
rect 259682 58046 259738 58102
rect 259558 57922 259614 57978
rect 259682 57922 259738 57978
rect 66954 40294 67010 40350
rect 67078 40294 67134 40350
rect 67202 40294 67258 40350
rect 67326 40294 67382 40350
rect 66954 40170 67010 40226
rect 67078 40170 67134 40226
rect 67202 40170 67258 40226
rect 67326 40170 67382 40226
rect 66954 40046 67010 40102
rect 67078 40046 67134 40102
rect 67202 40046 67258 40102
rect 67326 40046 67382 40102
rect 66954 39922 67010 39978
rect 67078 39922 67134 39978
rect 67202 39922 67258 39978
rect 67326 39922 67382 39978
rect 66954 22294 67010 22350
rect 67078 22294 67134 22350
rect 67202 22294 67258 22350
rect 67326 22294 67382 22350
rect 66954 22170 67010 22226
rect 67078 22170 67134 22226
rect 67202 22170 67258 22226
rect 67326 22170 67382 22226
rect 66954 22046 67010 22102
rect 67078 22046 67134 22102
rect 67202 22046 67258 22102
rect 67326 22046 67382 22102
rect 66954 21922 67010 21978
rect 67078 21922 67134 21978
rect 67202 21922 67258 21978
rect 67326 21922 67382 21978
rect 60844 4922 60900 4978
rect 55132 4742 55188 4798
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 39954 -1176 40010 -1120
rect 40078 -1176 40134 -1120
rect 40202 -1176 40258 -1120
rect 40326 -1176 40382 -1120
rect 39954 -1300 40010 -1244
rect 40078 -1300 40134 -1244
rect 40202 -1300 40258 -1244
rect 40326 -1300 40382 -1244
rect 39954 -1424 40010 -1368
rect 40078 -1424 40134 -1368
rect 40202 -1424 40258 -1368
rect 40326 -1424 40382 -1368
rect 39954 -1548 40010 -1492
rect 40078 -1548 40134 -1492
rect 40202 -1548 40258 -1492
rect 40326 -1548 40382 -1492
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 70674 46294 70730 46350
rect 70798 46294 70854 46350
rect 70922 46294 70978 46350
rect 71046 46294 71102 46350
rect 70674 46170 70730 46226
rect 70798 46170 70854 46226
rect 70922 46170 70978 46226
rect 71046 46170 71102 46226
rect 70674 46046 70730 46102
rect 70798 46046 70854 46102
rect 70922 46046 70978 46102
rect 71046 46046 71102 46102
rect 70674 45922 70730 45978
rect 70798 45922 70854 45978
rect 70922 45922 70978 45978
rect 71046 45922 71102 45978
rect 70674 28294 70730 28350
rect 70798 28294 70854 28350
rect 70922 28294 70978 28350
rect 71046 28294 71102 28350
rect 70674 28170 70730 28226
rect 70798 28170 70854 28226
rect 70922 28170 70978 28226
rect 71046 28170 71102 28226
rect 70674 28046 70730 28102
rect 70798 28046 70854 28102
rect 70922 28046 70978 28102
rect 71046 28046 71102 28102
rect 70674 27922 70730 27978
rect 70798 27922 70854 27978
rect 70922 27922 70978 27978
rect 71046 27922 71102 27978
rect 70674 10294 70730 10350
rect 70798 10294 70854 10350
rect 70922 10294 70978 10350
rect 71046 10294 71102 10350
rect 70674 10170 70730 10226
rect 70798 10170 70854 10226
rect 70922 10170 70978 10226
rect 71046 10170 71102 10226
rect 70674 10046 70730 10102
rect 70798 10046 70854 10102
rect 70922 10046 70978 10102
rect 71046 10046 71102 10102
rect 70674 9922 70730 9978
rect 70798 9922 70854 9978
rect 70922 9922 70978 9978
rect 71046 9922 71102 9978
rect 97674 40294 97730 40350
rect 97798 40294 97854 40350
rect 97922 40294 97978 40350
rect 98046 40294 98102 40350
rect 97674 40170 97730 40226
rect 97798 40170 97854 40226
rect 97922 40170 97978 40226
rect 98046 40170 98102 40226
rect 97674 40046 97730 40102
rect 97798 40046 97854 40102
rect 97922 40046 97978 40102
rect 98046 40046 98102 40102
rect 97674 39922 97730 39978
rect 97798 39922 97854 39978
rect 97922 39922 97978 39978
rect 98046 39922 98102 39978
rect 97674 22294 97730 22350
rect 97798 22294 97854 22350
rect 97922 22294 97978 22350
rect 98046 22294 98102 22350
rect 97674 22170 97730 22226
rect 97798 22170 97854 22226
rect 97922 22170 97978 22226
rect 98046 22170 98102 22226
rect 97674 22046 97730 22102
rect 97798 22046 97854 22102
rect 97922 22046 97978 22102
rect 98046 22046 98102 22102
rect 97674 21922 97730 21978
rect 97798 21922 97854 21978
rect 97922 21922 97978 21978
rect 98046 21922 98102 21978
rect 91532 4922 91588 4978
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 70674 -1176 70730 -1120
rect 70798 -1176 70854 -1120
rect 70922 -1176 70978 -1120
rect 71046 -1176 71102 -1120
rect 70674 -1300 70730 -1244
rect 70798 -1300 70854 -1244
rect 70922 -1300 70978 -1244
rect 71046 -1300 71102 -1244
rect 70674 -1424 70730 -1368
rect 70798 -1424 70854 -1368
rect 70922 -1424 70978 -1368
rect 71046 -1424 71102 -1368
rect 70674 -1548 70730 -1492
rect 70798 -1548 70854 -1492
rect 70922 -1548 70978 -1492
rect 71046 -1548 71102 -1492
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 101394 46294 101450 46350
rect 101518 46294 101574 46350
rect 101642 46294 101698 46350
rect 101766 46294 101822 46350
rect 101394 46170 101450 46226
rect 101518 46170 101574 46226
rect 101642 46170 101698 46226
rect 101766 46170 101822 46226
rect 101394 46046 101450 46102
rect 101518 46046 101574 46102
rect 101642 46046 101698 46102
rect 101766 46046 101822 46102
rect 101394 45922 101450 45978
rect 101518 45922 101574 45978
rect 101642 45922 101698 45978
rect 101766 45922 101822 45978
rect 101394 28294 101450 28350
rect 101518 28294 101574 28350
rect 101642 28294 101698 28350
rect 101766 28294 101822 28350
rect 101394 28170 101450 28226
rect 101518 28170 101574 28226
rect 101642 28170 101698 28226
rect 101766 28170 101822 28226
rect 101394 28046 101450 28102
rect 101518 28046 101574 28102
rect 101642 28046 101698 28102
rect 101766 28046 101822 28102
rect 101394 27922 101450 27978
rect 101518 27922 101574 27978
rect 101642 27922 101698 27978
rect 101766 27922 101822 27978
rect 101394 10294 101450 10350
rect 101518 10294 101574 10350
rect 101642 10294 101698 10350
rect 101766 10294 101822 10350
rect 101394 10170 101450 10226
rect 101518 10170 101574 10226
rect 101642 10170 101698 10226
rect 101766 10170 101822 10226
rect 101394 10046 101450 10102
rect 101518 10046 101574 10102
rect 101642 10046 101698 10102
rect 101766 10046 101822 10102
rect 101394 9922 101450 9978
rect 101518 9922 101574 9978
rect 101642 9922 101698 9978
rect 101766 9922 101822 9978
rect 101394 -1176 101450 -1120
rect 101518 -1176 101574 -1120
rect 101642 -1176 101698 -1120
rect 101766 -1176 101822 -1120
rect 101394 -1300 101450 -1244
rect 101518 -1300 101574 -1244
rect 101642 -1300 101698 -1244
rect 101766 -1300 101822 -1244
rect 101394 -1424 101450 -1368
rect 101518 -1424 101574 -1368
rect 101642 -1424 101698 -1368
rect 101766 -1424 101822 -1368
rect 101394 -1548 101450 -1492
rect 101518 -1548 101574 -1492
rect 101642 -1548 101698 -1492
rect 101766 -1548 101822 -1492
rect 128394 40294 128450 40350
rect 128518 40294 128574 40350
rect 128642 40294 128698 40350
rect 128766 40294 128822 40350
rect 128394 40170 128450 40226
rect 128518 40170 128574 40226
rect 128642 40170 128698 40226
rect 128766 40170 128822 40226
rect 128394 40046 128450 40102
rect 128518 40046 128574 40102
rect 128642 40046 128698 40102
rect 128766 40046 128822 40102
rect 128394 39922 128450 39978
rect 128518 39922 128574 39978
rect 128642 39922 128698 39978
rect 128766 39922 128822 39978
rect 128394 22294 128450 22350
rect 128518 22294 128574 22350
rect 128642 22294 128698 22350
rect 128766 22294 128822 22350
rect 128394 22170 128450 22226
rect 128518 22170 128574 22226
rect 128642 22170 128698 22226
rect 128766 22170 128822 22226
rect 128394 22046 128450 22102
rect 128518 22046 128574 22102
rect 128642 22046 128698 22102
rect 128766 22046 128822 22102
rect 128394 21922 128450 21978
rect 128518 21922 128574 21978
rect 128642 21922 128698 21978
rect 128766 21922 128822 21978
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 132114 46294 132170 46350
rect 132238 46294 132294 46350
rect 132362 46294 132418 46350
rect 132486 46294 132542 46350
rect 132114 46170 132170 46226
rect 132238 46170 132294 46226
rect 132362 46170 132418 46226
rect 132486 46170 132542 46226
rect 132114 46046 132170 46102
rect 132238 46046 132294 46102
rect 132362 46046 132418 46102
rect 132486 46046 132542 46102
rect 132114 45922 132170 45978
rect 132238 45922 132294 45978
rect 132362 45922 132418 45978
rect 132486 45922 132542 45978
rect 132114 28294 132170 28350
rect 132238 28294 132294 28350
rect 132362 28294 132418 28350
rect 132486 28294 132542 28350
rect 132114 28170 132170 28226
rect 132238 28170 132294 28226
rect 132362 28170 132418 28226
rect 132486 28170 132542 28226
rect 132114 28046 132170 28102
rect 132238 28046 132294 28102
rect 132362 28046 132418 28102
rect 132486 28046 132542 28102
rect 132114 27922 132170 27978
rect 132238 27922 132294 27978
rect 132362 27922 132418 27978
rect 132486 27922 132542 27978
rect 132114 10294 132170 10350
rect 132238 10294 132294 10350
rect 132362 10294 132418 10350
rect 132486 10294 132542 10350
rect 132114 10170 132170 10226
rect 132238 10170 132294 10226
rect 132362 10170 132418 10226
rect 132486 10170 132542 10226
rect 132114 10046 132170 10102
rect 132238 10046 132294 10102
rect 132362 10046 132418 10102
rect 132486 10046 132542 10102
rect 132114 9922 132170 9978
rect 132238 9922 132294 9978
rect 132362 9922 132418 9978
rect 132486 9922 132542 9978
rect 159114 40294 159170 40350
rect 159238 40294 159294 40350
rect 159362 40294 159418 40350
rect 159486 40294 159542 40350
rect 159114 40170 159170 40226
rect 159238 40170 159294 40226
rect 159362 40170 159418 40226
rect 159486 40170 159542 40226
rect 159114 40046 159170 40102
rect 159238 40046 159294 40102
rect 159362 40046 159418 40102
rect 159486 40046 159542 40102
rect 159114 39922 159170 39978
rect 159238 39922 159294 39978
rect 159362 39922 159418 39978
rect 159486 39922 159542 39978
rect 159114 22294 159170 22350
rect 159238 22294 159294 22350
rect 159362 22294 159418 22350
rect 159486 22294 159542 22350
rect 159114 22170 159170 22226
rect 159238 22170 159294 22226
rect 159362 22170 159418 22226
rect 159486 22170 159542 22226
rect 159114 22046 159170 22102
rect 159238 22046 159294 22102
rect 159362 22046 159418 22102
rect 159486 22046 159542 22102
rect 159114 21922 159170 21978
rect 159238 21922 159294 21978
rect 159362 21922 159418 21978
rect 159486 21922 159542 21978
rect 142940 4742 142996 4798
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 132114 -1176 132170 -1120
rect 132238 -1176 132294 -1120
rect 132362 -1176 132418 -1120
rect 132486 -1176 132542 -1120
rect 132114 -1300 132170 -1244
rect 132238 -1300 132294 -1244
rect 132362 -1300 132418 -1244
rect 132486 -1300 132542 -1244
rect 132114 -1424 132170 -1368
rect 132238 -1424 132294 -1368
rect 132362 -1424 132418 -1368
rect 132486 -1424 132542 -1368
rect 132114 -1548 132170 -1492
rect 132238 -1548 132294 -1492
rect 132362 -1548 132418 -1492
rect 132486 -1548 132542 -1492
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 162834 46294 162890 46350
rect 162958 46294 163014 46350
rect 163082 46294 163138 46350
rect 163206 46294 163262 46350
rect 162834 46170 162890 46226
rect 162958 46170 163014 46226
rect 163082 46170 163138 46226
rect 163206 46170 163262 46226
rect 162834 46046 162890 46102
rect 162958 46046 163014 46102
rect 163082 46046 163138 46102
rect 163206 46046 163262 46102
rect 162834 45922 162890 45978
rect 162958 45922 163014 45978
rect 163082 45922 163138 45978
rect 163206 45922 163262 45978
rect 162834 28294 162890 28350
rect 162958 28294 163014 28350
rect 163082 28294 163138 28350
rect 163206 28294 163262 28350
rect 162834 28170 162890 28226
rect 162958 28170 163014 28226
rect 163082 28170 163138 28226
rect 163206 28170 163262 28226
rect 162834 28046 162890 28102
rect 162958 28046 163014 28102
rect 163082 28046 163138 28102
rect 163206 28046 163262 28102
rect 162834 27922 162890 27978
rect 162958 27922 163014 27978
rect 163082 27922 163138 27978
rect 163206 27922 163262 27978
rect 162834 10294 162890 10350
rect 162958 10294 163014 10350
rect 163082 10294 163138 10350
rect 163206 10294 163262 10350
rect 162834 10170 162890 10226
rect 162958 10170 163014 10226
rect 163082 10170 163138 10226
rect 163206 10170 163262 10226
rect 162834 10046 162890 10102
rect 162958 10046 163014 10102
rect 163082 10046 163138 10102
rect 163206 10046 163262 10102
rect 162834 9922 162890 9978
rect 162958 9922 163014 9978
rect 163082 9922 163138 9978
rect 163206 9922 163262 9978
rect 172956 47762 173012 47818
rect 189834 40294 189890 40350
rect 189958 40294 190014 40350
rect 190082 40294 190138 40350
rect 190206 40294 190262 40350
rect 189834 40170 189890 40226
rect 189958 40170 190014 40226
rect 190082 40170 190138 40226
rect 190206 40170 190262 40226
rect 189834 40046 189890 40102
rect 189958 40046 190014 40102
rect 190082 40046 190138 40102
rect 190206 40046 190262 40102
rect 189834 39922 189890 39978
rect 189958 39922 190014 39978
rect 190082 39922 190138 39978
rect 190206 39922 190262 39978
rect 189834 22294 189890 22350
rect 189958 22294 190014 22350
rect 190082 22294 190138 22350
rect 190206 22294 190262 22350
rect 189834 22170 189890 22226
rect 189958 22170 190014 22226
rect 190082 22170 190138 22226
rect 190206 22170 190262 22226
rect 189834 22046 189890 22102
rect 189958 22046 190014 22102
rect 190082 22046 190138 22102
rect 190206 22046 190262 22102
rect 189834 21922 189890 21978
rect 189958 21922 190014 21978
rect 190082 21922 190138 21978
rect 190206 21922 190262 21978
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 162834 -1176 162890 -1120
rect 162958 -1176 163014 -1120
rect 163082 -1176 163138 -1120
rect 163206 -1176 163262 -1120
rect 162834 -1300 162890 -1244
rect 162958 -1300 163014 -1244
rect 163082 -1300 163138 -1244
rect 163206 -1300 163262 -1244
rect 162834 -1424 162890 -1368
rect 162958 -1424 163014 -1368
rect 163082 -1424 163138 -1368
rect 163206 -1424 163262 -1368
rect 162834 -1548 162890 -1492
rect 162958 -1548 163014 -1492
rect 163082 -1548 163138 -1492
rect 163206 -1548 163262 -1492
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 193554 46294 193610 46350
rect 193678 46294 193734 46350
rect 193802 46294 193858 46350
rect 193926 46294 193982 46350
rect 193554 46170 193610 46226
rect 193678 46170 193734 46226
rect 193802 46170 193858 46226
rect 193926 46170 193982 46226
rect 193554 46046 193610 46102
rect 193678 46046 193734 46102
rect 193802 46046 193858 46102
rect 193926 46046 193982 46102
rect 193554 45922 193610 45978
rect 193678 45922 193734 45978
rect 193802 45922 193858 45978
rect 193926 45922 193982 45978
rect 193554 28294 193610 28350
rect 193678 28294 193734 28350
rect 193802 28294 193858 28350
rect 193926 28294 193982 28350
rect 193554 28170 193610 28226
rect 193678 28170 193734 28226
rect 193802 28170 193858 28226
rect 193926 28170 193982 28226
rect 193554 28046 193610 28102
rect 193678 28046 193734 28102
rect 193802 28046 193858 28102
rect 193926 28046 193982 28102
rect 193554 27922 193610 27978
rect 193678 27922 193734 27978
rect 193802 27922 193858 27978
rect 193926 27922 193982 27978
rect 193554 10294 193610 10350
rect 193678 10294 193734 10350
rect 193802 10294 193858 10350
rect 193926 10294 193982 10350
rect 193554 10170 193610 10226
rect 193678 10170 193734 10226
rect 193802 10170 193858 10226
rect 193926 10170 193982 10226
rect 193554 10046 193610 10102
rect 193678 10046 193734 10102
rect 193802 10046 193858 10102
rect 193926 10046 193982 10102
rect 193554 9922 193610 9978
rect 193678 9922 193734 9978
rect 193802 9922 193858 9978
rect 193926 9922 193982 9978
rect 209132 47942 209188 47998
rect 220554 40294 220610 40350
rect 220678 40294 220734 40350
rect 220802 40294 220858 40350
rect 220926 40294 220982 40350
rect 220554 40170 220610 40226
rect 220678 40170 220734 40226
rect 220802 40170 220858 40226
rect 220926 40170 220982 40226
rect 220554 40046 220610 40102
rect 220678 40046 220734 40102
rect 220802 40046 220858 40102
rect 220926 40046 220982 40102
rect 220554 39922 220610 39978
rect 220678 39922 220734 39978
rect 220802 39922 220858 39978
rect 220926 39922 220982 39978
rect 220554 22294 220610 22350
rect 220678 22294 220734 22350
rect 220802 22294 220858 22350
rect 220926 22294 220982 22350
rect 220554 22170 220610 22226
rect 220678 22170 220734 22226
rect 220802 22170 220858 22226
rect 220926 22170 220982 22226
rect 220554 22046 220610 22102
rect 220678 22046 220734 22102
rect 220802 22046 220858 22102
rect 220926 22046 220982 22102
rect 220554 21922 220610 21978
rect 220678 21922 220734 21978
rect 220802 21922 220858 21978
rect 220926 21922 220982 21978
rect 193554 -1176 193610 -1120
rect 193678 -1176 193734 -1120
rect 193802 -1176 193858 -1120
rect 193926 -1176 193982 -1120
rect 193554 -1300 193610 -1244
rect 193678 -1300 193734 -1244
rect 193802 -1300 193858 -1244
rect 193926 -1300 193982 -1244
rect 193554 -1424 193610 -1368
rect 193678 -1424 193734 -1368
rect 193802 -1424 193858 -1368
rect 193926 -1424 193982 -1368
rect 193554 -1548 193610 -1492
rect 193678 -1548 193734 -1492
rect 193802 -1548 193858 -1492
rect 193926 -1548 193982 -1492
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 224274 46294 224330 46350
rect 224398 46294 224454 46350
rect 224522 46294 224578 46350
rect 224646 46294 224702 46350
rect 224274 46170 224330 46226
rect 224398 46170 224454 46226
rect 224522 46170 224578 46226
rect 224646 46170 224702 46226
rect 224274 46046 224330 46102
rect 224398 46046 224454 46102
rect 224522 46046 224578 46102
rect 224646 46046 224702 46102
rect 224274 45922 224330 45978
rect 224398 45922 224454 45978
rect 224522 45922 224578 45978
rect 224646 45922 224702 45978
rect 224274 28294 224330 28350
rect 224398 28294 224454 28350
rect 224522 28294 224578 28350
rect 224646 28294 224702 28350
rect 224274 28170 224330 28226
rect 224398 28170 224454 28226
rect 224522 28170 224578 28226
rect 224646 28170 224702 28226
rect 224274 28046 224330 28102
rect 224398 28046 224454 28102
rect 224522 28046 224578 28102
rect 224646 28046 224702 28102
rect 224274 27922 224330 27978
rect 224398 27922 224454 27978
rect 224522 27922 224578 27978
rect 224646 27922 224702 27978
rect 224274 10294 224330 10350
rect 224398 10294 224454 10350
rect 224522 10294 224578 10350
rect 224646 10294 224702 10350
rect 224274 10170 224330 10226
rect 224398 10170 224454 10226
rect 224522 10170 224578 10226
rect 224646 10170 224702 10226
rect 224274 10046 224330 10102
rect 224398 10046 224454 10102
rect 224522 10046 224578 10102
rect 224646 10046 224702 10102
rect 224274 9922 224330 9978
rect 224398 9922 224454 9978
rect 224522 9922 224578 9978
rect 224646 9922 224702 9978
rect 224274 -1176 224330 -1120
rect 224398 -1176 224454 -1120
rect 224522 -1176 224578 -1120
rect 224646 -1176 224702 -1120
rect 224274 -1300 224330 -1244
rect 224398 -1300 224454 -1244
rect 224522 -1300 224578 -1244
rect 224646 -1300 224702 -1244
rect 224274 -1424 224330 -1368
rect 224398 -1424 224454 -1368
rect 224522 -1424 224578 -1368
rect 224646 -1424 224702 -1368
rect 224274 -1548 224330 -1492
rect 224398 -1548 224454 -1492
rect 224522 -1548 224578 -1492
rect 224646 -1548 224702 -1492
rect 251274 40294 251330 40350
rect 251398 40294 251454 40350
rect 251522 40294 251578 40350
rect 251646 40294 251702 40350
rect 251274 40170 251330 40226
rect 251398 40170 251454 40226
rect 251522 40170 251578 40226
rect 251646 40170 251702 40226
rect 251274 40046 251330 40102
rect 251398 40046 251454 40102
rect 251522 40046 251578 40102
rect 251646 40046 251702 40102
rect 251274 39922 251330 39978
rect 251398 39922 251454 39978
rect 251522 39922 251578 39978
rect 251646 39922 251702 39978
rect 251274 22294 251330 22350
rect 251398 22294 251454 22350
rect 251522 22294 251578 22350
rect 251646 22294 251702 22350
rect 251274 22170 251330 22226
rect 251398 22170 251454 22226
rect 251522 22170 251578 22226
rect 251646 22170 251702 22226
rect 251274 22046 251330 22102
rect 251398 22046 251454 22102
rect 251522 22046 251578 22102
rect 251646 22046 251702 22102
rect 251274 21922 251330 21978
rect 251398 21922 251454 21978
rect 251522 21922 251578 21978
rect 251646 21922 251702 21978
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 254994 46294 255050 46350
rect 255118 46294 255174 46350
rect 255242 46294 255298 46350
rect 255366 46294 255422 46350
rect 254994 46170 255050 46226
rect 255118 46170 255174 46226
rect 255242 46170 255298 46226
rect 255366 46170 255422 46226
rect 254994 46046 255050 46102
rect 255118 46046 255174 46102
rect 255242 46046 255298 46102
rect 255366 46046 255422 46102
rect 254994 45922 255050 45978
rect 255118 45922 255174 45978
rect 255242 45922 255298 45978
rect 255366 45922 255422 45978
rect 254994 28294 255050 28350
rect 255118 28294 255174 28350
rect 255242 28294 255298 28350
rect 255366 28294 255422 28350
rect 254994 28170 255050 28226
rect 255118 28170 255174 28226
rect 255242 28170 255298 28226
rect 255366 28170 255422 28226
rect 254994 28046 255050 28102
rect 255118 28046 255174 28102
rect 255242 28046 255298 28102
rect 255366 28046 255422 28102
rect 254994 27922 255050 27978
rect 255118 27922 255174 27978
rect 255242 27922 255298 27978
rect 255366 27922 255422 27978
rect 268604 136862 268660 136918
rect 268716 133442 268772 133498
rect 269724 231362 269780 231418
rect 269836 227762 269892 227818
rect 270508 234422 270564 234478
rect 270844 231182 270900 231238
rect 272524 153636 272580 153658
rect 272524 153602 272580 153636
rect 275548 237122 275604 237178
rect 254994 10294 255050 10350
rect 255118 10294 255174 10350
rect 255242 10294 255298 10350
rect 255366 10294 255422 10350
rect 254994 10170 255050 10226
rect 255118 10170 255174 10226
rect 255242 10170 255298 10226
rect 255366 10170 255422 10226
rect 254994 10046 255050 10102
rect 255118 10046 255174 10102
rect 255242 10046 255298 10102
rect 255366 10046 255422 10102
rect 254994 9922 255050 9978
rect 255118 9922 255174 9978
rect 255242 9922 255298 9978
rect 255366 9922 255422 9978
rect 275660 236942 275716 236998
rect 281372 240542 281428 240598
rect 279692 239282 279748 239338
rect 278012 150362 278068 150418
rect 284956 240722 285012 240778
rect 281994 238294 282050 238350
rect 282118 238294 282174 238350
rect 282242 238294 282298 238350
rect 282366 238294 282422 238350
rect 281994 238170 282050 238226
rect 282118 238170 282174 238226
rect 282242 238170 282298 238226
rect 282366 238170 282422 238226
rect 281994 238046 282050 238102
rect 282118 238046 282174 238102
rect 282242 238046 282298 238102
rect 282366 238046 282422 238102
rect 281994 237922 282050 237978
rect 282118 237922 282174 237978
rect 282242 237922 282298 237978
rect 282366 237922 282422 237978
rect 284732 240362 284788 240418
rect 281994 220294 282050 220350
rect 282118 220294 282174 220350
rect 282242 220294 282298 220350
rect 282366 220294 282422 220350
rect 281994 220170 282050 220226
rect 282118 220170 282174 220226
rect 282242 220170 282298 220226
rect 282366 220170 282422 220226
rect 281994 220046 282050 220102
rect 282118 220046 282174 220102
rect 282242 220046 282298 220102
rect 282366 220046 282422 220102
rect 281994 219922 282050 219978
rect 282118 219922 282174 219978
rect 282242 219922 282298 219978
rect 282366 219922 282422 219978
rect 281994 202294 282050 202350
rect 282118 202294 282174 202350
rect 282242 202294 282298 202350
rect 282366 202294 282422 202350
rect 281994 202170 282050 202226
rect 282118 202170 282174 202226
rect 282242 202170 282298 202226
rect 282366 202170 282422 202226
rect 281994 202046 282050 202102
rect 282118 202046 282174 202102
rect 282242 202046 282298 202102
rect 282366 202046 282422 202102
rect 281994 201922 282050 201978
rect 282118 201922 282174 201978
rect 282242 201922 282298 201978
rect 282366 201922 282422 201978
rect 281994 184294 282050 184350
rect 282118 184294 282174 184350
rect 282242 184294 282298 184350
rect 282366 184294 282422 184350
rect 281994 184170 282050 184226
rect 282118 184170 282174 184226
rect 282242 184170 282298 184226
rect 282366 184170 282422 184226
rect 281994 184046 282050 184102
rect 282118 184046 282174 184102
rect 282242 184046 282298 184102
rect 282366 184046 282422 184102
rect 281994 183922 282050 183978
rect 282118 183922 282174 183978
rect 282242 183922 282298 183978
rect 282366 183922 282422 183978
rect 281994 166294 282050 166350
rect 282118 166294 282174 166350
rect 282242 166294 282298 166350
rect 282366 166294 282422 166350
rect 281994 166170 282050 166226
rect 282118 166170 282174 166226
rect 282242 166170 282298 166226
rect 282366 166170 282422 166226
rect 281994 166046 282050 166102
rect 282118 166046 282174 166102
rect 282242 166046 282298 166102
rect 282366 166046 282422 166102
rect 281994 165922 282050 165978
rect 282118 165922 282174 165978
rect 282242 165922 282298 165978
rect 282366 165922 282422 165978
rect 281994 148294 282050 148350
rect 282118 148294 282174 148350
rect 282242 148294 282298 148350
rect 282366 148294 282422 148350
rect 281994 148170 282050 148226
rect 282118 148170 282174 148226
rect 282242 148170 282298 148226
rect 282366 148170 282422 148226
rect 281994 148046 282050 148102
rect 282118 148046 282174 148102
rect 282242 148046 282298 148102
rect 282366 148046 282422 148102
rect 281994 147922 282050 147978
rect 282118 147922 282174 147978
rect 282242 147922 282298 147978
rect 282366 147922 282422 147978
rect 281994 130294 282050 130350
rect 282118 130294 282174 130350
rect 282242 130294 282298 130350
rect 282366 130294 282422 130350
rect 281994 130170 282050 130226
rect 282118 130170 282174 130226
rect 282242 130170 282298 130226
rect 282366 130170 282422 130226
rect 281994 130046 282050 130102
rect 282118 130046 282174 130102
rect 282242 130046 282298 130102
rect 282366 130046 282422 130102
rect 281994 129922 282050 129978
rect 282118 129922 282174 129978
rect 282242 129922 282298 129978
rect 282366 129922 282422 129978
rect 281994 112294 282050 112350
rect 282118 112294 282174 112350
rect 282242 112294 282298 112350
rect 282366 112294 282422 112350
rect 281994 112170 282050 112226
rect 282118 112170 282174 112226
rect 282242 112170 282298 112226
rect 282366 112170 282422 112226
rect 281994 112046 282050 112102
rect 282118 112046 282174 112102
rect 282242 112046 282298 112102
rect 282366 112046 282422 112102
rect 281994 111922 282050 111978
rect 282118 111922 282174 111978
rect 282242 111922 282298 111978
rect 282366 111922 282422 111978
rect 281994 94294 282050 94350
rect 282118 94294 282174 94350
rect 282242 94294 282298 94350
rect 282366 94294 282422 94350
rect 281994 94170 282050 94226
rect 282118 94170 282174 94226
rect 282242 94170 282298 94226
rect 282366 94170 282422 94226
rect 281994 94046 282050 94102
rect 282118 94046 282174 94102
rect 282242 94046 282298 94102
rect 282366 94046 282422 94102
rect 281994 93922 282050 93978
rect 282118 93922 282174 93978
rect 282242 93922 282298 93978
rect 282366 93922 282422 93978
rect 281994 76294 282050 76350
rect 282118 76294 282174 76350
rect 282242 76294 282298 76350
rect 282366 76294 282422 76350
rect 281994 76170 282050 76226
rect 282118 76170 282174 76226
rect 282242 76170 282298 76226
rect 282366 76170 282422 76226
rect 281994 76046 282050 76102
rect 282118 76046 282174 76102
rect 282242 76046 282298 76102
rect 282366 76046 282422 76102
rect 281994 75922 282050 75978
rect 282118 75922 282174 75978
rect 282242 75922 282298 75978
rect 282366 75922 282422 75978
rect 281994 58294 282050 58350
rect 282118 58294 282174 58350
rect 282242 58294 282298 58350
rect 282366 58294 282422 58350
rect 281994 58170 282050 58226
rect 282118 58170 282174 58226
rect 282242 58170 282298 58226
rect 282366 58170 282422 58226
rect 281994 58046 282050 58102
rect 282118 58046 282174 58102
rect 282242 58046 282298 58102
rect 282366 58046 282422 58102
rect 281994 57922 282050 57978
rect 282118 57922 282174 57978
rect 282242 57922 282298 57978
rect 282366 57922 282422 57978
rect 281994 40294 282050 40350
rect 282118 40294 282174 40350
rect 282242 40294 282298 40350
rect 282366 40294 282422 40350
rect 281994 40170 282050 40226
rect 282118 40170 282174 40226
rect 282242 40170 282298 40226
rect 282366 40170 282422 40226
rect 281994 40046 282050 40102
rect 282118 40046 282174 40102
rect 282242 40046 282298 40102
rect 282366 40046 282422 40102
rect 281994 39922 282050 39978
rect 282118 39922 282174 39978
rect 282242 39922 282298 39978
rect 282366 39922 282422 39978
rect 281994 22294 282050 22350
rect 282118 22294 282174 22350
rect 282242 22294 282298 22350
rect 282366 22294 282422 22350
rect 281994 22170 282050 22226
rect 282118 22170 282174 22226
rect 282242 22170 282298 22226
rect 282366 22170 282422 22226
rect 281994 22046 282050 22102
rect 282118 22046 282174 22102
rect 282242 22046 282298 22102
rect 282366 22046 282422 22102
rect 281994 21922 282050 21978
rect 282118 21922 282174 21978
rect 282242 21922 282298 21978
rect 282366 21922 282422 21978
rect 254994 -1176 255050 -1120
rect 255118 -1176 255174 -1120
rect 255242 -1176 255298 -1120
rect 255366 -1176 255422 -1120
rect 254994 -1300 255050 -1244
rect 255118 -1300 255174 -1244
rect 255242 -1300 255298 -1244
rect 255366 -1300 255422 -1244
rect 254994 -1424 255050 -1368
rect 255118 -1424 255174 -1368
rect 255242 -1424 255298 -1368
rect 255366 -1424 255422 -1368
rect 254994 -1548 255050 -1492
rect 255118 -1548 255174 -1492
rect 255242 -1548 255298 -1492
rect 255366 -1548 255422 -1492
rect 283052 234422 283108 234478
rect 284732 4742 284788 4798
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 285180 236042 285236 236098
rect 312714 238294 312770 238350
rect 312838 238294 312894 238350
rect 312962 238294 313018 238350
rect 313086 238294 313142 238350
rect 312714 238170 312770 238226
rect 312838 238170 312894 238226
rect 312962 238170 313018 238226
rect 313086 238170 313142 238226
rect 312714 238046 312770 238102
rect 312838 238046 312894 238102
rect 312962 238046 313018 238102
rect 313086 238046 313142 238102
rect 312714 237922 312770 237978
rect 312838 237922 312894 237978
rect 312962 237922 313018 237978
rect 313086 237922 313142 237978
rect 285714 226294 285770 226350
rect 285838 226294 285894 226350
rect 285962 226294 286018 226350
rect 286086 226294 286142 226350
rect 285714 226170 285770 226226
rect 285838 226170 285894 226226
rect 285962 226170 286018 226226
rect 286086 226170 286142 226226
rect 285714 226046 285770 226102
rect 285838 226046 285894 226102
rect 285962 226046 286018 226102
rect 286086 226046 286142 226102
rect 285714 225922 285770 225978
rect 285838 225922 285894 225978
rect 285962 225922 286018 225978
rect 286086 225922 286142 225978
rect 289772 214442 289828 214498
rect 285714 208294 285770 208350
rect 285838 208294 285894 208350
rect 285962 208294 286018 208350
rect 286086 208294 286142 208350
rect 285714 208170 285770 208226
rect 285838 208170 285894 208226
rect 285962 208170 286018 208226
rect 286086 208170 286142 208226
rect 285714 208046 285770 208102
rect 285838 208046 285894 208102
rect 285962 208046 286018 208102
rect 286086 208046 286142 208102
rect 285714 207922 285770 207978
rect 285838 207922 285894 207978
rect 285962 207922 286018 207978
rect 286086 207922 286142 207978
rect 285714 190294 285770 190350
rect 285838 190294 285894 190350
rect 285962 190294 286018 190350
rect 286086 190294 286142 190350
rect 285714 190170 285770 190226
rect 285838 190170 285894 190226
rect 285962 190170 286018 190226
rect 286086 190170 286142 190226
rect 285714 190046 285770 190102
rect 285838 190046 285894 190102
rect 285962 190046 286018 190102
rect 286086 190046 286142 190102
rect 285714 189922 285770 189978
rect 285838 189922 285894 189978
rect 285962 189922 286018 189978
rect 286086 189922 286142 189978
rect 285714 172294 285770 172350
rect 285838 172294 285894 172350
rect 285962 172294 286018 172350
rect 286086 172294 286142 172350
rect 285714 172170 285770 172226
rect 285838 172170 285894 172226
rect 285962 172170 286018 172226
rect 286086 172170 286142 172226
rect 285714 172046 285770 172102
rect 285838 172046 285894 172102
rect 285962 172046 286018 172102
rect 286086 172046 286142 172102
rect 285714 171922 285770 171978
rect 285838 171922 285894 171978
rect 285962 171922 286018 171978
rect 286086 171922 286142 171978
rect 285714 154294 285770 154350
rect 285838 154294 285894 154350
rect 285962 154294 286018 154350
rect 286086 154294 286142 154350
rect 285714 154170 285770 154226
rect 285838 154170 285894 154226
rect 285962 154170 286018 154226
rect 286086 154170 286142 154226
rect 285714 154046 285770 154102
rect 285838 154046 285894 154102
rect 285962 154046 286018 154102
rect 286086 154046 286142 154102
rect 285714 153922 285770 153978
rect 285838 153922 285894 153978
rect 285962 153922 286018 153978
rect 286086 153922 286142 153978
rect 285714 136294 285770 136350
rect 285838 136294 285894 136350
rect 285962 136294 286018 136350
rect 286086 136294 286142 136350
rect 285714 136170 285770 136226
rect 285838 136170 285894 136226
rect 285962 136170 286018 136226
rect 286086 136170 286142 136226
rect 285714 136046 285770 136102
rect 285838 136046 285894 136102
rect 285962 136046 286018 136102
rect 286086 136046 286142 136102
rect 285714 135922 285770 135978
rect 285838 135922 285894 135978
rect 285962 135922 286018 135978
rect 286086 135922 286142 135978
rect 285714 118294 285770 118350
rect 285838 118294 285894 118350
rect 285962 118294 286018 118350
rect 286086 118294 286142 118350
rect 285714 118170 285770 118226
rect 285838 118170 285894 118226
rect 285962 118170 286018 118226
rect 286086 118170 286142 118226
rect 285714 118046 285770 118102
rect 285838 118046 285894 118102
rect 285962 118046 286018 118102
rect 286086 118046 286142 118102
rect 285714 117922 285770 117978
rect 285838 117922 285894 117978
rect 285962 117922 286018 117978
rect 286086 117922 286142 117978
rect 285714 100294 285770 100350
rect 285838 100294 285894 100350
rect 285962 100294 286018 100350
rect 286086 100294 286142 100350
rect 285714 100170 285770 100226
rect 285838 100170 285894 100226
rect 285962 100170 286018 100226
rect 286086 100170 286142 100226
rect 285714 100046 285770 100102
rect 285838 100046 285894 100102
rect 285962 100046 286018 100102
rect 286086 100046 286142 100102
rect 285714 99922 285770 99978
rect 285838 99922 285894 99978
rect 285962 99922 286018 99978
rect 286086 99922 286142 99978
rect 285714 82294 285770 82350
rect 285838 82294 285894 82350
rect 285962 82294 286018 82350
rect 286086 82294 286142 82350
rect 285714 82170 285770 82226
rect 285838 82170 285894 82226
rect 285962 82170 286018 82226
rect 286086 82170 286142 82226
rect 285714 82046 285770 82102
rect 285838 82046 285894 82102
rect 285962 82046 286018 82102
rect 286086 82046 286142 82102
rect 285714 81922 285770 81978
rect 285838 81922 285894 81978
rect 285962 81922 286018 81978
rect 286086 81922 286142 81978
rect 285714 64294 285770 64350
rect 285838 64294 285894 64350
rect 285962 64294 286018 64350
rect 286086 64294 286142 64350
rect 285714 64170 285770 64226
rect 285838 64170 285894 64226
rect 285962 64170 286018 64226
rect 286086 64170 286142 64226
rect 285714 64046 285770 64102
rect 285838 64046 285894 64102
rect 285962 64046 286018 64102
rect 286086 64046 286142 64102
rect 285714 63922 285770 63978
rect 285838 63922 285894 63978
rect 285962 63922 286018 63978
rect 286086 63922 286142 63978
rect 285714 46294 285770 46350
rect 285838 46294 285894 46350
rect 285962 46294 286018 46350
rect 286086 46294 286142 46350
rect 285714 46170 285770 46226
rect 285838 46170 285894 46226
rect 285962 46170 286018 46226
rect 286086 46170 286142 46226
rect 285714 46046 285770 46102
rect 285838 46046 285894 46102
rect 285962 46046 286018 46102
rect 286086 46046 286142 46102
rect 285714 45922 285770 45978
rect 285838 45922 285894 45978
rect 285962 45922 286018 45978
rect 286086 45922 286142 45978
rect 285714 28294 285770 28350
rect 285838 28294 285894 28350
rect 285962 28294 286018 28350
rect 286086 28294 286142 28350
rect 285714 28170 285770 28226
rect 285838 28170 285894 28226
rect 285962 28170 286018 28226
rect 286086 28170 286142 28226
rect 285714 28046 285770 28102
rect 285838 28046 285894 28102
rect 285962 28046 286018 28102
rect 286086 28046 286142 28102
rect 285714 27922 285770 27978
rect 285838 27922 285894 27978
rect 285962 27922 286018 27978
rect 286086 27922 286142 27978
rect 285714 10294 285770 10350
rect 285838 10294 285894 10350
rect 285962 10294 286018 10350
rect 286086 10294 286142 10350
rect 285714 10170 285770 10226
rect 285838 10170 285894 10226
rect 285962 10170 286018 10226
rect 286086 10170 286142 10226
rect 285714 10046 285770 10102
rect 285838 10046 285894 10102
rect 285962 10046 286018 10102
rect 286086 10046 286142 10102
rect 285714 9922 285770 9978
rect 285838 9922 285894 9978
rect 285962 9922 286018 9978
rect 286086 9922 286142 9978
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 288092 211382 288148 211438
rect 293804 160442 293860 160498
rect 293916 158642 293972 158698
rect 295596 155402 295652 155458
rect 298956 160622 299012 160678
rect 300636 158822 300692 158878
rect 298172 124262 298228 124318
rect 304892 124082 304948 124138
rect 306572 123902 306628 123958
rect 311612 231002 311668 231058
rect 307356 146042 307412 146098
rect 306796 123542 306852 123598
rect 299528 82091 299584 82147
rect 299632 82091 299688 82147
rect 299736 82091 299792 82147
rect 299528 81987 299584 82043
rect 299632 81987 299688 82043
rect 299736 81987 299792 82043
rect 299528 81883 299584 81939
rect 299632 81883 299688 81939
rect 299736 81883 299792 81939
rect 295412 76294 295468 76350
rect 295536 76294 295592 76350
rect 295412 76170 295468 76226
rect 295536 76170 295592 76226
rect 295412 76046 295468 76102
rect 295536 76046 295592 76102
rect 295412 75922 295468 75978
rect 295536 75922 295592 75978
rect 303728 76294 303784 76350
rect 303852 76294 303908 76350
rect 303728 76170 303784 76226
rect 303852 76170 303908 76226
rect 303728 76046 303784 76102
rect 303852 76046 303908 76102
rect 303728 75922 303784 75978
rect 303852 75922 303908 75978
rect 299570 64294 299626 64350
rect 299694 64294 299750 64350
rect 299570 64170 299626 64226
rect 299694 64170 299750 64226
rect 299570 64046 299626 64102
rect 299694 64046 299750 64102
rect 299570 63922 299626 63978
rect 299694 63922 299750 63978
rect 295412 58294 295468 58350
rect 295536 58294 295592 58350
rect 295412 58170 295468 58226
rect 295536 58170 295592 58226
rect 295412 58046 295468 58102
rect 295536 58046 295592 58102
rect 295412 57922 295468 57978
rect 295536 57922 295592 57978
rect 303728 58294 303784 58350
rect 303852 58294 303908 58350
rect 303728 58170 303784 58226
rect 303852 58170 303908 58226
rect 303728 58046 303784 58102
rect 303852 58046 303908 58102
rect 303728 57922 303784 57978
rect 303852 57922 303908 57978
rect 308252 123722 308308 123778
rect 307844 82091 307900 82147
rect 307948 82091 308004 82147
rect 308052 82091 308108 82147
rect 307844 81987 307900 82043
rect 307948 81987 308004 82043
rect 308052 81987 308108 82043
rect 307844 81883 307900 81939
rect 307948 81883 308004 81939
rect 308052 81883 308108 81939
rect 307886 64294 307942 64350
rect 308010 64294 308066 64350
rect 307886 64170 307942 64226
rect 308010 64170 308066 64226
rect 307886 64046 307942 64102
rect 308010 64046 308066 64102
rect 307886 63922 307942 63978
rect 308010 63922 308066 63978
rect 311724 47762 311780 47818
rect 311836 230642 311892 230698
rect 312060 230462 312116 230518
rect 312044 76294 312100 76350
rect 312168 76294 312224 76350
rect 312044 76170 312100 76226
rect 312168 76170 312224 76226
rect 312044 76046 312100 76102
rect 312168 76046 312224 76102
rect 312044 75922 312100 75978
rect 312168 75922 312224 75978
rect 312044 58294 312100 58350
rect 312168 58294 312224 58350
rect 312044 58170 312100 58226
rect 312168 58170 312224 58226
rect 312044 58046 312100 58102
rect 312168 58046 312224 58102
rect 312044 57922 312100 57978
rect 312168 57922 312224 57978
rect 312396 47942 312452 47998
rect 312714 220294 312770 220350
rect 312838 220294 312894 220350
rect 312962 220294 313018 220350
rect 313086 220294 313142 220350
rect 312714 220170 312770 220226
rect 312838 220170 312894 220226
rect 312962 220170 313018 220226
rect 313086 220170 313142 220226
rect 312714 220046 312770 220102
rect 312838 220046 312894 220102
rect 312962 220046 313018 220102
rect 313086 220046 313142 220102
rect 312714 219922 312770 219978
rect 312838 219922 312894 219978
rect 312962 219922 313018 219978
rect 313086 219922 313142 219978
rect 312714 202294 312770 202350
rect 312838 202294 312894 202350
rect 312962 202294 313018 202350
rect 313086 202294 313142 202350
rect 312714 202170 312770 202226
rect 312838 202170 312894 202226
rect 312962 202170 313018 202226
rect 313086 202170 313142 202226
rect 312714 202046 312770 202102
rect 312838 202046 312894 202102
rect 312962 202046 313018 202102
rect 313086 202046 313142 202102
rect 312714 201922 312770 201978
rect 312838 201922 312894 201978
rect 312962 201922 313018 201978
rect 313086 201922 313142 201978
rect 312714 184294 312770 184350
rect 312838 184294 312894 184350
rect 312962 184294 313018 184350
rect 313086 184294 313142 184350
rect 312714 184170 312770 184226
rect 312838 184170 312894 184226
rect 312962 184170 313018 184226
rect 313086 184170 313142 184226
rect 312714 184046 312770 184102
rect 312838 184046 312894 184102
rect 312962 184046 313018 184102
rect 313086 184046 313142 184102
rect 312714 183922 312770 183978
rect 312838 183922 312894 183978
rect 312962 183922 313018 183978
rect 313086 183922 313142 183978
rect 312714 166294 312770 166350
rect 312838 166294 312894 166350
rect 312962 166294 313018 166350
rect 313086 166294 313142 166350
rect 312714 166170 312770 166226
rect 312838 166170 312894 166226
rect 312962 166170 313018 166226
rect 313086 166170 313142 166226
rect 312714 166046 312770 166102
rect 312838 166046 312894 166102
rect 312962 166046 313018 166102
rect 313086 166046 313142 166102
rect 312714 165922 312770 165978
rect 312838 165922 312894 165978
rect 312962 165922 313018 165978
rect 313086 165922 313142 165978
rect 314972 234602 315028 234658
rect 312714 148294 312770 148350
rect 312838 148294 312894 148350
rect 312962 148294 313018 148350
rect 313086 148294 313142 148350
rect 312714 148170 312770 148226
rect 312838 148170 312894 148226
rect 312962 148170 313018 148226
rect 313086 148170 313142 148226
rect 312714 148046 312770 148102
rect 312838 148046 312894 148102
rect 312962 148046 313018 148102
rect 313086 148046 313142 148102
rect 312714 147922 312770 147978
rect 312838 147922 312894 147978
rect 312962 147922 313018 147978
rect 313086 147922 313142 147978
rect 312714 130294 312770 130350
rect 312838 130294 312894 130350
rect 312962 130294 313018 130350
rect 313086 130294 313142 130350
rect 312714 130170 312770 130226
rect 312838 130170 312894 130226
rect 312962 130170 313018 130226
rect 313086 130170 313142 130226
rect 312714 130046 312770 130102
rect 312838 130046 312894 130102
rect 312962 130046 313018 130102
rect 313086 130046 313142 130102
rect 312714 129922 312770 129978
rect 312838 129922 312894 129978
rect 312962 129922 313018 129978
rect 313086 129922 313142 129978
rect 312714 112294 312770 112350
rect 312838 112294 312894 112350
rect 312962 112294 313018 112350
rect 313086 112294 313142 112350
rect 312714 112170 312770 112226
rect 312838 112170 312894 112226
rect 312962 112170 313018 112226
rect 313086 112170 313142 112226
rect 312714 112046 312770 112102
rect 312838 112046 312894 112102
rect 312962 112046 313018 112102
rect 313086 112046 313142 112102
rect 312714 111922 312770 111978
rect 312838 111922 312894 111978
rect 312962 111922 313018 111978
rect 313086 111922 313142 111978
rect 312714 94294 312770 94350
rect 312838 94294 312894 94350
rect 312962 94294 313018 94350
rect 313086 94294 313142 94350
rect 312714 94170 312770 94226
rect 312838 94170 312894 94226
rect 312962 94170 313018 94226
rect 313086 94170 313142 94226
rect 312714 94046 312770 94102
rect 312838 94046 312894 94102
rect 312962 94046 313018 94102
rect 313086 94046 313142 94102
rect 312714 93922 312770 93978
rect 312838 93922 312894 93978
rect 312962 93922 313018 93978
rect 313086 93922 313142 93978
rect 312714 76294 312770 76350
rect 312838 76294 312894 76350
rect 312962 76294 313018 76350
rect 313086 76294 313142 76350
rect 312714 76170 312770 76226
rect 312838 76170 312894 76226
rect 312962 76170 313018 76226
rect 313086 76170 313142 76226
rect 312714 76046 312770 76102
rect 312838 76046 312894 76102
rect 312962 76046 313018 76102
rect 313086 76046 313142 76102
rect 312714 75922 312770 75978
rect 312838 75922 312894 75978
rect 312962 75922 313018 75978
rect 313086 75922 313142 75978
rect 312714 58294 312770 58350
rect 312838 58294 312894 58350
rect 312962 58294 313018 58350
rect 313086 58294 313142 58350
rect 312714 58170 312770 58226
rect 312838 58170 312894 58226
rect 312962 58170 313018 58226
rect 313086 58170 313142 58226
rect 312714 58046 312770 58102
rect 312838 58046 312894 58102
rect 312962 58046 313018 58102
rect 313086 58046 313142 58102
rect 312714 57922 312770 57978
rect 312838 57922 312894 57978
rect 312962 57922 313018 57978
rect 313086 57922 313142 57978
rect 312714 40294 312770 40350
rect 312838 40294 312894 40350
rect 312962 40294 313018 40350
rect 313086 40294 313142 40350
rect 312714 40170 312770 40226
rect 312838 40170 312894 40226
rect 312962 40170 313018 40226
rect 313086 40170 313142 40226
rect 312714 40046 312770 40102
rect 312838 40046 312894 40102
rect 312962 40046 313018 40102
rect 313086 40046 313142 40102
rect 312714 39922 312770 39978
rect 312838 39922 312894 39978
rect 312962 39922 313018 39978
rect 313086 39922 313142 39978
rect 312714 22294 312770 22350
rect 312838 22294 312894 22350
rect 312962 22294 313018 22350
rect 313086 22294 313142 22350
rect 312714 22170 312770 22226
rect 312838 22170 312894 22226
rect 312962 22170 313018 22226
rect 313086 22170 313142 22226
rect 312714 22046 312770 22102
rect 312838 22046 312894 22102
rect 312962 22046 313018 22102
rect 313086 22046 313142 22102
rect 312714 21922 312770 21978
rect 312838 21922 312894 21978
rect 312962 21922 313018 21978
rect 313086 21922 313142 21978
rect 285714 -1176 285770 -1120
rect 285838 -1176 285894 -1120
rect 285962 -1176 286018 -1120
rect 286086 -1176 286142 -1120
rect 285714 -1300 285770 -1244
rect 285838 -1300 285894 -1244
rect 285962 -1300 286018 -1244
rect 286086 -1300 286142 -1244
rect 285714 -1424 285770 -1368
rect 285838 -1424 285894 -1368
rect 285962 -1424 286018 -1368
rect 286086 -1424 286142 -1368
rect 285714 -1548 285770 -1492
rect 285838 -1548 285894 -1492
rect 285962 -1548 286018 -1492
rect 286086 -1548 286142 -1492
rect 315084 211202 315140 211258
rect 334236 241982 334292 242038
rect 335916 240722 335972 240778
rect 334124 240542 334180 240598
rect 320572 240212 320628 240238
rect 320572 240182 320628 240212
rect 319900 240044 319956 240058
rect 319900 240002 319956 240044
rect 316434 226294 316490 226350
rect 316558 226294 316614 226350
rect 316682 226294 316738 226350
rect 316806 226294 316862 226350
rect 316434 226170 316490 226226
rect 316558 226170 316614 226226
rect 316682 226170 316738 226226
rect 316806 226170 316862 226226
rect 316434 226046 316490 226102
rect 316558 226046 316614 226102
rect 316682 226046 316738 226102
rect 316806 226046 316862 226102
rect 316434 225922 316490 225978
rect 316558 225922 316614 225978
rect 316682 225922 316738 225978
rect 316806 225922 316862 225978
rect 316434 208294 316490 208350
rect 316558 208294 316614 208350
rect 316682 208294 316738 208350
rect 316806 208294 316862 208350
rect 316434 208170 316490 208226
rect 316558 208170 316614 208226
rect 316682 208170 316738 208226
rect 316806 208170 316862 208226
rect 316434 208046 316490 208102
rect 316558 208046 316614 208102
rect 316682 208046 316738 208102
rect 316806 208046 316862 208102
rect 316434 207922 316490 207978
rect 316558 207922 316614 207978
rect 316682 207922 316738 207978
rect 316806 207922 316862 207978
rect 315538 184294 315594 184350
rect 315662 184294 315718 184350
rect 315538 184170 315594 184226
rect 315662 184170 315718 184226
rect 315538 184046 315594 184102
rect 315662 184046 315718 184102
rect 315538 183922 315594 183978
rect 315662 183922 315718 183978
rect 315538 166294 315594 166350
rect 315662 166294 315718 166350
rect 315538 166170 315594 166226
rect 315662 166170 315718 166226
rect 315538 166046 315594 166102
rect 315662 166046 315718 166102
rect 315538 165922 315594 165978
rect 315662 165922 315718 165978
rect 321244 237662 321300 237718
rect 321916 237482 321972 237538
rect 320012 230642 320068 230698
rect 329196 230282 329252 230338
rect 336700 304802 336756 304858
rect 336588 241622 336644 241678
rect 338268 368702 338324 368758
rect 336924 308942 336980 308998
rect 338156 336302 338212 336358
rect 336812 252962 336868 253018
rect 336924 284642 336980 284698
rect 336812 241802 336868 241858
rect 337260 279602 337316 279658
rect 337036 277262 337092 277318
rect 337148 267182 337204 267238
rect 337260 253502 337316 253558
rect 337372 257822 337428 257878
rect 337260 244682 337316 244738
rect 337484 254762 337540 254818
rect 337596 246302 337652 246358
rect 337708 240362 337764 240418
rect 337484 234602 337540 234658
rect 343434 400294 343490 400350
rect 343558 400294 343614 400350
rect 343682 400294 343738 400350
rect 343806 400294 343862 400350
rect 343434 400170 343490 400226
rect 343558 400170 343614 400226
rect 343682 400170 343738 400226
rect 343806 400170 343862 400226
rect 343434 400046 343490 400102
rect 343558 400046 343614 400102
rect 343682 400046 343738 400102
rect 343806 400046 343862 400102
rect 343434 399922 343490 399978
rect 343558 399922 343614 399978
rect 343682 399922 343738 399978
rect 343806 399922 343862 399978
rect 341964 392282 342020 392338
rect 338828 313262 338884 313318
rect 339388 336302 339444 336358
rect 339388 313292 339444 313318
rect 339388 313262 339444 313292
rect 339276 305004 339332 305038
rect 339276 304982 339332 305004
rect 339388 284642 339444 284698
rect 339388 279636 339444 279658
rect 339388 279602 339444 279636
rect 339276 277262 339332 277318
rect 339276 267372 339332 267418
rect 339276 267362 339332 267372
rect 338716 264302 338772 264358
rect 338380 254582 338436 254638
rect 338604 258722 338660 258778
rect 338268 248642 338324 248698
rect 338380 239282 338436 239338
rect 339388 264302 339444 264358
rect 338828 255662 338884 255718
rect 338940 248822 338996 248878
rect 339052 248642 339108 248698
rect 339276 255662 339332 255718
rect 339276 254762 339332 254818
rect 339276 254582 339332 254638
rect 339500 258748 339556 258778
rect 339500 258722 339556 258748
rect 339500 257852 339556 257878
rect 339500 257822 339556 257852
rect 339276 248822 339332 248878
rect 339388 246316 339444 246358
rect 339388 246302 339444 246316
rect 339500 241802 339556 241858
rect 339724 227582 339780 227638
rect 340284 373742 340340 373798
rect 341180 244682 341236 244738
rect 340396 241622 340452 241678
rect 341516 224162 341572 224218
rect 341740 234242 341796 234298
rect 339948 193922 340004 193978
rect 339276 193202 339332 193258
rect 342076 373022 342132 373078
rect 342300 325862 342356 325918
rect 342860 378782 342916 378838
rect 342748 292562 342804 292618
rect 356188 408122 356244 408178
rect 358764 409922 358820 409978
rect 357308 409562 357364 409618
rect 358092 409382 358148 409438
rect 357644 409022 357700 409078
rect 357644 407582 357700 407638
rect 347154 406294 347210 406350
rect 347278 406294 347334 406350
rect 347402 406294 347458 406350
rect 347526 406294 347582 406350
rect 347154 406170 347210 406226
rect 347278 406170 347334 406226
rect 347402 406170 347458 406226
rect 347526 406170 347582 406226
rect 347154 406046 347210 406102
rect 347278 406046 347334 406102
rect 347402 406046 347458 406102
rect 347526 406046 347582 406102
rect 347154 405922 347210 405978
rect 347278 405922 347334 405978
rect 347402 405922 347458 405978
rect 347526 405922 347582 405978
rect 343434 382294 343490 382350
rect 343558 382294 343614 382350
rect 343682 382294 343738 382350
rect 343806 382294 343862 382350
rect 343434 382170 343490 382226
rect 343558 382170 343614 382226
rect 343682 382170 343738 382226
rect 343806 382170 343862 382226
rect 343434 382046 343490 382102
rect 343558 382046 343614 382102
rect 343682 382046 343738 382102
rect 343806 382046 343862 382102
rect 343434 381922 343490 381978
rect 343558 381922 343614 381978
rect 343682 381922 343738 381978
rect 343806 381922 343862 381978
rect 344092 398222 344148 398278
rect 345548 396602 345604 396658
rect 344204 395342 344260 395398
rect 343434 364294 343490 364350
rect 343558 364294 343614 364350
rect 343682 364294 343738 364350
rect 343806 364294 343862 364350
rect 343434 364170 343490 364226
rect 343558 364170 343614 364226
rect 343682 364170 343738 364226
rect 343806 364170 343862 364226
rect 343434 364046 343490 364102
rect 343558 364046 343614 364102
rect 343682 364046 343738 364102
rect 343806 364046 343862 364102
rect 343434 363922 343490 363978
rect 343558 363922 343614 363978
rect 343682 363922 343738 363978
rect 343806 363922 343862 363978
rect 343434 346294 343490 346350
rect 343558 346294 343614 346350
rect 343682 346294 343738 346350
rect 343806 346294 343862 346350
rect 343434 346170 343490 346226
rect 343558 346170 343614 346226
rect 343682 346170 343738 346226
rect 343806 346170 343862 346226
rect 343434 346046 343490 346102
rect 343558 346046 343614 346102
rect 343682 346046 343738 346102
rect 343806 346046 343862 346102
rect 343434 345922 343490 345978
rect 343558 345922 343614 345978
rect 343682 345922 343738 345978
rect 343806 345922 343862 345978
rect 344428 366362 344484 366418
rect 343434 328294 343490 328350
rect 343558 328294 343614 328350
rect 343682 328294 343738 328350
rect 343806 328294 343862 328350
rect 343434 328170 343490 328226
rect 343558 328170 343614 328226
rect 343682 328170 343738 328226
rect 343806 328170 343862 328226
rect 343434 328046 343490 328102
rect 343558 328046 343614 328102
rect 343682 328046 343738 328102
rect 343806 328046 343862 328102
rect 343434 327922 343490 327978
rect 343558 327922 343614 327978
rect 343682 327922 343738 327978
rect 343806 327922 343862 327978
rect 343434 310294 343490 310350
rect 343558 310294 343614 310350
rect 343682 310294 343738 310350
rect 343806 310294 343862 310350
rect 343434 310170 343490 310226
rect 343558 310170 343614 310226
rect 343682 310170 343738 310226
rect 343806 310170 343862 310226
rect 343434 310046 343490 310102
rect 343558 310046 343614 310102
rect 343682 310046 343738 310102
rect 343806 310046 343862 310102
rect 343434 309922 343490 309978
rect 343558 309922 343614 309978
rect 343682 309922 343738 309978
rect 343806 309922 343862 309978
rect 343434 292294 343490 292350
rect 343558 292294 343614 292350
rect 343682 292294 343738 292350
rect 343806 292294 343862 292350
rect 343434 292170 343490 292226
rect 343558 292170 343614 292226
rect 343682 292170 343738 292226
rect 343806 292170 343862 292226
rect 343434 292046 343490 292102
rect 343558 292046 343614 292102
rect 343682 292046 343738 292102
rect 343806 292046 343862 292102
rect 343434 291922 343490 291978
rect 343558 291922 343614 291978
rect 343682 291922 343738 291978
rect 343806 291922 343862 291978
rect 342748 287342 342804 287398
rect 343434 274294 343490 274350
rect 343558 274294 343614 274350
rect 343682 274294 343738 274350
rect 343806 274294 343862 274350
rect 343434 274170 343490 274226
rect 343558 274170 343614 274226
rect 343682 274170 343738 274226
rect 343806 274170 343862 274226
rect 343434 274046 343490 274102
rect 343558 274046 343614 274102
rect 343682 274046 343738 274102
rect 343806 274046 343862 274102
rect 343434 273922 343490 273978
rect 343558 273922 343614 273978
rect 343682 273922 343738 273978
rect 343806 273922 343862 273978
rect 342860 236042 342916 236098
rect 343434 256294 343490 256350
rect 343558 256294 343614 256350
rect 343682 256294 343738 256350
rect 343806 256294 343862 256350
rect 343434 256170 343490 256226
rect 343558 256170 343614 256226
rect 343682 256170 343738 256226
rect 343806 256170 343862 256226
rect 343434 256046 343490 256102
rect 343558 256046 343614 256102
rect 343682 256046 343738 256102
rect 343806 256046 343862 256102
rect 343434 255922 343490 255978
rect 343558 255922 343614 255978
rect 343682 255922 343738 255978
rect 343806 255922 343862 255978
rect 343084 241082 343140 241138
rect 342972 234422 343028 234478
rect 343434 238294 343490 238350
rect 343558 238294 343614 238350
rect 343682 238294 343738 238350
rect 343806 238294 343862 238350
rect 343434 238170 343490 238226
rect 343558 238170 343614 238226
rect 343682 238170 343738 238226
rect 343806 238170 343862 238226
rect 343434 238046 343490 238102
rect 343558 238046 343614 238102
rect 343682 238046 343738 238102
rect 343806 238046 343862 238102
rect 343434 237922 343490 237978
rect 343558 237922 343614 237978
rect 343682 237922 343738 237978
rect 343806 237922 343862 237978
rect 342636 231002 342692 231058
rect 343434 220294 343490 220350
rect 343558 220294 343614 220350
rect 343682 220294 343738 220350
rect 343806 220294 343862 220350
rect 343434 220170 343490 220226
rect 343558 220170 343614 220226
rect 343682 220170 343738 220226
rect 343806 220170 343862 220226
rect 343434 220046 343490 220102
rect 343558 220046 343614 220102
rect 343682 220046 343738 220102
rect 343806 220046 343862 220102
rect 343434 219922 343490 219978
rect 343558 219922 343614 219978
rect 343682 219922 343738 219978
rect 343806 219922 343862 219978
rect 342972 211022 343028 211078
rect 343434 202294 343490 202350
rect 343558 202294 343614 202350
rect 343682 202294 343738 202350
rect 343806 202294 343862 202350
rect 343434 202170 343490 202226
rect 343558 202170 343614 202226
rect 343682 202170 343738 202226
rect 343806 202170 343862 202226
rect 343434 202046 343490 202102
rect 343558 202046 343614 202102
rect 343682 202046 343738 202102
rect 343806 202046 343862 202102
rect 343434 201922 343490 201978
rect 343558 201922 343614 201978
rect 343682 201922 343738 201978
rect 343806 201922 343862 201978
rect 341852 192482 341908 192538
rect 344316 192662 344372 192718
rect 345100 252962 345156 253018
rect 344876 191762 344932 191818
rect 344092 191582 344148 191638
rect 319822 190294 319878 190350
rect 319946 190294 320002 190350
rect 319822 190170 319878 190226
rect 319946 190170 320002 190226
rect 319822 190046 319878 190102
rect 319946 190046 320002 190102
rect 319822 189922 319878 189978
rect 319946 189922 320002 189978
rect 328390 190294 328446 190350
rect 328514 190294 328570 190350
rect 328390 190170 328446 190226
rect 328514 190170 328570 190226
rect 328390 190046 328446 190102
rect 328514 190046 328570 190102
rect 328390 189922 328446 189978
rect 328514 189922 328570 189978
rect 336958 190294 337014 190350
rect 337082 190294 337138 190350
rect 336958 190170 337014 190226
rect 337082 190170 337138 190226
rect 336958 190046 337014 190102
rect 337082 190046 337138 190102
rect 336958 189922 337014 189978
rect 337082 189922 337138 189978
rect 324106 184294 324162 184350
rect 324230 184294 324286 184350
rect 324106 184170 324162 184226
rect 324230 184170 324286 184226
rect 324106 184046 324162 184102
rect 324230 184046 324286 184102
rect 324106 183922 324162 183978
rect 324230 183922 324286 183978
rect 332674 184294 332730 184350
rect 332798 184294 332854 184350
rect 332674 184170 332730 184226
rect 332798 184170 332854 184226
rect 332674 184046 332730 184102
rect 332798 184046 332854 184102
rect 332674 183922 332730 183978
rect 332798 183922 332854 183978
rect 341242 184294 341298 184350
rect 341366 184294 341422 184350
rect 341242 184170 341298 184226
rect 341366 184170 341422 184226
rect 341242 184046 341298 184102
rect 341366 184046 341422 184102
rect 341242 183922 341298 183978
rect 341366 183922 341422 183978
rect 357756 406862 357812 406918
rect 347154 388294 347210 388350
rect 347278 388294 347334 388350
rect 347402 388294 347458 388350
rect 347526 388294 347582 388350
rect 347154 388170 347210 388226
rect 347278 388170 347334 388226
rect 347402 388170 347458 388226
rect 347526 388170 347582 388226
rect 347154 388046 347210 388102
rect 347278 388046 347334 388102
rect 347402 388046 347458 388102
rect 347526 388046 347582 388102
rect 347154 387922 347210 387978
rect 347278 387922 347334 387978
rect 347402 387922 347458 387978
rect 347526 387922 347582 387978
rect 345436 195722 345492 195778
rect 345324 192302 345380 192358
rect 345526 190294 345582 190350
rect 345650 190294 345706 190350
rect 345526 190170 345582 190226
rect 345650 190170 345706 190226
rect 345526 190046 345582 190102
rect 345650 190046 345706 190102
rect 345526 189922 345582 189978
rect 345650 189922 345706 189978
rect 345996 196622 346052 196678
rect 345884 175202 345940 175258
rect 345212 173942 345268 173998
rect 319822 172294 319878 172350
rect 319946 172294 320002 172350
rect 319822 172170 319878 172226
rect 319946 172170 320002 172226
rect 319822 172046 319878 172102
rect 319946 172046 320002 172102
rect 319822 171922 319878 171978
rect 319946 171922 320002 171978
rect 328390 172294 328446 172350
rect 328514 172294 328570 172350
rect 328390 172170 328446 172226
rect 328514 172170 328570 172226
rect 328390 172046 328446 172102
rect 328514 172046 328570 172102
rect 328390 171922 328446 171978
rect 328514 171922 328570 171978
rect 336958 172294 337014 172350
rect 337082 172294 337138 172350
rect 336958 172170 337014 172226
rect 337082 172170 337138 172226
rect 336958 172046 337014 172102
rect 337082 172046 337138 172102
rect 336958 171922 337014 171978
rect 337082 171922 337138 171978
rect 345526 172294 345582 172350
rect 345650 172294 345706 172350
rect 345526 172170 345582 172226
rect 345650 172170 345706 172226
rect 345526 172046 345582 172102
rect 345650 172046 345706 172102
rect 345526 171922 345582 171978
rect 345650 171922 345706 171978
rect 324106 166294 324162 166350
rect 324230 166294 324286 166350
rect 324106 166170 324162 166226
rect 324230 166170 324286 166226
rect 324106 166046 324162 166102
rect 324230 166046 324286 166102
rect 324106 165922 324162 165978
rect 324230 165922 324286 165978
rect 332674 166294 332730 166350
rect 332798 166294 332854 166350
rect 332674 166170 332730 166226
rect 332798 166170 332854 166226
rect 332674 166046 332730 166102
rect 332798 166046 332854 166102
rect 332674 165922 332730 165978
rect 332798 165922 332854 165978
rect 341242 166294 341298 166350
rect 341366 166294 341422 166350
rect 341242 166170 341298 166226
rect 341366 166170 341422 166226
rect 341242 166046 341298 166102
rect 341366 166046 341422 166102
rect 341242 165922 341298 165978
rect 341366 165922 341422 165978
rect 324380 157742 324436 157798
rect 330652 157562 330708 157618
rect 332220 157382 332276 157438
rect 316434 154294 316490 154350
rect 316558 154294 316614 154350
rect 316682 154294 316738 154350
rect 316806 154294 316862 154350
rect 316434 154170 316490 154226
rect 316558 154170 316614 154226
rect 316682 154170 316738 154226
rect 316806 154170 316862 154226
rect 316434 154046 316490 154102
rect 316558 154046 316614 154102
rect 316682 154046 316738 154102
rect 316806 154046 316862 154102
rect 316434 153922 316490 153978
rect 316558 153922 316614 153978
rect 316682 153922 316738 153978
rect 316806 153922 316862 153978
rect 347154 370294 347210 370350
rect 347278 370294 347334 370350
rect 347402 370294 347458 370350
rect 347526 370294 347582 370350
rect 347154 370170 347210 370226
rect 347278 370170 347334 370226
rect 347402 370170 347458 370226
rect 347526 370170 347582 370226
rect 347154 370046 347210 370102
rect 347278 370046 347334 370102
rect 347402 370046 347458 370102
rect 347526 370046 347582 370102
rect 347154 369922 347210 369978
rect 347278 369922 347334 369978
rect 347402 369922 347458 369978
rect 347526 369922 347582 369978
rect 347154 352294 347210 352350
rect 347278 352294 347334 352350
rect 347402 352294 347458 352350
rect 347526 352294 347582 352350
rect 347154 352170 347210 352226
rect 347278 352170 347334 352226
rect 347402 352170 347458 352226
rect 347526 352170 347582 352226
rect 347154 352046 347210 352102
rect 347278 352046 347334 352102
rect 347402 352046 347458 352102
rect 347526 352046 347582 352102
rect 347154 351922 347210 351978
rect 347278 351922 347334 351978
rect 347402 351922 347458 351978
rect 347526 351922 347582 351978
rect 347154 334294 347210 334350
rect 347278 334294 347334 334350
rect 347402 334294 347458 334350
rect 347526 334294 347582 334350
rect 347154 334170 347210 334226
rect 347278 334170 347334 334226
rect 347402 334170 347458 334226
rect 347526 334170 347582 334226
rect 347154 334046 347210 334102
rect 347278 334046 347334 334102
rect 347402 334046 347458 334102
rect 347526 334046 347582 334102
rect 347154 333922 347210 333978
rect 347278 333922 347334 333978
rect 347402 333922 347458 333978
rect 347526 333922 347582 333978
rect 346220 243062 346276 243118
rect 346332 193202 346388 193258
rect 346108 157562 346164 157618
rect 346220 191582 346276 191638
rect 347154 316294 347210 316350
rect 347278 316294 347334 316350
rect 347402 316294 347458 316350
rect 347526 316294 347582 316350
rect 347154 316170 347210 316226
rect 347278 316170 347334 316226
rect 347402 316170 347458 316226
rect 347526 316170 347582 316226
rect 347154 316046 347210 316102
rect 347278 316046 347334 316102
rect 347402 316046 347458 316102
rect 347526 316046 347582 316102
rect 347154 315922 347210 315978
rect 347278 315922 347334 315978
rect 347402 315922 347458 315978
rect 347526 315922 347582 315978
rect 347154 298294 347210 298350
rect 347278 298294 347334 298350
rect 347402 298294 347458 298350
rect 347526 298294 347582 298350
rect 347154 298170 347210 298226
rect 347278 298170 347334 298226
rect 347402 298170 347458 298226
rect 347526 298170 347582 298226
rect 347154 298046 347210 298102
rect 347278 298046 347334 298102
rect 347402 298046 347458 298102
rect 347526 298046 347582 298102
rect 347154 297922 347210 297978
rect 347278 297922 347334 297978
rect 347402 297922 347458 297978
rect 347526 297922 347582 297978
rect 343434 148294 343490 148350
rect 343558 148294 343614 148350
rect 343682 148294 343738 148350
rect 343806 148294 343862 148350
rect 343434 148170 343490 148226
rect 343558 148170 343614 148226
rect 343682 148170 343738 148226
rect 343806 148170 343862 148226
rect 343434 148046 343490 148102
rect 343558 148046 343614 148102
rect 343682 148046 343738 148102
rect 343806 148046 343862 148102
rect 343434 147922 343490 147978
rect 343558 147922 343614 147978
rect 343682 147922 343738 147978
rect 343806 147922 343862 147978
rect 316434 136294 316490 136350
rect 316558 136294 316614 136350
rect 316682 136294 316738 136350
rect 316806 136294 316862 136350
rect 316434 136170 316490 136226
rect 316558 136170 316614 136226
rect 316682 136170 316738 136226
rect 316806 136170 316862 136226
rect 316434 136046 316490 136102
rect 316558 136046 316614 136102
rect 316682 136046 316738 136102
rect 316806 136046 316862 136102
rect 316434 135922 316490 135978
rect 316558 135922 316614 135978
rect 316682 135922 316738 135978
rect 316806 135922 316862 135978
rect 316434 118294 316490 118350
rect 316558 118294 316614 118350
rect 316682 118294 316738 118350
rect 316806 118294 316862 118350
rect 316434 118170 316490 118226
rect 316558 118170 316614 118226
rect 316682 118170 316738 118226
rect 316806 118170 316862 118226
rect 316434 118046 316490 118102
rect 316558 118046 316614 118102
rect 316682 118046 316738 118102
rect 316806 118046 316862 118102
rect 316434 117922 316490 117978
rect 316558 117922 316614 117978
rect 316682 117922 316738 117978
rect 316806 117922 316862 117978
rect 316434 100294 316490 100350
rect 316558 100294 316614 100350
rect 316682 100294 316738 100350
rect 316806 100294 316862 100350
rect 316434 100170 316490 100226
rect 316558 100170 316614 100226
rect 316682 100170 316738 100226
rect 316806 100170 316862 100226
rect 316434 100046 316490 100102
rect 316558 100046 316614 100102
rect 316682 100046 316738 100102
rect 316806 100046 316862 100102
rect 316434 99922 316490 99978
rect 316558 99922 316614 99978
rect 316682 99922 316738 99978
rect 316806 99922 316862 99978
rect 330092 146942 330148 146998
rect 343434 130294 343490 130350
rect 343558 130294 343614 130350
rect 343682 130294 343738 130350
rect 343806 130294 343862 130350
rect 343434 130170 343490 130226
rect 343558 130170 343614 130226
rect 343682 130170 343738 130226
rect 343806 130170 343862 130226
rect 343434 130046 343490 130102
rect 343558 130046 343614 130102
rect 343682 130046 343738 130102
rect 343806 130046 343862 130102
rect 343434 129922 343490 129978
rect 343558 129922 343614 129978
rect 343682 129922 343738 129978
rect 343806 129922 343862 129978
rect 347154 280294 347210 280350
rect 347278 280294 347334 280350
rect 347402 280294 347458 280350
rect 347526 280294 347582 280350
rect 347154 280170 347210 280226
rect 347278 280170 347334 280226
rect 347402 280170 347458 280226
rect 347526 280170 347582 280226
rect 347154 280046 347210 280102
rect 347278 280046 347334 280102
rect 347402 280046 347458 280102
rect 347526 280046 347582 280102
rect 347154 279922 347210 279978
rect 347278 279922 347334 279978
rect 347402 279922 347458 279978
rect 347526 279922 347582 279978
rect 347154 262294 347210 262350
rect 347278 262294 347334 262350
rect 347402 262294 347458 262350
rect 347526 262294 347582 262350
rect 347154 262170 347210 262226
rect 347278 262170 347334 262226
rect 347402 262170 347458 262226
rect 347526 262170 347582 262226
rect 347154 262046 347210 262102
rect 347278 262046 347334 262102
rect 347402 262046 347458 262102
rect 347526 262046 347582 262102
rect 347154 261922 347210 261978
rect 347278 261922 347334 261978
rect 347402 261922 347458 261978
rect 347526 261922 347582 261978
rect 347154 244294 347210 244350
rect 347278 244294 347334 244350
rect 347402 244294 347458 244350
rect 347526 244294 347582 244350
rect 347154 244170 347210 244226
rect 347278 244170 347334 244226
rect 347402 244170 347458 244226
rect 347526 244170 347582 244226
rect 347154 244046 347210 244102
rect 347278 244046 347334 244102
rect 347402 244046 347458 244102
rect 347526 244046 347582 244102
rect 347154 243922 347210 243978
rect 347278 243922 347334 243978
rect 347402 243922 347458 243978
rect 347526 243922 347582 243978
rect 347154 226294 347210 226350
rect 347278 226294 347334 226350
rect 347402 226294 347458 226350
rect 347526 226294 347582 226350
rect 347154 226170 347210 226226
rect 347278 226170 347334 226226
rect 347402 226170 347458 226226
rect 347526 226170 347582 226226
rect 347154 226046 347210 226102
rect 347278 226046 347334 226102
rect 347402 226046 347458 226102
rect 347526 226046 347582 226102
rect 347154 225922 347210 225978
rect 347278 225922 347334 225978
rect 347402 225922 347458 225978
rect 347526 225922 347582 225978
rect 347154 208294 347210 208350
rect 347278 208294 347334 208350
rect 347402 208294 347458 208350
rect 347526 208294 347582 208350
rect 347154 208170 347210 208226
rect 347278 208170 347334 208226
rect 347402 208170 347458 208226
rect 347526 208170 347582 208226
rect 347154 208046 347210 208102
rect 347278 208046 347334 208102
rect 347402 208046 347458 208102
rect 347526 208046 347582 208102
rect 347154 207922 347210 207978
rect 347278 207922 347334 207978
rect 347402 207922 347458 207978
rect 347526 207922 347582 207978
rect 347004 191762 347060 191818
rect 347004 173762 347060 173818
rect 348572 375362 348628 375418
rect 347788 157382 347844 157438
rect 348460 241982 348516 242038
rect 347154 154294 347210 154350
rect 347278 154294 347334 154350
rect 347402 154294 347458 154350
rect 347526 154294 347582 154350
rect 347154 154170 347210 154226
rect 347278 154170 347334 154226
rect 347402 154170 347458 154226
rect 347526 154170 347582 154226
rect 347154 154046 347210 154102
rect 347278 154046 347334 154102
rect 347402 154046 347458 154102
rect 347526 154046 347582 154102
rect 347154 153922 347210 153978
rect 347278 153922 347334 153978
rect 347402 153922 347458 153978
rect 347526 153922 347582 153978
rect 347154 136294 347210 136350
rect 347278 136294 347334 136350
rect 347402 136294 347458 136350
rect 347526 136294 347582 136350
rect 347154 136170 347210 136226
rect 347278 136170 347334 136226
rect 347402 136170 347458 136226
rect 347526 136170 347582 136226
rect 347154 136046 347210 136102
rect 347278 136046 347334 136102
rect 347402 136046 347458 136102
rect 347526 136046 347582 136102
rect 347154 135922 347210 135978
rect 347278 135922 347334 135978
rect 347402 135922 347458 135978
rect 347526 135922 347582 135978
rect 343434 112294 343490 112350
rect 343558 112294 343614 112350
rect 343682 112294 343738 112350
rect 343806 112294 343862 112350
rect 343434 112170 343490 112226
rect 343558 112170 343614 112226
rect 343682 112170 343738 112226
rect 343806 112170 343862 112226
rect 343434 112046 343490 112102
rect 343558 112046 343614 112102
rect 343682 112046 343738 112102
rect 343806 112046 343862 112102
rect 343434 111922 343490 111978
rect 343558 111922 343614 111978
rect 343682 111922 343738 111978
rect 343806 111922 343862 111978
rect 343434 94294 343490 94350
rect 343558 94294 343614 94350
rect 343682 94294 343738 94350
rect 343806 94294 343862 94350
rect 343434 94170 343490 94226
rect 343558 94170 343614 94226
rect 343682 94170 343738 94226
rect 343806 94170 343862 94226
rect 343434 94046 343490 94102
rect 343558 94046 343614 94102
rect 343682 94046 343738 94102
rect 343806 94046 343862 94102
rect 343434 93922 343490 93978
rect 343558 93922 343614 93978
rect 343682 93922 343738 93978
rect 343806 93922 343862 93978
rect 316160 82091 316216 82147
rect 316264 82091 316320 82147
rect 316368 82091 316424 82147
rect 316160 81987 316216 82043
rect 316264 81987 316320 82043
rect 316368 81987 316424 82043
rect 316160 81883 316216 81939
rect 316264 81883 316320 81939
rect 316368 81883 316424 81939
rect 324476 82091 324532 82147
rect 324580 82091 324636 82147
rect 324684 82091 324740 82147
rect 324476 81987 324532 82043
rect 324580 81987 324636 82043
rect 324684 81987 324740 82043
rect 324476 81883 324532 81939
rect 324580 81883 324636 81939
rect 324684 81883 324740 81939
rect 320360 76294 320416 76350
rect 320484 76294 320540 76350
rect 320360 76170 320416 76226
rect 320484 76170 320540 76226
rect 320360 76046 320416 76102
rect 320484 76046 320540 76102
rect 320360 75922 320416 75978
rect 320484 75922 320540 75978
rect 343434 76294 343490 76350
rect 343558 76294 343614 76350
rect 343682 76294 343738 76350
rect 343806 76294 343862 76350
rect 343434 76170 343490 76226
rect 343558 76170 343614 76226
rect 343682 76170 343738 76226
rect 343806 76170 343862 76226
rect 343434 76046 343490 76102
rect 343558 76046 343614 76102
rect 343682 76046 343738 76102
rect 343806 76046 343862 76102
rect 343434 75922 343490 75978
rect 343558 75922 343614 75978
rect 343682 75922 343738 75978
rect 343806 75922 343862 75978
rect 316202 64294 316258 64350
rect 316326 64294 316382 64350
rect 316202 64170 316258 64226
rect 316326 64170 316382 64226
rect 316202 64046 316258 64102
rect 316326 64046 316382 64102
rect 316202 63922 316258 63978
rect 316326 63922 316382 63978
rect 324518 64294 324574 64350
rect 324642 64294 324698 64350
rect 324518 64170 324574 64226
rect 324642 64170 324698 64226
rect 324518 64046 324574 64102
rect 324642 64046 324698 64102
rect 324518 63922 324574 63978
rect 324642 63922 324698 63978
rect 320360 58294 320416 58350
rect 320484 58294 320540 58350
rect 320360 58170 320416 58226
rect 320484 58170 320540 58226
rect 320360 58046 320416 58102
rect 320484 58046 320540 58102
rect 320360 57922 320416 57978
rect 320484 57922 320540 57978
rect 343434 58294 343490 58350
rect 343558 58294 343614 58350
rect 343682 58294 343738 58350
rect 343806 58294 343862 58350
rect 343434 58170 343490 58226
rect 343558 58170 343614 58226
rect 343682 58170 343738 58226
rect 343806 58170 343862 58226
rect 343434 58046 343490 58102
rect 343558 58046 343614 58102
rect 343682 58046 343738 58102
rect 343806 58046 343862 58102
rect 343434 57922 343490 57978
rect 343558 57922 343614 57978
rect 343682 57922 343738 57978
rect 343806 57922 343862 57978
rect 314972 4922 315028 4978
rect 316434 46294 316490 46350
rect 316558 46294 316614 46350
rect 316682 46294 316738 46350
rect 316806 46294 316862 46350
rect 316434 46170 316490 46226
rect 316558 46170 316614 46226
rect 316682 46170 316738 46226
rect 316806 46170 316862 46226
rect 316434 46046 316490 46102
rect 316558 46046 316614 46102
rect 316682 46046 316738 46102
rect 316806 46046 316862 46102
rect 316434 45922 316490 45978
rect 316558 45922 316614 45978
rect 316682 45922 316738 45978
rect 316806 45922 316862 45978
rect 316434 28294 316490 28350
rect 316558 28294 316614 28350
rect 316682 28294 316738 28350
rect 316806 28294 316862 28350
rect 316434 28170 316490 28226
rect 316558 28170 316614 28226
rect 316682 28170 316738 28226
rect 316806 28170 316862 28226
rect 316434 28046 316490 28102
rect 316558 28046 316614 28102
rect 316682 28046 316738 28102
rect 316806 28046 316862 28102
rect 316434 27922 316490 27978
rect 316558 27922 316614 27978
rect 316682 27922 316738 27978
rect 316806 27922 316862 27978
rect 316434 10294 316490 10350
rect 316558 10294 316614 10350
rect 316682 10294 316738 10350
rect 316806 10294 316862 10350
rect 316434 10170 316490 10226
rect 316558 10170 316614 10226
rect 316682 10170 316738 10226
rect 316806 10170 316862 10226
rect 316434 10046 316490 10102
rect 316558 10046 316614 10102
rect 316682 10046 316738 10102
rect 316806 10046 316862 10102
rect 316434 9922 316490 9978
rect 316558 9922 316614 9978
rect 316682 9922 316738 9978
rect 316806 9922 316862 9978
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 316434 -1176 316490 -1120
rect 316558 -1176 316614 -1120
rect 316682 -1176 316738 -1120
rect 316806 -1176 316862 -1120
rect 316434 -1300 316490 -1244
rect 316558 -1300 316614 -1244
rect 316682 -1300 316738 -1244
rect 316806 -1300 316862 -1244
rect 316434 -1424 316490 -1368
rect 316558 -1424 316614 -1368
rect 316682 -1424 316738 -1368
rect 316806 -1424 316862 -1368
rect 316434 -1548 316490 -1492
rect 316558 -1548 316614 -1492
rect 316682 -1548 316738 -1492
rect 316806 -1548 316862 -1492
rect 343434 40294 343490 40350
rect 343558 40294 343614 40350
rect 343682 40294 343738 40350
rect 343806 40294 343862 40350
rect 343434 40170 343490 40226
rect 343558 40170 343614 40226
rect 343682 40170 343738 40226
rect 343806 40170 343862 40226
rect 343434 40046 343490 40102
rect 343558 40046 343614 40102
rect 343682 40046 343738 40102
rect 343806 40046 343862 40102
rect 343434 39922 343490 39978
rect 343558 39922 343614 39978
rect 343682 39922 343738 39978
rect 343806 39922 343862 39978
rect 343434 22294 343490 22350
rect 343558 22294 343614 22350
rect 343682 22294 343738 22350
rect 343806 22294 343862 22350
rect 343434 22170 343490 22226
rect 343558 22170 343614 22226
rect 343682 22170 343738 22226
rect 343806 22170 343862 22226
rect 343434 22046 343490 22102
rect 343558 22046 343614 22102
rect 343682 22046 343738 22102
rect 343806 22046 343862 22102
rect 343434 21922 343490 21978
rect 343558 21922 343614 21978
rect 343682 21922 343738 21978
rect 343806 21922 343862 21978
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 349020 397142 349076 397198
rect 353500 396962 353556 397018
rect 349020 240002 349076 240058
rect 348908 237482 348964 237538
rect 347154 118294 347210 118350
rect 347278 118294 347334 118350
rect 347402 118294 347458 118350
rect 347526 118294 347582 118350
rect 347154 118170 347210 118226
rect 347278 118170 347334 118226
rect 347402 118170 347458 118226
rect 347526 118170 347582 118226
rect 347154 118046 347210 118102
rect 347278 118046 347334 118102
rect 347402 118046 347458 118102
rect 347526 118046 347582 118102
rect 347154 117922 347210 117978
rect 347278 117922 347334 117978
rect 347402 117922 347458 117978
rect 347526 117922 347582 117978
rect 347154 100294 347210 100350
rect 347278 100294 347334 100350
rect 347402 100294 347458 100350
rect 347526 100294 347582 100350
rect 347154 100170 347210 100226
rect 347278 100170 347334 100226
rect 347402 100170 347458 100226
rect 347526 100170 347582 100226
rect 347154 100046 347210 100102
rect 347278 100046 347334 100102
rect 347402 100046 347458 100102
rect 347526 100046 347582 100102
rect 347154 99922 347210 99978
rect 347278 99922 347334 99978
rect 347402 99922 347458 99978
rect 347526 99922 347582 99978
rect 347154 82294 347210 82350
rect 347278 82294 347334 82350
rect 347402 82294 347458 82350
rect 347526 82294 347582 82350
rect 347154 82170 347210 82226
rect 347278 82170 347334 82226
rect 347402 82170 347458 82226
rect 347526 82170 347582 82226
rect 347154 82046 347210 82102
rect 347278 82046 347334 82102
rect 347402 82046 347458 82102
rect 347526 82046 347582 82102
rect 347154 81922 347210 81978
rect 347278 81922 347334 81978
rect 347402 81922 347458 81978
rect 347526 81922 347582 81978
rect 347154 64294 347210 64350
rect 347278 64294 347334 64350
rect 347402 64294 347458 64350
rect 347526 64294 347582 64350
rect 347154 64170 347210 64226
rect 347278 64170 347334 64226
rect 347402 64170 347458 64226
rect 347526 64170 347582 64226
rect 347154 64046 347210 64102
rect 347278 64046 347334 64102
rect 347402 64046 347458 64102
rect 347526 64046 347582 64102
rect 347154 63922 347210 63978
rect 347278 63922 347334 63978
rect 347402 63922 347458 63978
rect 347526 63922 347582 63978
rect 347154 46294 347210 46350
rect 347278 46294 347334 46350
rect 347402 46294 347458 46350
rect 347526 46294 347582 46350
rect 347154 46170 347210 46226
rect 347278 46170 347334 46226
rect 347402 46170 347458 46226
rect 347526 46170 347582 46226
rect 347154 46046 347210 46102
rect 347278 46046 347334 46102
rect 347402 46046 347458 46102
rect 347526 46046 347582 46102
rect 347154 45922 347210 45978
rect 347278 45922 347334 45978
rect 347402 45922 347458 45978
rect 347526 45922 347582 45978
rect 350252 379682 350308 379738
rect 349468 157742 349524 157798
rect 350588 372122 350644 372178
rect 350812 196622 350868 196678
rect 351372 192662 351428 192718
rect 350812 170522 350868 170578
rect 355852 396782 355908 396838
rect 354396 394802 354452 394858
rect 354284 368702 354340 368758
rect 353500 240182 353556 240238
rect 352716 192482 352772 192538
rect 352940 150542 352996 150598
rect 355404 366542 355460 366598
rect 354396 237662 354452 237718
rect 354508 235142 354564 235198
rect 354396 214262 354452 214318
rect 355180 210842 355236 210898
rect 356524 356102 356580 356158
rect 356188 325862 356244 325918
rect 356524 296702 356580 296758
rect 355852 242702 355908 242758
rect 355852 235142 355908 235198
rect 357084 369062 357140 369118
rect 356188 153422 356244 153478
rect 356972 180962 357028 181018
rect 357308 308942 357364 308998
rect 357868 383102 357924 383158
rect 357420 147662 357476 147718
rect 357420 146942 357476 146998
rect 357868 230282 357924 230338
rect 358540 192302 358596 192358
rect 358428 173042 358484 173098
rect 358988 406862 359044 406918
rect 358764 168722 358820 168778
rect 359324 255662 359380 255718
rect 359100 230282 359156 230338
rect 359212 214082 359268 214138
rect 359212 176282 359268 176338
rect 360444 407042 360500 407098
rect 362124 395522 362180 395578
rect 361900 391922 361956 391978
rect 361676 391382 361732 391438
rect 375452 395522 375508 395578
rect 527754 580294 527810 580350
rect 527878 580294 527934 580350
rect 528002 580294 528058 580350
rect 528126 580294 528182 580350
rect 527754 580170 527810 580226
rect 527878 580170 527934 580226
rect 528002 580170 528058 580226
rect 528126 580170 528182 580226
rect 527754 580046 527810 580102
rect 527878 580046 527934 580102
rect 528002 580046 528058 580102
rect 528126 580046 528182 580102
rect 527754 579922 527810 579978
rect 527878 579922 527934 579978
rect 528002 579922 528058 579978
rect 528126 579922 528182 579978
rect 527754 562294 527810 562350
rect 527878 562294 527934 562350
rect 528002 562294 528058 562350
rect 528126 562294 528182 562350
rect 527754 562170 527810 562226
rect 527878 562170 527934 562226
rect 528002 562170 528058 562226
rect 528126 562170 528182 562226
rect 527754 562046 527810 562102
rect 527878 562046 527934 562102
rect 528002 562046 528058 562102
rect 528126 562046 528182 562102
rect 527754 561922 527810 561978
rect 527878 561922 527934 561978
rect 528002 561922 528058 561978
rect 528126 561922 528182 561978
rect 517078 550294 517134 550350
rect 517202 550294 517258 550350
rect 517078 550170 517134 550226
rect 517202 550170 517258 550226
rect 517078 550046 517134 550102
rect 517202 550046 517258 550102
rect 517078 549922 517134 549978
rect 517202 549922 517258 549978
rect 527754 544294 527810 544350
rect 527878 544294 527934 544350
rect 528002 544294 528058 544350
rect 528126 544294 528182 544350
rect 527754 544170 527810 544226
rect 527878 544170 527934 544226
rect 528002 544170 528058 544226
rect 528126 544170 528182 544226
rect 527754 544046 527810 544102
rect 527878 544046 527934 544102
rect 528002 544046 528058 544102
rect 528126 544046 528182 544102
rect 527754 543922 527810 543978
rect 527878 543922 527934 543978
rect 528002 543922 528058 543978
rect 528126 543922 528182 543978
rect 517078 532294 517134 532350
rect 517202 532294 517258 532350
rect 517078 532170 517134 532226
rect 517202 532170 517258 532226
rect 517078 532046 517134 532102
rect 517202 532046 517258 532102
rect 517078 531922 517134 531978
rect 517202 531922 517258 531978
rect 527754 526294 527810 526350
rect 527878 526294 527934 526350
rect 528002 526294 528058 526350
rect 528126 526294 528182 526350
rect 527754 526170 527810 526226
rect 527878 526170 527934 526226
rect 528002 526170 528058 526226
rect 528126 526170 528182 526226
rect 527754 526046 527810 526102
rect 527878 526046 527934 526102
rect 528002 526046 528058 526102
rect 528126 526046 528182 526102
rect 527754 525922 527810 525978
rect 527878 525922 527934 525978
rect 528002 525922 528058 525978
rect 528126 525922 528182 525978
rect 517078 514294 517134 514350
rect 517202 514294 517258 514350
rect 517078 514170 517134 514226
rect 517202 514170 517258 514226
rect 517078 514046 517134 514102
rect 517202 514046 517258 514102
rect 517078 513922 517134 513978
rect 517202 513922 517258 513978
rect 527754 508294 527810 508350
rect 527878 508294 527934 508350
rect 528002 508294 528058 508350
rect 528126 508294 528182 508350
rect 527754 508170 527810 508226
rect 527878 508170 527934 508226
rect 528002 508170 528058 508226
rect 528126 508170 528182 508226
rect 527754 508046 527810 508102
rect 527878 508046 527934 508102
rect 528002 508046 528058 508102
rect 528126 508046 528182 508102
rect 527754 507922 527810 507978
rect 527878 507922 527934 507978
rect 528002 507922 528058 507978
rect 528126 507922 528182 507978
rect 517078 496294 517134 496350
rect 517202 496294 517258 496350
rect 517078 496170 517134 496226
rect 517202 496170 517258 496226
rect 517078 496046 517134 496102
rect 517202 496046 517258 496102
rect 517078 495922 517134 495978
rect 517202 495922 517258 495978
rect 527754 490294 527810 490350
rect 527878 490294 527934 490350
rect 528002 490294 528058 490350
rect 528126 490294 528182 490350
rect 527754 490170 527810 490226
rect 527878 490170 527934 490226
rect 528002 490170 528058 490226
rect 528126 490170 528182 490226
rect 527754 490046 527810 490102
rect 527878 490046 527934 490102
rect 528002 490046 528058 490102
rect 528126 490046 528182 490102
rect 527754 489922 527810 489978
rect 527878 489922 527934 489978
rect 528002 489922 528058 489978
rect 528126 489922 528182 489978
rect 517078 478294 517134 478350
rect 517202 478294 517258 478350
rect 517078 478170 517134 478226
rect 517202 478170 517258 478226
rect 517078 478046 517134 478102
rect 517202 478046 517258 478102
rect 517078 477922 517134 477978
rect 517202 477922 517258 477978
rect 527754 472294 527810 472350
rect 527878 472294 527934 472350
rect 528002 472294 528058 472350
rect 528126 472294 528182 472350
rect 527754 472170 527810 472226
rect 527878 472170 527934 472226
rect 528002 472170 528058 472226
rect 528126 472170 528182 472226
rect 527754 472046 527810 472102
rect 527878 472046 527934 472102
rect 528002 472046 528058 472102
rect 528126 472046 528182 472102
rect 527754 471922 527810 471978
rect 527878 471922 527934 471978
rect 528002 471922 528058 471978
rect 528126 471922 528182 471978
rect 517078 460294 517134 460350
rect 517202 460294 517258 460350
rect 517078 460170 517134 460226
rect 517202 460170 517258 460226
rect 517078 460046 517134 460102
rect 517202 460046 517258 460102
rect 517078 459922 517134 459978
rect 517202 459922 517258 459978
rect 527754 454294 527810 454350
rect 527878 454294 527934 454350
rect 528002 454294 528058 454350
rect 528126 454294 528182 454350
rect 527754 454170 527810 454226
rect 527878 454170 527934 454226
rect 528002 454170 528058 454226
rect 528126 454170 528182 454226
rect 527754 454046 527810 454102
rect 527878 454046 527934 454102
rect 528002 454046 528058 454102
rect 528126 454046 528182 454102
rect 527754 453922 527810 453978
rect 527878 453922 527934 453978
rect 528002 453922 528058 453978
rect 528126 453922 528182 453978
rect 517078 442294 517134 442350
rect 517202 442294 517258 442350
rect 517078 442170 517134 442226
rect 517202 442170 517258 442226
rect 517078 442046 517134 442102
rect 517202 442046 517258 442102
rect 517078 441922 517134 441978
rect 517202 441922 517258 441978
rect 527754 436294 527810 436350
rect 527878 436294 527934 436350
rect 528002 436294 528058 436350
rect 528126 436294 528182 436350
rect 527754 436170 527810 436226
rect 527878 436170 527934 436226
rect 528002 436170 528058 436226
rect 528126 436170 528182 436226
rect 527754 436046 527810 436102
rect 527878 436046 527934 436102
rect 528002 436046 528058 436102
rect 528126 436046 528182 436102
rect 527754 435922 527810 435978
rect 527878 435922 527934 435978
rect 528002 435922 528058 435978
rect 528126 435922 528182 435978
rect 517078 424294 517134 424350
rect 517202 424294 517258 424350
rect 517078 424170 517134 424226
rect 517202 424170 517258 424226
rect 517078 424046 517134 424102
rect 517202 424046 517258 424102
rect 517078 423922 517134 423978
rect 517202 423922 517258 423978
rect 527754 418294 527810 418350
rect 527878 418294 527934 418350
rect 528002 418294 528058 418350
rect 528126 418294 528182 418350
rect 527754 418170 527810 418226
rect 527878 418170 527934 418226
rect 528002 418170 528058 418226
rect 528126 418170 528182 418226
rect 527754 418046 527810 418102
rect 527878 418046 527934 418102
rect 528002 418046 528058 418102
rect 528126 418046 528182 418102
rect 527754 417922 527810 417978
rect 527878 417922 527934 417978
rect 528002 417922 528058 417978
rect 528126 417922 528182 417978
rect 514892 409562 514948 409618
rect 519148 409922 519204 409978
rect 527754 400294 527810 400350
rect 527878 400294 527934 400350
rect 528002 400294 528058 400350
rect 528126 400294 528182 400350
rect 527754 400170 527810 400226
rect 527878 400170 527934 400226
rect 528002 400170 528058 400226
rect 528126 400170 528182 400226
rect 527754 400046 527810 400102
rect 527878 400046 527934 400102
rect 528002 400046 528058 400102
rect 528126 400046 528182 400102
rect 527754 399922 527810 399978
rect 527878 399922 527934 399978
rect 528002 399922 528058 399978
rect 528126 399922 528182 399978
rect 526428 397142 526484 397198
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 531474 568294 531530 568350
rect 531598 568294 531654 568350
rect 531722 568294 531778 568350
rect 531846 568294 531902 568350
rect 531474 568170 531530 568226
rect 531598 568170 531654 568226
rect 531722 568170 531778 568226
rect 531846 568170 531902 568226
rect 531474 568046 531530 568102
rect 531598 568046 531654 568102
rect 531722 568046 531778 568102
rect 531846 568046 531902 568102
rect 531474 567922 531530 567978
rect 531598 567922 531654 567978
rect 531722 567922 531778 567978
rect 531846 567922 531902 567978
rect 558474 597156 558530 597212
rect 558598 597156 558654 597212
rect 558722 597156 558778 597212
rect 558846 597156 558902 597212
rect 558474 597032 558530 597088
rect 558598 597032 558654 597088
rect 558722 597032 558778 597088
rect 558846 597032 558902 597088
rect 558474 596908 558530 596964
rect 558598 596908 558654 596964
rect 558722 596908 558778 596964
rect 558846 596908 558902 596964
rect 558474 596784 558530 596840
rect 558598 596784 558654 596840
rect 558722 596784 558778 596840
rect 558846 596784 558902 596840
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 558474 580294 558530 580350
rect 558598 580294 558654 580350
rect 558722 580294 558778 580350
rect 558846 580294 558902 580350
rect 558474 580170 558530 580226
rect 558598 580170 558654 580226
rect 558722 580170 558778 580226
rect 558846 580170 558902 580226
rect 558474 580046 558530 580102
rect 558598 580046 558654 580102
rect 558722 580046 558778 580102
rect 558846 580046 558902 580102
rect 558474 579922 558530 579978
rect 558598 579922 558654 579978
rect 558722 579922 558778 579978
rect 558846 579922 558902 579978
rect 532438 562294 532494 562350
rect 532562 562294 532618 562350
rect 532438 562170 532494 562226
rect 532562 562170 532618 562226
rect 532438 562046 532494 562102
rect 532562 562046 532618 562102
rect 532438 561922 532494 561978
rect 532562 561922 532618 561978
rect 531474 550294 531530 550350
rect 531598 550294 531654 550350
rect 531722 550294 531778 550350
rect 531846 550294 531902 550350
rect 531474 550170 531530 550226
rect 531598 550170 531654 550226
rect 531722 550170 531778 550226
rect 531846 550170 531902 550226
rect 531474 550046 531530 550102
rect 531598 550046 531654 550102
rect 531722 550046 531778 550102
rect 531846 550046 531902 550102
rect 531474 549922 531530 549978
rect 531598 549922 531654 549978
rect 531722 549922 531778 549978
rect 531846 549922 531902 549978
rect 547798 550294 547854 550350
rect 547922 550294 547978 550350
rect 547798 550170 547854 550226
rect 547922 550170 547978 550226
rect 547798 550046 547854 550102
rect 547922 550046 547978 550102
rect 547798 549922 547854 549978
rect 547922 549922 547978 549978
rect 532438 544294 532494 544350
rect 532562 544294 532618 544350
rect 532438 544170 532494 544226
rect 532562 544170 532618 544226
rect 532438 544046 532494 544102
rect 532562 544046 532618 544102
rect 532438 543922 532494 543978
rect 532562 543922 532618 543978
rect 531474 532294 531530 532350
rect 531598 532294 531654 532350
rect 531722 532294 531778 532350
rect 531846 532294 531902 532350
rect 531474 532170 531530 532226
rect 531598 532170 531654 532226
rect 531722 532170 531778 532226
rect 531846 532170 531902 532226
rect 531474 532046 531530 532102
rect 531598 532046 531654 532102
rect 531722 532046 531778 532102
rect 531846 532046 531902 532102
rect 531474 531922 531530 531978
rect 531598 531922 531654 531978
rect 531722 531922 531778 531978
rect 531846 531922 531902 531978
rect 547798 532294 547854 532350
rect 547922 532294 547978 532350
rect 547798 532170 547854 532226
rect 547922 532170 547978 532226
rect 547798 532046 547854 532102
rect 547922 532046 547978 532102
rect 547798 531922 547854 531978
rect 547922 531922 547978 531978
rect 532438 526294 532494 526350
rect 532562 526294 532618 526350
rect 532438 526170 532494 526226
rect 532562 526170 532618 526226
rect 532438 526046 532494 526102
rect 532562 526046 532618 526102
rect 532438 525922 532494 525978
rect 532562 525922 532618 525978
rect 531474 514294 531530 514350
rect 531598 514294 531654 514350
rect 531722 514294 531778 514350
rect 531846 514294 531902 514350
rect 531474 514170 531530 514226
rect 531598 514170 531654 514226
rect 531722 514170 531778 514226
rect 531846 514170 531902 514226
rect 531474 514046 531530 514102
rect 531598 514046 531654 514102
rect 531722 514046 531778 514102
rect 531846 514046 531902 514102
rect 531474 513922 531530 513978
rect 531598 513922 531654 513978
rect 531722 513922 531778 513978
rect 531846 513922 531902 513978
rect 547798 514294 547854 514350
rect 547922 514294 547978 514350
rect 547798 514170 547854 514226
rect 547922 514170 547978 514226
rect 547798 514046 547854 514102
rect 547922 514046 547978 514102
rect 547798 513922 547854 513978
rect 547922 513922 547978 513978
rect 532438 508294 532494 508350
rect 532562 508294 532618 508350
rect 532438 508170 532494 508226
rect 532562 508170 532618 508226
rect 532438 508046 532494 508102
rect 532562 508046 532618 508102
rect 532438 507922 532494 507978
rect 532562 507922 532618 507978
rect 531474 496294 531530 496350
rect 531598 496294 531654 496350
rect 531722 496294 531778 496350
rect 531846 496294 531902 496350
rect 531474 496170 531530 496226
rect 531598 496170 531654 496226
rect 531722 496170 531778 496226
rect 531846 496170 531902 496226
rect 531474 496046 531530 496102
rect 531598 496046 531654 496102
rect 531722 496046 531778 496102
rect 531846 496046 531902 496102
rect 531474 495922 531530 495978
rect 531598 495922 531654 495978
rect 531722 495922 531778 495978
rect 531846 495922 531902 495978
rect 547798 496294 547854 496350
rect 547922 496294 547978 496350
rect 547798 496170 547854 496226
rect 547922 496170 547978 496226
rect 547798 496046 547854 496102
rect 547922 496046 547978 496102
rect 547798 495922 547854 495978
rect 547922 495922 547978 495978
rect 532438 490294 532494 490350
rect 532562 490294 532618 490350
rect 532438 490170 532494 490226
rect 532562 490170 532618 490226
rect 532438 490046 532494 490102
rect 532562 490046 532618 490102
rect 532438 489922 532494 489978
rect 532562 489922 532618 489978
rect 531474 478294 531530 478350
rect 531598 478294 531654 478350
rect 531722 478294 531778 478350
rect 531846 478294 531902 478350
rect 531474 478170 531530 478226
rect 531598 478170 531654 478226
rect 531722 478170 531778 478226
rect 531846 478170 531902 478226
rect 531474 478046 531530 478102
rect 531598 478046 531654 478102
rect 531722 478046 531778 478102
rect 531846 478046 531902 478102
rect 531474 477922 531530 477978
rect 531598 477922 531654 477978
rect 531722 477922 531778 477978
rect 531846 477922 531902 477978
rect 547798 478294 547854 478350
rect 547922 478294 547978 478350
rect 547798 478170 547854 478226
rect 547922 478170 547978 478226
rect 547798 478046 547854 478102
rect 547922 478046 547978 478102
rect 547798 477922 547854 477978
rect 547922 477922 547978 477978
rect 532438 472294 532494 472350
rect 532562 472294 532618 472350
rect 532438 472170 532494 472226
rect 532562 472170 532618 472226
rect 532438 472046 532494 472102
rect 532562 472046 532618 472102
rect 532438 471922 532494 471978
rect 532562 471922 532618 471978
rect 531474 460294 531530 460350
rect 531598 460294 531654 460350
rect 531722 460294 531778 460350
rect 531846 460294 531902 460350
rect 531474 460170 531530 460226
rect 531598 460170 531654 460226
rect 531722 460170 531778 460226
rect 531846 460170 531902 460226
rect 531474 460046 531530 460102
rect 531598 460046 531654 460102
rect 531722 460046 531778 460102
rect 531846 460046 531902 460102
rect 531474 459922 531530 459978
rect 531598 459922 531654 459978
rect 531722 459922 531778 459978
rect 531846 459922 531902 459978
rect 547798 460294 547854 460350
rect 547922 460294 547978 460350
rect 547798 460170 547854 460226
rect 547922 460170 547978 460226
rect 547798 460046 547854 460102
rect 547922 460046 547978 460102
rect 547798 459922 547854 459978
rect 547922 459922 547978 459978
rect 532438 454294 532494 454350
rect 532562 454294 532618 454350
rect 532438 454170 532494 454226
rect 532562 454170 532618 454226
rect 532438 454046 532494 454102
rect 532562 454046 532618 454102
rect 532438 453922 532494 453978
rect 532562 453922 532618 453978
rect 531474 442294 531530 442350
rect 531598 442294 531654 442350
rect 531722 442294 531778 442350
rect 531846 442294 531902 442350
rect 531474 442170 531530 442226
rect 531598 442170 531654 442226
rect 531722 442170 531778 442226
rect 531846 442170 531902 442226
rect 531474 442046 531530 442102
rect 531598 442046 531654 442102
rect 531722 442046 531778 442102
rect 531846 442046 531902 442102
rect 531474 441922 531530 441978
rect 531598 441922 531654 441978
rect 531722 441922 531778 441978
rect 531846 441922 531902 441978
rect 547798 442294 547854 442350
rect 547922 442294 547978 442350
rect 547798 442170 547854 442226
rect 547922 442170 547978 442226
rect 547798 442046 547854 442102
rect 547922 442046 547978 442102
rect 547798 441922 547854 441978
rect 547922 441922 547978 441978
rect 532438 436294 532494 436350
rect 532562 436294 532618 436350
rect 532438 436170 532494 436226
rect 532562 436170 532618 436226
rect 532438 436046 532494 436102
rect 532562 436046 532618 436102
rect 532438 435922 532494 435978
rect 532562 435922 532618 435978
rect 531474 424294 531530 424350
rect 531598 424294 531654 424350
rect 531722 424294 531778 424350
rect 531846 424294 531902 424350
rect 531474 424170 531530 424226
rect 531598 424170 531654 424226
rect 531722 424170 531778 424226
rect 531846 424170 531902 424226
rect 531474 424046 531530 424102
rect 531598 424046 531654 424102
rect 531722 424046 531778 424102
rect 531846 424046 531902 424102
rect 531474 423922 531530 423978
rect 531598 423922 531654 423978
rect 531722 423922 531778 423978
rect 531846 423922 531902 423978
rect 547798 424294 547854 424350
rect 547922 424294 547978 424350
rect 547798 424170 547854 424226
rect 547922 424170 547978 424226
rect 547798 424046 547854 424102
rect 547922 424046 547978 424102
rect 547798 423922 547854 423978
rect 547922 423922 547978 423978
rect 532438 418294 532494 418350
rect 532562 418294 532618 418350
rect 532438 418170 532494 418226
rect 532562 418170 532618 418226
rect 532438 418046 532494 418102
rect 532562 418046 532618 418102
rect 532438 417922 532494 417978
rect 532562 417922 532618 417978
rect 533820 407042 533876 407098
rect 539196 406862 539252 406918
rect 531474 406294 531530 406350
rect 531598 406294 531654 406350
rect 531722 406294 531778 406350
rect 531846 406294 531902 406350
rect 531474 406170 531530 406226
rect 531598 406170 531654 406226
rect 531722 406170 531778 406226
rect 531846 406170 531902 406226
rect 531474 406046 531530 406102
rect 531598 406046 531654 406102
rect 531722 406046 531778 406102
rect 531846 406046 531902 406102
rect 531474 405922 531530 405978
rect 531598 405922 531654 405978
rect 531722 405922 531778 405978
rect 531846 405922 531902 405978
rect 549388 400562 549444 400618
rect 551180 407402 551236 407458
rect 558474 562294 558530 562350
rect 558598 562294 558654 562350
rect 558722 562294 558778 562350
rect 558846 562294 558902 562350
rect 558474 562170 558530 562226
rect 558598 562170 558654 562226
rect 558722 562170 558778 562226
rect 558846 562170 558902 562226
rect 558474 562046 558530 562102
rect 558598 562046 558654 562102
rect 558722 562046 558778 562102
rect 558846 562046 558902 562102
rect 558474 561922 558530 561978
rect 558598 561922 558654 561978
rect 558722 561922 558778 561978
rect 558846 561922 558902 561978
rect 556108 410822 556164 410878
rect 558474 544294 558530 544350
rect 558598 544294 558654 544350
rect 558722 544294 558778 544350
rect 558846 544294 558902 544350
rect 558474 544170 558530 544226
rect 558598 544170 558654 544226
rect 558722 544170 558778 544226
rect 558846 544170 558902 544226
rect 558474 544046 558530 544102
rect 558598 544046 558654 544102
rect 558722 544046 558778 544102
rect 558846 544046 558902 544102
rect 558474 543922 558530 543978
rect 558598 543922 558654 543978
rect 558722 543922 558778 543978
rect 558846 543922 558902 543978
rect 556220 409202 556276 409258
rect 552748 405602 552804 405658
rect 556444 410642 556500 410698
rect 558474 526294 558530 526350
rect 558598 526294 558654 526350
rect 558722 526294 558778 526350
rect 558846 526294 558902 526350
rect 558474 526170 558530 526226
rect 558598 526170 558654 526226
rect 558722 526170 558778 526226
rect 558846 526170 558902 526226
rect 558474 526046 558530 526102
rect 558598 526046 558654 526102
rect 558722 526046 558778 526102
rect 558846 526046 558902 526102
rect 558474 525922 558530 525978
rect 558598 525922 558654 525978
rect 558722 525922 558778 525978
rect 558846 525922 558902 525978
rect 558474 508294 558530 508350
rect 558598 508294 558654 508350
rect 558722 508294 558778 508350
rect 558846 508294 558902 508350
rect 558474 508170 558530 508226
rect 558598 508170 558654 508226
rect 558722 508170 558778 508226
rect 558846 508170 558902 508226
rect 558474 508046 558530 508102
rect 558598 508046 558654 508102
rect 558722 508046 558778 508102
rect 558846 508046 558902 508102
rect 558474 507922 558530 507978
rect 558598 507922 558654 507978
rect 558722 507922 558778 507978
rect 558846 507922 558902 507978
rect 558474 490294 558530 490350
rect 558598 490294 558654 490350
rect 558722 490294 558778 490350
rect 558846 490294 558902 490350
rect 558474 490170 558530 490226
rect 558598 490170 558654 490226
rect 558722 490170 558778 490226
rect 558846 490170 558902 490226
rect 558474 490046 558530 490102
rect 558598 490046 558654 490102
rect 558722 490046 558778 490102
rect 558846 490046 558902 490102
rect 558474 489922 558530 489978
rect 558598 489922 558654 489978
rect 558722 489922 558778 489978
rect 558846 489922 558902 489978
rect 558474 472294 558530 472350
rect 558598 472294 558654 472350
rect 558722 472294 558778 472350
rect 558846 472294 558902 472350
rect 558474 472170 558530 472226
rect 558598 472170 558654 472226
rect 558722 472170 558778 472226
rect 558846 472170 558902 472226
rect 558474 472046 558530 472102
rect 558598 472046 558654 472102
rect 558722 472046 558778 472102
rect 558846 472046 558902 472102
rect 558474 471922 558530 471978
rect 558598 471922 558654 471978
rect 558722 471922 558778 471978
rect 558846 471922 558902 471978
rect 558474 454294 558530 454350
rect 558598 454294 558654 454350
rect 558722 454294 558778 454350
rect 558846 454294 558902 454350
rect 558474 454170 558530 454226
rect 558598 454170 558654 454226
rect 558722 454170 558778 454226
rect 558846 454170 558902 454226
rect 558474 454046 558530 454102
rect 558598 454046 558654 454102
rect 558722 454046 558778 454102
rect 558846 454046 558902 454102
rect 558474 453922 558530 453978
rect 558598 453922 558654 453978
rect 558722 453922 558778 453978
rect 558846 453922 558902 453978
rect 558474 436294 558530 436350
rect 558598 436294 558654 436350
rect 558722 436294 558778 436350
rect 558846 436294 558902 436350
rect 558474 436170 558530 436226
rect 558598 436170 558654 436226
rect 558722 436170 558778 436226
rect 558846 436170 558902 436226
rect 558474 436046 558530 436102
rect 558598 436046 558654 436102
rect 558722 436046 558778 436102
rect 558846 436046 558902 436102
rect 558474 435922 558530 435978
rect 558598 435922 558654 435978
rect 558722 435922 558778 435978
rect 558846 435922 558902 435978
rect 558474 418294 558530 418350
rect 558598 418294 558654 418350
rect 558722 418294 558778 418350
rect 558846 418294 558902 418350
rect 558474 418170 558530 418226
rect 558598 418170 558654 418226
rect 558722 418170 558778 418226
rect 558846 418170 558902 418226
rect 558474 418046 558530 418102
rect 558598 418046 558654 418102
rect 558722 418046 558778 418102
rect 558846 418046 558902 418102
rect 558474 417922 558530 417978
rect 558598 417922 558654 417978
rect 558722 417922 558778 417978
rect 558846 417922 558902 417978
rect 557788 406682 557844 406738
rect 556332 399302 556388 399358
rect 560252 404522 560308 404578
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 562194 568294 562250 568350
rect 562318 568294 562374 568350
rect 562442 568294 562498 568350
rect 562566 568294 562622 568350
rect 562194 568170 562250 568226
rect 562318 568170 562374 568226
rect 562442 568170 562498 568226
rect 562566 568170 562622 568226
rect 562194 568046 562250 568102
rect 562318 568046 562374 568102
rect 562442 568046 562498 568102
rect 562566 568046 562622 568102
rect 562194 567922 562250 567978
rect 562318 567922 562374 567978
rect 562442 567922 562498 567978
rect 562566 567922 562622 567978
rect 562194 550294 562250 550350
rect 562318 550294 562374 550350
rect 562442 550294 562498 550350
rect 562566 550294 562622 550350
rect 562194 550170 562250 550226
rect 562318 550170 562374 550226
rect 562442 550170 562498 550226
rect 562566 550170 562622 550226
rect 562194 550046 562250 550102
rect 562318 550046 562374 550102
rect 562442 550046 562498 550102
rect 562566 550046 562622 550102
rect 562194 549922 562250 549978
rect 562318 549922 562374 549978
rect 562442 549922 562498 549978
rect 562566 549922 562622 549978
rect 562194 532294 562250 532350
rect 562318 532294 562374 532350
rect 562442 532294 562498 532350
rect 562566 532294 562622 532350
rect 562194 532170 562250 532226
rect 562318 532170 562374 532226
rect 562442 532170 562498 532226
rect 562566 532170 562622 532226
rect 562194 532046 562250 532102
rect 562318 532046 562374 532102
rect 562442 532046 562498 532102
rect 562566 532046 562622 532102
rect 562194 531922 562250 531978
rect 562318 531922 562374 531978
rect 562442 531922 562498 531978
rect 562566 531922 562622 531978
rect 562194 514294 562250 514350
rect 562318 514294 562374 514350
rect 562442 514294 562498 514350
rect 562566 514294 562622 514350
rect 562194 514170 562250 514226
rect 562318 514170 562374 514226
rect 562442 514170 562498 514226
rect 562566 514170 562622 514226
rect 562194 514046 562250 514102
rect 562318 514046 562374 514102
rect 562442 514046 562498 514102
rect 562566 514046 562622 514102
rect 562194 513922 562250 513978
rect 562318 513922 562374 513978
rect 562442 513922 562498 513978
rect 562566 513922 562622 513978
rect 562194 496294 562250 496350
rect 562318 496294 562374 496350
rect 562442 496294 562498 496350
rect 562566 496294 562622 496350
rect 562194 496170 562250 496226
rect 562318 496170 562374 496226
rect 562442 496170 562498 496226
rect 562566 496170 562622 496226
rect 562194 496046 562250 496102
rect 562318 496046 562374 496102
rect 562442 496046 562498 496102
rect 562566 496046 562622 496102
rect 562194 495922 562250 495978
rect 562318 495922 562374 495978
rect 562442 495922 562498 495978
rect 562566 495922 562622 495978
rect 562194 478294 562250 478350
rect 562318 478294 562374 478350
rect 562442 478294 562498 478350
rect 562566 478294 562622 478350
rect 562194 478170 562250 478226
rect 562318 478170 562374 478226
rect 562442 478170 562498 478226
rect 562566 478170 562622 478226
rect 562194 478046 562250 478102
rect 562318 478046 562374 478102
rect 562442 478046 562498 478102
rect 562566 478046 562622 478102
rect 562194 477922 562250 477978
rect 562318 477922 562374 477978
rect 562442 477922 562498 477978
rect 562566 477922 562622 477978
rect 562194 460294 562250 460350
rect 562318 460294 562374 460350
rect 562442 460294 562498 460350
rect 562566 460294 562622 460350
rect 562194 460170 562250 460226
rect 562318 460170 562374 460226
rect 562442 460170 562498 460226
rect 562566 460170 562622 460226
rect 562194 460046 562250 460102
rect 562318 460046 562374 460102
rect 562442 460046 562498 460102
rect 562566 460046 562622 460102
rect 562194 459922 562250 459978
rect 562318 459922 562374 459978
rect 562442 459922 562498 459978
rect 562566 459922 562622 459978
rect 562194 442294 562250 442350
rect 562318 442294 562374 442350
rect 562442 442294 562498 442350
rect 562566 442294 562622 442350
rect 562194 442170 562250 442226
rect 562318 442170 562374 442226
rect 562442 442170 562498 442226
rect 562566 442170 562622 442226
rect 562194 442046 562250 442102
rect 562318 442046 562374 442102
rect 562442 442046 562498 442102
rect 562566 442046 562622 442102
rect 562194 441922 562250 441978
rect 562318 441922 562374 441978
rect 562442 441922 562498 441978
rect 562566 441922 562622 441978
rect 562194 424294 562250 424350
rect 562318 424294 562374 424350
rect 562442 424294 562498 424350
rect 562566 424294 562622 424350
rect 562194 424170 562250 424226
rect 562318 424170 562374 424226
rect 562442 424170 562498 424226
rect 562566 424170 562622 424226
rect 562194 424046 562250 424102
rect 562318 424046 562374 424102
rect 562442 424046 562498 424102
rect 562566 424046 562622 424102
rect 562194 423922 562250 423978
rect 562318 423922 562374 423978
rect 562442 423922 562498 423978
rect 562566 423922 562622 423978
rect 562194 406294 562250 406350
rect 562318 406294 562374 406350
rect 562442 406294 562498 406350
rect 562566 406294 562622 406350
rect 562194 406170 562250 406226
rect 562318 406170 562374 406226
rect 562442 406170 562498 406226
rect 562566 406170 562622 406226
rect 562194 406046 562250 406102
rect 562318 406046 562374 406102
rect 562442 406046 562498 406102
rect 562566 406046 562622 406102
rect 562194 405922 562250 405978
rect 562318 405922 562374 405978
rect 562442 405922 562498 405978
rect 562566 405922 562622 405978
rect 558474 400294 558530 400350
rect 558598 400294 558654 400350
rect 558722 400294 558778 400350
rect 558846 400294 558902 400350
rect 558474 400170 558530 400226
rect 558598 400170 558654 400226
rect 558722 400170 558778 400226
rect 558846 400170 558902 400226
rect 558474 400046 558530 400102
rect 558598 400046 558654 400102
rect 558722 400046 558778 400102
rect 558846 400046 558902 400102
rect 558474 399922 558530 399978
rect 558598 399922 558654 399978
rect 558722 399922 558778 399978
rect 558846 399922 558902 399978
rect 551068 399122 551124 399178
rect 549500 398942 549556 398998
rect 532476 396962 532532 397018
rect 556668 396782 556724 396838
rect 550620 396602 550676 396658
rect 538524 394828 538580 394858
rect 538524 394802 538580 394828
rect 559468 398222 559524 398278
rect 441756 392282 441812 392338
rect 362124 391742 362180 391798
rect 379878 388294 379934 388350
rect 380002 388294 380058 388350
rect 379878 388170 379934 388226
rect 380002 388170 380058 388226
rect 379878 388046 379934 388102
rect 380002 388046 380058 388102
rect 379878 387922 379934 387978
rect 380002 387922 380058 387978
rect 410598 388294 410654 388350
rect 410722 388294 410778 388350
rect 410598 388170 410654 388226
rect 410722 388170 410778 388226
rect 410598 388046 410654 388102
rect 410722 388046 410778 388102
rect 410598 387922 410654 387978
rect 410722 387922 410778 387978
rect 441318 388294 441374 388350
rect 441442 388294 441498 388350
rect 441318 388170 441374 388226
rect 441442 388170 441498 388226
rect 441318 388046 441374 388102
rect 441442 388046 441498 388102
rect 441318 387922 441374 387978
rect 441442 387922 441498 387978
rect 472038 388294 472094 388350
rect 472162 388294 472218 388350
rect 472038 388170 472094 388226
rect 472162 388170 472218 388226
rect 472038 388046 472094 388102
rect 472162 388046 472218 388102
rect 472038 387922 472094 387978
rect 472162 387922 472218 387978
rect 502758 388294 502814 388350
rect 502882 388294 502938 388350
rect 502758 388170 502814 388226
rect 502882 388170 502938 388226
rect 502758 388046 502814 388102
rect 502882 388046 502938 388102
rect 502758 387922 502814 387978
rect 502882 387922 502938 387978
rect 533478 388294 533534 388350
rect 533602 388294 533658 388350
rect 533478 388170 533534 388226
rect 533602 388170 533658 388226
rect 533478 388046 533534 388102
rect 533602 388046 533658 388102
rect 533478 387922 533534 387978
rect 533602 387922 533658 387978
rect 362124 383102 362180 383158
rect 364518 382294 364574 382350
rect 364642 382294 364698 382350
rect 364518 382170 364574 382226
rect 364642 382170 364698 382226
rect 364518 382046 364574 382102
rect 364642 382046 364698 382102
rect 364518 381922 364574 381978
rect 364642 381922 364698 381978
rect 395238 382294 395294 382350
rect 395362 382294 395418 382350
rect 395238 382170 395294 382226
rect 395362 382170 395418 382226
rect 395238 382046 395294 382102
rect 395362 382046 395418 382102
rect 395238 381922 395294 381978
rect 395362 381922 395418 381978
rect 425958 382294 426014 382350
rect 426082 382294 426138 382350
rect 425958 382170 426014 382226
rect 426082 382170 426138 382226
rect 425958 382046 426014 382102
rect 426082 382046 426138 382102
rect 425958 381922 426014 381978
rect 426082 381922 426138 381978
rect 456678 382294 456734 382350
rect 456802 382294 456858 382350
rect 456678 382170 456734 382226
rect 456802 382170 456858 382226
rect 456678 382046 456734 382102
rect 456802 382046 456858 382102
rect 456678 381922 456734 381978
rect 456802 381922 456858 381978
rect 487398 382294 487454 382350
rect 487522 382294 487578 382350
rect 487398 382170 487454 382226
rect 487522 382170 487578 382226
rect 487398 382046 487454 382102
rect 487522 382046 487578 382102
rect 487398 381922 487454 381978
rect 487522 381922 487578 381978
rect 518118 382294 518174 382350
rect 518242 382294 518298 382350
rect 518118 382170 518174 382226
rect 518242 382170 518298 382226
rect 518118 382046 518174 382102
rect 518242 382046 518298 382102
rect 518118 381922 518174 381978
rect 518242 381922 518298 381978
rect 548838 382294 548894 382350
rect 548962 382294 549018 382350
rect 548838 382170 548894 382226
rect 548962 382170 549018 382226
rect 548838 382046 548894 382102
rect 548962 382046 549018 382102
rect 548838 381922 548894 381978
rect 548962 381922 549018 381978
rect 379878 370294 379934 370350
rect 380002 370294 380058 370350
rect 379878 370170 379934 370226
rect 380002 370170 380058 370226
rect 379878 370046 379934 370102
rect 380002 370046 380058 370102
rect 379878 369922 379934 369978
rect 380002 369922 380058 369978
rect 410598 370294 410654 370350
rect 410722 370294 410778 370350
rect 410598 370170 410654 370226
rect 410722 370170 410778 370226
rect 410598 370046 410654 370102
rect 410722 370046 410778 370102
rect 410598 369922 410654 369978
rect 410722 369922 410778 369978
rect 441318 370294 441374 370350
rect 441442 370294 441498 370350
rect 441318 370170 441374 370226
rect 441442 370170 441498 370226
rect 441318 370046 441374 370102
rect 441442 370046 441498 370102
rect 441318 369922 441374 369978
rect 441442 369922 441498 369978
rect 472038 370294 472094 370350
rect 472162 370294 472218 370350
rect 472038 370170 472094 370226
rect 472162 370170 472218 370226
rect 472038 370046 472094 370102
rect 472162 370046 472218 370102
rect 472038 369922 472094 369978
rect 472162 369922 472218 369978
rect 502758 370294 502814 370350
rect 502882 370294 502938 370350
rect 502758 370170 502814 370226
rect 502882 370170 502938 370226
rect 502758 370046 502814 370102
rect 502882 370046 502938 370102
rect 502758 369922 502814 369978
rect 502882 369922 502938 369978
rect 533478 370294 533534 370350
rect 533602 370294 533658 370350
rect 533478 370170 533534 370226
rect 533602 370170 533658 370226
rect 533478 370046 533534 370102
rect 533602 370046 533658 370102
rect 533478 369922 533534 369978
rect 533602 369922 533658 369978
rect 364518 364294 364574 364350
rect 364642 364294 364698 364350
rect 364518 364170 364574 364226
rect 364642 364170 364698 364226
rect 364518 364046 364574 364102
rect 364642 364046 364698 364102
rect 364518 363922 364574 363978
rect 364642 363922 364698 363978
rect 395238 364294 395294 364350
rect 395362 364294 395418 364350
rect 395238 364170 395294 364226
rect 395362 364170 395418 364226
rect 395238 364046 395294 364102
rect 395362 364046 395418 364102
rect 395238 363922 395294 363978
rect 395362 363922 395418 363978
rect 425958 364294 426014 364350
rect 426082 364294 426138 364350
rect 425958 364170 426014 364226
rect 426082 364170 426138 364226
rect 425958 364046 426014 364102
rect 426082 364046 426138 364102
rect 425958 363922 426014 363978
rect 426082 363922 426138 363978
rect 456678 364294 456734 364350
rect 456802 364294 456858 364350
rect 456678 364170 456734 364226
rect 456802 364170 456858 364226
rect 456678 364046 456734 364102
rect 456802 364046 456858 364102
rect 456678 363922 456734 363978
rect 456802 363922 456858 363978
rect 487398 364294 487454 364350
rect 487522 364294 487578 364350
rect 487398 364170 487454 364226
rect 487522 364170 487578 364226
rect 487398 364046 487454 364102
rect 487522 364046 487578 364102
rect 487398 363922 487454 363978
rect 487522 363922 487578 363978
rect 518118 364294 518174 364350
rect 518242 364294 518298 364350
rect 518118 364170 518174 364226
rect 518242 364170 518298 364226
rect 518118 364046 518174 364102
rect 518242 364046 518298 364102
rect 518118 363922 518174 363978
rect 518242 363922 518298 363978
rect 548838 364294 548894 364350
rect 548962 364294 549018 364350
rect 548838 364170 548894 364226
rect 548962 364170 549018 364226
rect 548838 364046 548894 364102
rect 548962 364046 549018 364102
rect 548838 363922 548894 363978
rect 548962 363922 549018 363978
rect 379878 352294 379934 352350
rect 380002 352294 380058 352350
rect 379878 352170 379934 352226
rect 380002 352170 380058 352226
rect 379878 352046 379934 352102
rect 380002 352046 380058 352102
rect 379878 351922 379934 351978
rect 380002 351922 380058 351978
rect 410598 352294 410654 352350
rect 410722 352294 410778 352350
rect 410598 352170 410654 352226
rect 410722 352170 410778 352226
rect 410598 352046 410654 352102
rect 410722 352046 410778 352102
rect 410598 351922 410654 351978
rect 410722 351922 410778 351978
rect 441318 352294 441374 352350
rect 441442 352294 441498 352350
rect 441318 352170 441374 352226
rect 441442 352170 441498 352226
rect 441318 352046 441374 352102
rect 441442 352046 441498 352102
rect 441318 351922 441374 351978
rect 441442 351922 441498 351978
rect 472038 352294 472094 352350
rect 472162 352294 472218 352350
rect 472038 352170 472094 352226
rect 472162 352170 472218 352226
rect 472038 352046 472094 352102
rect 472162 352046 472218 352102
rect 472038 351922 472094 351978
rect 472162 351922 472218 351978
rect 502758 352294 502814 352350
rect 502882 352294 502938 352350
rect 502758 352170 502814 352226
rect 502882 352170 502938 352226
rect 502758 352046 502814 352102
rect 502882 352046 502938 352102
rect 502758 351922 502814 351978
rect 502882 351922 502938 351978
rect 533478 352294 533534 352350
rect 533602 352294 533658 352350
rect 533478 352170 533534 352226
rect 533602 352170 533658 352226
rect 533478 352046 533534 352102
rect 533602 352046 533658 352102
rect 533478 351922 533534 351978
rect 533602 351922 533658 351978
rect 364518 346294 364574 346350
rect 364642 346294 364698 346350
rect 364518 346170 364574 346226
rect 364642 346170 364698 346226
rect 364518 346046 364574 346102
rect 364642 346046 364698 346102
rect 364518 345922 364574 345978
rect 364642 345922 364698 345978
rect 395238 346294 395294 346350
rect 395362 346294 395418 346350
rect 395238 346170 395294 346226
rect 395362 346170 395418 346226
rect 395238 346046 395294 346102
rect 395362 346046 395418 346102
rect 395238 345922 395294 345978
rect 395362 345922 395418 345978
rect 425958 346294 426014 346350
rect 426082 346294 426138 346350
rect 425958 346170 426014 346226
rect 426082 346170 426138 346226
rect 425958 346046 426014 346102
rect 426082 346046 426138 346102
rect 425958 345922 426014 345978
rect 426082 345922 426138 345978
rect 456678 346294 456734 346350
rect 456802 346294 456858 346350
rect 456678 346170 456734 346226
rect 456802 346170 456858 346226
rect 456678 346046 456734 346102
rect 456802 346046 456858 346102
rect 456678 345922 456734 345978
rect 456802 345922 456858 345978
rect 487398 346294 487454 346350
rect 487522 346294 487578 346350
rect 487398 346170 487454 346226
rect 487522 346170 487578 346226
rect 487398 346046 487454 346102
rect 487522 346046 487578 346102
rect 487398 345922 487454 345978
rect 487522 345922 487578 345978
rect 518118 346294 518174 346350
rect 518242 346294 518298 346350
rect 518118 346170 518174 346226
rect 518242 346170 518298 346226
rect 518118 346046 518174 346102
rect 518242 346046 518298 346102
rect 518118 345922 518174 345978
rect 518242 345922 518298 345978
rect 548838 346294 548894 346350
rect 548962 346294 549018 346350
rect 548838 346170 548894 346226
rect 548962 346170 549018 346226
rect 548838 346046 548894 346102
rect 548962 346046 549018 346102
rect 548838 345922 548894 345978
rect 548962 345922 549018 345978
rect 379878 334294 379934 334350
rect 380002 334294 380058 334350
rect 379878 334170 379934 334226
rect 380002 334170 380058 334226
rect 379878 334046 379934 334102
rect 380002 334046 380058 334102
rect 379878 333922 379934 333978
rect 380002 333922 380058 333978
rect 410598 334294 410654 334350
rect 410722 334294 410778 334350
rect 410598 334170 410654 334226
rect 410722 334170 410778 334226
rect 410598 334046 410654 334102
rect 410722 334046 410778 334102
rect 410598 333922 410654 333978
rect 410722 333922 410778 333978
rect 441318 334294 441374 334350
rect 441442 334294 441498 334350
rect 441318 334170 441374 334226
rect 441442 334170 441498 334226
rect 441318 334046 441374 334102
rect 441442 334046 441498 334102
rect 441318 333922 441374 333978
rect 441442 333922 441498 333978
rect 472038 334294 472094 334350
rect 472162 334294 472218 334350
rect 472038 334170 472094 334226
rect 472162 334170 472218 334226
rect 472038 334046 472094 334102
rect 472162 334046 472218 334102
rect 472038 333922 472094 333978
rect 472162 333922 472218 333978
rect 502758 334294 502814 334350
rect 502882 334294 502938 334350
rect 502758 334170 502814 334226
rect 502882 334170 502938 334226
rect 502758 334046 502814 334102
rect 502882 334046 502938 334102
rect 502758 333922 502814 333978
rect 502882 333922 502938 333978
rect 533478 334294 533534 334350
rect 533602 334294 533658 334350
rect 533478 334170 533534 334226
rect 533602 334170 533658 334226
rect 533478 334046 533534 334102
rect 533602 334046 533658 334102
rect 533478 333922 533534 333978
rect 533602 333922 533658 333978
rect 364518 328294 364574 328350
rect 364642 328294 364698 328350
rect 364518 328170 364574 328226
rect 364642 328170 364698 328226
rect 364518 328046 364574 328102
rect 364642 328046 364698 328102
rect 364518 327922 364574 327978
rect 364642 327922 364698 327978
rect 395238 328294 395294 328350
rect 395362 328294 395418 328350
rect 395238 328170 395294 328226
rect 395362 328170 395418 328226
rect 395238 328046 395294 328102
rect 395362 328046 395418 328102
rect 395238 327922 395294 327978
rect 395362 327922 395418 327978
rect 425958 328294 426014 328350
rect 426082 328294 426138 328350
rect 425958 328170 426014 328226
rect 426082 328170 426138 328226
rect 425958 328046 426014 328102
rect 426082 328046 426138 328102
rect 425958 327922 426014 327978
rect 426082 327922 426138 327978
rect 456678 328294 456734 328350
rect 456802 328294 456858 328350
rect 456678 328170 456734 328226
rect 456802 328170 456858 328226
rect 456678 328046 456734 328102
rect 456802 328046 456858 328102
rect 456678 327922 456734 327978
rect 456802 327922 456858 327978
rect 487398 328294 487454 328350
rect 487522 328294 487578 328350
rect 487398 328170 487454 328226
rect 487522 328170 487578 328226
rect 487398 328046 487454 328102
rect 487522 328046 487578 328102
rect 487398 327922 487454 327978
rect 487522 327922 487578 327978
rect 518118 328294 518174 328350
rect 518242 328294 518298 328350
rect 518118 328170 518174 328226
rect 518242 328170 518298 328226
rect 518118 328046 518174 328102
rect 518242 328046 518298 328102
rect 518118 327922 518174 327978
rect 518242 327922 518298 327978
rect 548838 328294 548894 328350
rect 548962 328294 549018 328350
rect 548838 328170 548894 328226
rect 548962 328170 549018 328226
rect 548838 328046 548894 328102
rect 548962 328046 549018 328102
rect 548838 327922 548894 327978
rect 548962 327922 549018 327978
rect 379878 316294 379934 316350
rect 380002 316294 380058 316350
rect 379878 316170 379934 316226
rect 380002 316170 380058 316226
rect 379878 316046 379934 316102
rect 380002 316046 380058 316102
rect 379878 315922 379934 315978
rect 380002 315922 380058 315978
rect 410598 316294 410654 316350
rect 410722 316294 410778 316350
rect 410598 316170 410654 316226
rect 410722 316170 410778 316226
rect 410598 316046 410654 316102
rect 410722 316046 410778 316102
rect 410598 315922 410654 315978
rect 410722 315922 410778 315978
rect 441318 316294 441374 316350
rect 441442 316294 441498 316350
rect 441318 316170 441374 316226
rect 441442 316170 441498 316226
rect 441318 316046 441374 316102
rect 441442 316046 441498 316102
rect 441318 315922 441374 315978
rect 441442 315922 441498 315978
rect 472038 316294 472094 316350
rect 472162 316294 472218 316350
rect 472038 316170 472094 316226
rect 472162 316170 472218 316226
rect 472038 316046 472094 316102
rect 472162 316046 472218 316102
rect 472038 315922 472094 315978
rect 472162 315922 472218 315978
rect 502758 316294 502814 316350
rect 502882 316294 502938 316350
rect 502758 316170 502814 316226
rect 502882 316170 502938 316226
rect 502758 316046 502814 316102
rect 502882 316046 502938 316102
rect 502758 315922 502814 315978
rect 502882 315922 502938 315978
rect 533478 316294 533534 316350
rect 533602 316294 533658 316350
rect 533478 316170 533534 316226
rect 533602 316170 533658 316226
rect 533478 316046 533534 316102
rect 533602 316046 533658 316102
rect 533478 315922 533534 315978
rect 533602 315922 533658 315978
rect 364518 310294 364574 310350
rect 364642 310294 364698 310350
rect 364518 310170 364574 310226
rect 364642 310170 364698 310226
rect 364518 310046 364574 310102
rect 364642 310046 364698 310102
rect 364518 309922 364574 309978
rect 364642 309922 364698 309978
rect 395238 310294 395294 310350
rect 395362 310294 395418 310350
rect 395238 310170 395294 310226
rect 395362 310170 395418 310226
rect 395238 310046 395294 310102
rect 395362 310046 395418 310102
rect 395238 309922 395294 309978
rect 395362 309922 395418 309978
rect 425958 310294 426014 310350
rect 426082 310294 426138 310350
rect 425958 310170 426014 310226
rect 426082 310170 426138 310226
rect 425958 310046 426014 310102
rect 426082 310046 426138 310102
rect 425958 309922 426014 309978
rect 426082 309922 426138 309978
rect 456678 310294 456734 310350
rect 456802 310294 456858 310350
rect 456678 310170 456734 310226
rect 456802 310170 456858 310226
rect 456678 310046 456734 310102
rect 456802 310046 456858 310102
rect 456678 309922 456734 309978
rect 456802 309922 456858 309978
rect 487398 310294 487454 310350
rect 487522 310294 487578 310350
rect 487398 310170 487454 310226
rect 487522 310170 487578 310226
rect 487398 310046 487454 310102
rect 487522 310046 487578 310102
rect 487398 309922 487454 309978
rect 487522 309922 487578 309978
rect 518118 310294 518174 310350
rect 518242 310294 518298 310350
rect 518118 310170 518174 310226
rect 518242 310170 518298 310226
rect 518118 310046 518174 310102
rect 518242 310046 518298 310102
rect 518118 309922 518174 309978
rect 518242 309922 518298 309978
rect 548838 310294 548894 310350
rect 548962 310294 549018 310350
rect 548838 310170 548894 310226
rect 548962 310170 549018 310226
rect 548838 310046 548894 310102
rect 548962 310046 549018 310102
rect 548838 309922 548894 309978
rect 548962 309922 549018 309978
rect 359884 308582 359940 308638
rect 360108 308582 360164 308638
rect 360108 308402 360164 308458
rect 360332 308222 360388 308278
rect 359660 235900 359716 235918
rect 359660 235862 359716 235900
rect 359996 287342 360052 287398
rect 359996 235862 360052 235918
rect 359772 191762 359828 191818
rect 359772 186002 359828 186058
rect 359772 185642 359828 185698
rect 359996 185822 360052 185878
rect 360220 296702 360276 296758
rect 360220 185642 360276 185698
rect 379878 298294 379934 298350
rect 380002 298294 380058 298350
rect 379878 298170 379934 298226
rect 380002 298170 380058 298226
rect 379878 298046 379934 298102
rect 380002 298046 380058 298102
rect 379878 297922 379934 297978
rect 380002 297922 380058 297978
rect 410598 298294 410654 298350
rect 410722 298294 410778 298350
rect 410598 298170 410654 298226
rect 410722 298170 410778 298226
rect 410598 298046 410654 298102
rect 410722 298046 410778 298102
rect 410598 297922 410654 297978
rect 410722 297922 410778 297978
rect 441318 298294 441374 298350
rect 441442 298294 441498 298350
rect 441318 298170 441374 298226
rect 441442 298170 441498 298226
rect 441318 298046 441374 298102
rect 441442 298046 441498 298102
rect 441318 297922 441374 297978
rect 441442 297922 441498 297978
rect 472038 298294 472094 298350
rect 472162 298294 472218 298350
rect 472038 298170 472094 298226
rect 472162 298170 472218 298226
rect 472038 298046 472094 298102
rect 472162 298046 472218 298102
rect 472038 297922 472094 297978
rect 472162 297922 472218 297978
rect 502758 298294 502814 298350
rect 502882 298294 502938 298350
rect 502758 298170 502814 298226
rect 502882 298170 502938 298226
rect 502758 298046 502814 298102
rect 502882 298046 502938 298102
rect 502758 297922 502814 297978
rect 502882 297922 502938 297978
rect 533478 298294 533534 298350
rect 533602 298294 533658 298350
rect 533478 298170 533534 298226
rect 533602 298170 533658 298226
rect 533478 298046 533534 298102
rect 533602 298046 533658 298102
rect 533478 297922 533534 297978
rect 533602 297922 533658 297978
rect 362012 292562 362068 292618
rect 360444 255662 360500 255718
rect 360108 157022 360164 157078
rect 361788 235862 361844 235918
rect 360556 191762 360612 191818
rect 361228 184562 361284 184618
rect 361900 193922 361956 193978
rect 361900 184562 361956 184618
rect 361564 180962 361620 181018
rect 361452 176282 361508 176338
rect 364518 292294 364574 292350
rect 364642 292294 364698 292350
rect 364518 292170 364574 292226
rect 364642 292170 364698 292226
rect 364518 292046 364574 292102
rect 364642 292046 364698 292102
rect 364518 291922 364574 291978
rect 364642 291922 364698 291978
rect 395238 292294 395294 292350
rect 395362 292294 395418 292350
rect 395238 292170 395294 292226
rect 395362 292170 395418 292226
rect 395238 292046 395294 292102
rect 395362 292046 395418 292102
rect 395238 291922 395294 291978
rect 395362 291922 395418 291978
rect 425958 292294 426014 292350
rect 426082 292294 426138 292350
rect 425958 292170 426014 292226
rect 426082 292170 426138 292226
rect 425958 292046 426014 292102
rect 426082 292046 426138 292102
rect 425958 291922 426014 291978
rect 426082 291922 426138 291978
rect 456678 292294 456734 292350
rect 456802 292294 456858 292350
rect 456678 292170 456734 292226
rect 456802 292170 456858 292226
rect 456678 292046 456734 292102
rect 456802 292046 456858 292102
rect 456678 291922 456734 291978
rect 456802 291922 456858 291978
rect 487398 292294 487454 292350
rect 487522 292294 487578 292350
rect 487398 292170 487454 292226
rect 487522 292170 487578 292226
rect 487398 292046 487454 292102
rect 487522 292046 487578 292102
rect 487398 291922 487454 291978
rect 487522 291922 487578 291978
rect 518118 292294 518174 292350
rect 518242 292294 518298 292350
rect 518118 292170 518174 292226
rect 518242 292170 518298 292226
rect 518118 292046 518174 292102
rect 518242 292046 518298 292102
rect 518118 291922 518174 291978
rect 518242 291922 518298 291978
rect 548838 292294 548894 292350
rect 548962 292294 549018 292350
rect 548838 292170 548894 292226
rect 548962 292170 549018 292226
rect 548838 292046 548894 292102
rect 548962 292046 549018 292102
rect 548838 291922 548894 291978
rect 548962 291922 549018 291978
rect 379878 280294 379934 280350
rect 380002 280294 380058 280350
rect 379878 280170 379934 280226
rect 380002 280170 380058 280226
rect 379878 280046 379934 280102
rect 380002 280046 380058 280102
rect 379878 279922 379934 279978
rect 380002 279922 380058 279978
rect 410598 280294 410654 280350
rect 410722 280294 410778 280350
rect 410598 280170 410654 280226
rect 410722 280170 410778 280226
rect 410598 280046 410654 280102
rect 410722 280046 410778 280102
rect 410598 279922 410654 279978
rect 410722 279922 410778 279978
rect 441318 280294 441374 280350
rect 441442 280294 441498 280350
rect 441318 280170 441374 280226
rect 441442 280170 441498 280226
rect 441318 280046 441374 280102
rect 441442 280046 441498 280102
rect 441318 279922 441374 279978
rect 441442 279922 441498 279978
rect 472038 280294 472094 280350
rect 472162 280294 472218 280350
rect 472038 280170 472094 280226
rect 472162 280170 472218 280226
rect 472038 280046 472094 280102
rect 472162 280046 472218 280102
rect 472038 279922 472094 279978
rect 472162 279922 472218 279978
rect 502758 280294 502814 280350
rect 502882 280294 502938 280350
rect 502758 280170 502814 280226
rect 502882 280170 502938 280226
rect 502758 280046 502814 280102
rect 502882 280046 502938 280102
rect 502758 279922 502814 279978
rect 502882 279922 502938 279978
rect 533478 280294 533534 280350
rect 533602 280294 533658 280350
rect 533478 280170 533534 280226
rect 533602 280170 533658 280226
rect 533478 280046 533534 280102
rect 533602 280046 533658 280102
rect 533478 279922 533534 279978
rect 533602 279922 533658 279978
rect 364518 274294 364574 274350
rect 364642 274294 364698 274350
rect 364518 274170 364574 274226
rect 364642 274170 364698 274226
rect 364518 274046 364574 274102
rect 364642 274046 364698 274102
rect 364518 273922 364574 273978
rect 364642 273922 364698 273978
rect 395238 274294 395294 274350
rect 395362 274294 395418 274350
rect 395238 274170 395294 274226
rect 395362 274170 395418 274226
rect 395238 274046 395294 274102
rect 395362 274046 395418 274102
rect 395238 273922 395294 273978
rect 395362 273922 395418 273978
rect 425958 274294 426014 274350
rect 426082 274294 426138 274350
rect 425958 274170 426014 274226
rect 426082 274170 426138 274226
rect 425958 274046 426014 274102
rect 426082 274046 426138 274102
rect 425958 273922 426014 273978
rect 426082 273922 426138 273978
rect 456678 274294 456734 274350
rect 456802 274294 456858 274350
rect 456678 274170 456734 274226
rect 456802 274170 456858 274226
rect 456678 274046 456734 274102
rect 456802 274046 456858 274102
rect 456678 273922 456734 273978
rect 456802 273922 456858 273978
rect 487398 274294 487454 274350
rect 487522 274294 487578 274350
rect 487398 274170 487454 274226
rect 487522 274170 487578 274226
rect 487398 274046 487454 274102
rect 487522 274046 487578 274102
rect 487398 273922 487454 273978
rect 487522 273922 487578 273978
rect 518118 274294 518174 274350
rect 518242 274294 518298 274350
rect 518118 274170 518174 274226
rect 518242 274170 518298 274226
rect 518118 274046 518174 274102
rect 518242 274046 518298 274102
rect 518118 273922 518174 273978
rect 518242 273922 518298 273978
rect 548838 274294 548894 274350
rect 548962 274294 549018 274350
rect 548838 274170 548894 274226
rect 548962 274170 549018 274226
rect 548838 274046 548894 274102
rect 548962 274046 549018 274102
rect 548838 273922 548894 273978
rect 548962 273922 549018 273978
rect 379878 262294 379934 262350
rect 380002 262294 380058 262350
rect 379878 262170 379934 262226
rect 380002 262170 380058 262226
rect 379878 262046 379934 262102
rect 380002 262046 380058 262102
rect 379878 261922 379934 261978
rect 380002 261922 380058 261978
rect 410598 262294 410654 262350
rect 410722 262294 410778 262350
rect 410598 262170 410654 262226
rect 410722 262170 410778 262226
rect 410598 262046 410654 262102
rect 410722 262046 410778 262102
rect 410598 261922 410654 261978
rect 410722 261922 410778 261978
rect 441318 262294 441374 262350
rect 441442 262294 441498 262350
rect 441318 262170 441374 262226
rect 441442 262170 441498 262226
rect 441318 262046 441374 262102
rect 441442 262046 441498 262102
rect 441318 261922 441374 261978
rect 441442 261922 441498 261978
rect 472038 262294 472094 262350
rect 472162 262294 472218 262350
rect 472038 262170 472094 262226
rect 472162 262170 472218 262226
rect 472038 262046 472094 262102
rect 472162 262046 472218 262102
rect 472038 261922 472094 261978
rect 472162 261922 472218 261978
rect 502758 262294 502814 262350
rect 502882 262294 502938 262350
rect 502758 262170 502814 262226
rect 502882 262170 502938 262226
rect 502758 262046 502814 262102
rect 502882 262046 502938 262102
rect 502758 261922 502814 261978
rect 502882 261922 502938 261978
rect 533478 262294 533534 262350
rect 533602 262294 533658 262350
rect 533478 262170 533534 262226
rect 533602 262170 533658 262226
rect 533478 262046 533534 262102
rect 533602 262046 533658 262102
rect 533478 261922 533534 261978
rect 533602 261922 533658 261978
rect 364518 256294 364574 256350
rect 364642 256294 364698 256350
rect 364518 256170 364574 256226
rect 364642 256170 364698 256226
rect 364518 256046 364574 256102
rect 364642 256046 364698 256102
rect 364518 255922 364574 255978
rect 364642 255922 364698 255978
rect 395238 256294 395294 256350
rect 395362 256294 395418 256350
rect 395238 256170 395294 256226
rect 395362 256170 395418 256226
rect 395238 256046 395294 256102
rect 395362 256046 395418 256102
rect 395238 255922 395294 255978
rect 395362 255922 395418 255978
rect 425958 256294 426014 256350
rect 426082 256294 426138 256350
rect 425958 256170 426014 256226
rect 426082 256170 426138 256226
rect 425958 256046 426014 256102
rect 426082 256046 426138 256102
rect 425958 255922 426014 255978
rect 426082 255922 426138 255978
rect 456678 256294 456734 256350
rect 456802 256294 456858 256350
rect 456678 256170 456734 256226
rect 456802 256170 456858 256226
rect 456678 256046 456734 256102
rect 456802 256046 456858 256102
rect 456678 255922 456734 255978
rect 456802 255922 456858 255978
rect 487398 256294 487454 256350
rect 487522 256294 487578 256350
rect 487398 256170 487454 256226
rect 487522 256170 487578 256226
rect 487398 256046 487454 256102
rect 487522 256046 487578 256102
rect 487398 255922 487454 255978
rect 487522 255922 487578 255978
rect 518118 256294 518174 256350
rect 518242 256294 518298 256350
rect 518118 256170 518174 256226
rect 518242 256170 518298 256226
rect 518118 256046 518174 256102
rect 518242 256046 518298 256102
rect 518118 255922 518174 255978
rect 518242 255922 518298 255978
rect 548838 256294 548894 256350
rect 548962 256294 549018 256350
rect 548838 256170 548894 256226
rect 548962 256170 549018 256226
rect 548838 256046 548894 256102
rect 548962 256046 549018 256102
rect 548838 255922 548894 255978
rect 548962 255922 549018 255978
rect 379878 244294 379934 244350
rect 380002 244294 380058 244350
rect 379878 244170 379934 244226
rect 380002 244170 380058 244226
rect 379878 244046 379934 244102
rect 380002 244046 380058 244102
rect 379878 243922 379934 243978
rect 380002 243922 380058 243978
rect 410598 244294 410654 244350
rect 410722 244294 410778 244350
rect 410598 244170 410654 244226
rect 410722 244170 410778 244226
rect 410598 244046 410654 244102
rect 410722 244046 410778 244102
rect 410598 243922 410654 243978
rect 410722 243922 410778 243978
rect 441318 244294 441374 244350
rect 441442 244294 441498 244350
rect 441318 244170 441374 244226
rect 441442 244170 441498 244226
rect 441318 244046 441374 244102
rect 441442 244046 441498 244102
rect 441318 243922 441374 243978
rect 441442 243922 441498 243978
rect 472038 244294 472094 244350
rect 472162 244294 472218 244350
rect 472038 244170 472094 244226
rect 472162 244170 472218 244226
rect 472038 244046 472094 244102
rect 472162 244046 472218 244102
rect 472038 243922 472094 243978
rect 472162 243922 472218 243978
rect 502758 244294 502814 244350
rect 502882 244294 502938 244350
rect 502758 244170 502814 244226
rect 502882 244170 502938 244226
rect 502758 244046 502814 244102
rect 502882 244046 502938 244102
rect 502758 243922 502814 243978
rect 502882 243922 502938 243978
rect 533478 244294 533534 244350
rect 533602 244294 533658 244350
rect 533478 244170 533534 244226
rect 533602 244170 533658 244226
rect 533478 244046 533534 244102
rect 533602 244046 533658 244102
rect 533478 243922 533534 243978
rect 533602 243922 533658 243978
rect 364518 238294 364574 238350
rect 364642 238294 364698 238350
rect 364518 238170 364574 238226
rect 364642 238170 364698 238226
rect 364518 238046 364574 238102
rect 364642 238046 364698 238102
rect 364518 237922 364574 237978
rect 364642 237922 364698 237978
rect 395238 238294 395294 238350
rect 395362 238294 395418 238350
rect 395238 238170 395294 238226
rect 395362 238170 395418 238226
rect 395238 238046 395294 238102
rect 395362 238046 395418 238102
rect 395238 237922 395294 237978
rect 395362 237922 395418 237978
rect 425958 238294 426014 238350
rect 426082 238294 426138 238350
rect 425958 238170 426014 238226
rect 426082 238170 426138 238226
rect 425958 238046 426014 238102
rect 426082 238046 426138 238102
rect 425958 237922 426014 237978
rect 426082 237922 426138 237978
rect 456678 238294 456734 238350
rect 456802 238294 456858 238350
rect 456678 238170 456734 238226
rect 456802 238170 456858 238226
rect 456678 238046 456734 238102
rect 456802 238046 456858 238102
rect 456678 237922 456734 237978
rect 456802 237922 456858 237978
rect 487398 238294 487454 238350
rect 487522 238294 487578 238350
rect 487398 238170 487454 238226
rect 487522 238170 487578 238226
rect 487398 238046 487454 238102
rect 487522 238046 487578 238102
rect 487398 237922 487454 237978
rect 487522 237922 487578 237978
rect 518118 238294 518174 238350
rect 518242 238294 518298 238350
rect 518118 238170 518174 238226
rect 518242 238170 518298 238226
rect 518118 238046 518174 238102
rect 518242 238046 518298 238102
rect 518118 237922 518174 237978
rect 518242 237922 518298 237978
rect 548838 238294 548894 238350
rect 548962 238294 549018 238350
rect 548838 238170 548894 238226
rect 548962 238170 549018 238226
rect 548838 238046 548894 238102
rect 548962 238046 549018 238102
rect 548838 237922 548894 237978
rect 548962 237922 549018 237978
rect 379878 226294 379934 226350
rect 380002 226294 380058 226350
rect 379878 226170 379934 226226
rect 380002 226170 380058 226226
rect 379878 226046 379934 226102
rect 380002 226046 380058 226102
rect 379878 225922 379934 225978
rect 380002 225922 380058 225978
rect 410598 226294 410654 226350
rect 410722 226294 410778 226350
rect 410598 226170 410654 226226
rect 410722 226170 410778 226226
rect 410598 226046 410654 226102
rect 410722 226046 410778 226102
rect 410598 225922 410654 225978
rect 410722 225922 410778 225978
rect 441318 226294 441374 226350
rect 441442 226294 441498 226350
rect 441318 226170 441374 226226
rect 441442 226170 441498 226226
rect 441318 226046 441374 226102
rect 441442 226046 441498 226102
rect 441318 225922 441374 225978
rect 441442 225922 441498 225978
rect 472038 226294 472094 226350
rect 472162 226294 472218 226350
rect 472038 226170 472094 226226
rect 472162 226170 472218 226226
rect 472038 226046 472094 226102
rect 472162 226046 472218 226102
rect 472038 225922 472094 225978
rect 472162 225922 472218 225978
rect 502758 226294 502814 226350
rect 502882 226294 502938 226350
rect 502758 226170 502814 226226
rect 502882 226170 502938 226226
rect 502758 226046 502814 226102
rect 502882 226046 502938 226102
rect 502758 225922 502814 225978
rect 502882 225922 502938 225978
rect 533478 226294 533534 226350
rect 533602 226294 533658 226350
rect 533478 226170 533534 226226
rect 533602 226170 533658 226226
rect 533478 226046 533534 226102
rect 533602 226046 533658 226102
rect 533478 225922 533534 225978
rect 533602 225922 533658 225978
rect 364518 220294 364574 220350
rect 364642 220294 364698 220350
rect 364518 220170 364574 220226
rect 364642 220170 364698 220226
rect 364518 220046 364574 220102
rect 364642 220046 364698 220102
rect 364518 219922 364574 219978
rect 364642 219922 364698 219978
rect 395238 220294 395294 220350
rect 395362 220294 395418 220350
rect 395238 220170 395294 220226
rect 395362 220170 395418 220226
rect 395238 220046 395294 220102
rect 395362 220046 395418 220102
rect 395238 219922 395294 219978
rect 395362 219922 395418 219978
rect 425958 220294 426014 220350
rect 426082 220294 426138 220350
rect 425958 220170 426014 220226
rect 426082 220170 426138 220226
rect 425958 220046 426014 220102
rect 426082 220046 426138 220102
rect 425958 219922 426014 219978
rect 426082 219922 426138 219978
rect 456678 220294 456734 220350
rect 456802 220294 456858 220350
rect 456678 220170 456734 220226
rect 456802 220170 456858 220226
rect 456678 220046 456734 220102
rect 456802 220046 456858 220102
rect 456678 219922 456734 219978
rect 456802 219922 456858 219978
rect 487398 220294 487454 220350
rect 487522 220294 487578 220350
rect 487398 220170 487454 220226
rect 487522 220170 487578 220226
rect 487398 220046 487454 220102
rect 487522 220046 487578 220102
rect 487398 219922 487454 219978
rect 487522 219922 487578 219978
rect 518118 220294 518174 220350
rect 518242 220294 518298 220350
rect 518118 220170 518174 220226
rect 518242 220170 518298 220226
rect 518118 220046 518174 220102
rect 518242 220046 518298 220102
rect 518118 219922 518174 219978
rect 518242 219922 518298 219978
rect 548838 220294 548894 220350
rect 548962 220294 549018 220350
rect 548838 220170 548894 220226
rect 548962 220170 549018 220226
rect 548838 220046 548894 220102
rect 548962 220046 549018 220102
rect 548838 219922 548894 219978
rect 548962 219922 549018 219978
rect 379878 208294 379934 208350
rect 380002 208294 380058 208350
rect 379878 208170 379934 208226
rect 380002 208170 380058 208226
rect 379878 208046 379934 208102
rect 380002 208046 380058 208102
rect 379878 207922 379934 207978
rect 380002 207922 380058 207978
rect 410598 208294 410654 208350
rect 410722 208294 410778 208350
rect 410598 208170 410654 208226
rect 410722 208170 410778 208226
rect 410598 208046 410654 208102
rect 410722 208046 410778 208102
rect 410598 207922 410654 207978
rect 410722 207922 410778 207978
rect 441318 208294 441374 208350
rect 441442 208294 441498 208350
rect 441318 208170 441374 208226
rect 441442 208170 441498 208226
rect 441318 208046 441374 208102
rect 441442 208046 441498 208102
rect 441318 207922 441374 207978
rect 441442 207922 441498 207978
rect 472038 208294 472094 208350
rect 472162 208294 472218 208350
rect 472038 208170 472094 208226
rect 472162 208170 472218 208226
rect 472038 208046 472094 208102
rect 472162 208046 472218 208102
rect 472038 207922 472094 207978
rect 472162 207922 472218 207978
rect 502758 208294 502814 208350
rect 502882 208294 502938 208350
rect 502758 208170 502814 208226
rect 502882 208170 502938 208226
rect 502758 208046 502814 208102
rect 502882 208046 502938 208102
rect 502758 207922 502814 207978
rect 502882 207922 502938 207978
rect 533478 208294 533534 208350
rect 533602 208294 533658 208350
rect 533478 208170 533534 208226
rect 533602 208170 533658 208226
rect 533478 208046 533534 208102
rect 533602 208046 533658 208102
rect 533478 207922 533534 207978
rect 533602 207922 533658 207978
rect 364518 202294 364574 202350
rect 364642 202294 364698 202350
rect 364518 202170 364574 202226
rect 364642 202170 364698 202226
rect 364518 202046 364574 202102
rect 364642 202046 364698 202102
rect 364518 201922 364574 201978
rect 364642 201922 364698 201978
rect 395238 202294 395294 202350
rect 395362 202294 395418 202350
rect 395238 202170 395294 202226
rect 395362 202170 395418 202226
rect 395238 202046 395294 202102
rect 395362 202046 395418 202102
rect 395238 201922 395294 201978
rect 395362 201922 395418 201978
rect 425958 202294 426014 202350
rect 426082 202294 426138 202350
rect 425958 202170 426014 202226
rect 426082 202170 426138 202226
rect 425958 202046 426014 202102
rect 426082 202046 426138 202102
rect 425958 201922 426014 201978
rect 426082 201922 426138 201978
rect 456678 202294 456734 202350
rect 456802 202294 456858 202350
rect 456678 202170 456734 202226
rect 456802 202170 456858 202226
rect 456678 202046 456734 202102
rect 456802 202046 456858 202102
rect 456678 201922 456734 201978
rect 456802 201922 456858 201978
rect 487398 202294 487454 202350
rect 487522 202294 487578 202350
rect 487398 202170 487454 202226
rect 487522 202170 487578 202226
rect 487398 202046 487454 202102
rect 487522 202046 487578 202102
rect 487398 201922 487454 201978
rect 487522 201922 487578 201978
rect 518118 202294 518174 202350
rect 518242 202294 518298 202350
rect 518118 202170 518174 202226
rect 518242 202170 518298 202226
rect 518118 202046 518174 202102
rect 518242 202046 518298 202102
rect 518118 201922 518174 201978
rect 518242 201922 518298 201978
rect 548838 202294 548894 202350
rect 548962 202294 549018 202350
rect 548838 202170 548894 202226
rect 548962 202170 549018 202226
rect 548838 202046 548894 202102
rect 548962 202046 549018 202102
rect 548838 201922 548894 201978
rect 548962 201922 549018 201978
rect 362124 195722 362180 195778
rect 379878 190294 379934 190350
rect 380002 190294 380058 190350
rect 379878 190170 379934 190226
rect 380002 190170 380058 190226
rect 379878 190046 379934 190102
rect 380002 190046 380058 190102
rect 379878 189922 379934 189978
rect 380002 189922 380058 189978
rect 410598 190294 410654 190350
rect 410722 190294 410778 190350
rect 410598 190170 410654 190226
rect 410722 190170 410778 190226
rect 410598 190046 410654 190102
rect 410722 190046 410778 190102
rect 410598 189922 410654 189978
rect 410722 189922 410778 189978
rect 441318 190294 441374 190350
rect 441442 190294 441498 190350
rect 441318 190170 441374 190226
rect 441442 190170 441498 190226
rect 441318 190046 441374 190102
rect 441442 190046 441498 190102
rect 441318 189922 441374 189978
rect 441442 189922 441498 189978
rect 472038 190294 472094 190350
rect 472162 190294 472218 190350
rect 472038 190170 472094 190226
rect 472162 190170 472218 190226
rect 472038 190046 472094 190102
rect 472162 190046 472218 190102
rect 472038 189922 472094 189978
rect 472162 189922 472218 189978
rect 502758 190294 502814 190350
rect 502882 190294 502938 190350
rect 502758 190170 502814 190226
rect 502882 190170 502938 190226
rect 502758 190046 502814 190102
rect 502882 190046 502938 190102
rect 502758 189922 502814 189978
rect 502882 189922 502938 189978
rect 533478 190294 533534 190350
rect 533602 190294 533658 190350
rect 533478 190170 533534 190226
rect 533602 190170 533658 190226
rect 533478 190046 533534 190102
rect 533602 190046 533658 190102
rect 533478 189922 533534 189978
rect 533602 189922 533658 189978
rect 364518 184294 364574 184350
rect 364642 184294 364698 184350
rect 364518 184170 364574 184226
rect 364642 184170 364698 184226
rect 364518 184046 364574 184102
rect 364642 184046 364698 184102
rect 364518 183922 364574 183978
rect 364642 183922 364698 183978
rect 395238 184294 395294 184350
rect 395362 184294 395418 184350
rect 395238 184170 395294 184226
rect 395362 184170 395418 184226
rect 395238 184046 395294 184102
rect 395362 184046 395418 184102
rect 395238 183922 395294 183978
rect 395362 183922 395418 183978
rect 425958 184294 426014 184350
rect 426082 184294 426138 184350
rect 425958 184170 426014 184226
rect 426082 184170 426138 184226
rect 425958 184046 426014 184102
rect 426082 184046 426138 184102
rect 425958 183922 426014 183978
rect 426082 183922 426138 183978
rect 456678 184294 456734 184350
rect 456802 184294 456858 184350
rect 456678 184170 456734 184226
rect 456802 184170 456858 184226
rect 456678 184046 456734 184102
rect 456802 184046 456858 184102
rect 456678 183922 456734 183978
rect 456802 183922 456858 183978
rect 487398 184294 487454 184350
rect 487522 184294 487578 184350
rect 487398 184170 487454 184226
rect 487522 184170 487578 184226
rect 487398 184046 487454 184102
rect 487522 184046 487578 184102
rect 487398 183922 487454 183978
rect 487522 183922 487578 183978
rect 518118 184294 518174 184350
rect 518242 184294 518298 184350
rect 518118 184170 518174 184226
rect 518242 184170 518298 184226
rect 518118 184046 518174 184102
rect 518242 184046 518298 184102
rect 518118 183922 518174 183978
rect 518242 183922 518298 183978
rect 548838 184294 548894 184350
rect 548962 184294 549018 184350
rect 548838 184170 548894 184226
rect 548962 184170 549018 184226
rect 548838 184046 548894 184102
rect 548962 184046 549018 184102
rect 548838 183922 548894 183978
rect 548962 183922 549018 183978
rect 375228 175252 375284 175258
rect 375228 175202 375284 175252
rect 417564 173942 417620 173998
rect 374154 166294 374210 166350
rect 374278 166294 374334 166350
rect 374402 166294 374458 166350
rect 374526 166294 374582 166350
rect 374154 166170 374210 166226
rect 374278 166170 374334 166226
rect 374402 166170 374458 166226
rect 374526 166170 374582 166226
rect 374154 166046 374210 166102
rect 374278 166046 374334 166102
rect 374402 166046 374458 166102
rect 374526 166046 374582 166102
rect 374154 165922 374210 165978
rect 374278 165922 374334 165978
rect 374402 165922 374458 165978
rect 374526 165922 374582 165978
rect 374154 148294 374210 148350
rect 374278 148294 374334 148350
rect 374402 148294 374458 148350
rect 374526 148294 374582 148350
rect 374154 148170 374210 148226
rect 374278 148170 374334 148226
rect 374402 148170 374458 148226
rect 374526 148170 374582 148226
rect 374154 148046 374210 148102
rect 374278 148046 374334 148102
rect 374402 148046 374458 148102
rect 374526 148046 374582 148102
rect 374154 147922 374210 147978
rect 374278 147922 374334 147978
rect 374402 147922 374458 147978
rect 374526 147922 374582 147978
rect 374154 130294 374210 130350
rect 374278 130294 374334 130350
rect 374402 130294 374458 130350
rect 374526 130294 374582 130350
rect 374154 130170 374210 130226
rect 374278 130170 374334 130226
rect 374402 130170 374458 130226
rect 374526 130170 374582 130226
rect 374154 130046 374210 130102
rect 374278 130046 374334 130102
rect 374402 130046 374458 130102
rect 374526 130046 374582 130102
rect 374154 129922 374210 129978
rect 374278 129922 374334 129978
rect 374402 129922 374458 129978
rect 374526 129922 374582 129978
rect 359884 115802 359940 115858
rect 377874 172294 377930 172350
rect 377998 172294 378054 172350
rect 378122 172294 378178 172350
rect 378246 172294 378302 172350
rect 377874 172170 377930 172226
rect 377998 172170 378054 172226
rect 378122 172170 378178 172226
rect 378246 172170 378302 172226
rect 377874 172046 377930 172102
rect 377998 172046 378054 172102
rect 378122 172046 378178 172102
rect 378246 172046 378302 172102
rect 377874 171922 377930 171978
rect 377998 171922 378054 171978
rect 378122 171922 378178 171978
rect 378246 171922 378302 171978
rect 377874 154294 377930 154350
rect 377998 154294 378054 154350
rect 378122 154294 378178 154350
rect 378246 154294 378302 154350
rect 377874 154170 377930 154226
rect 377998 154170 378054 154226
rect 378122 154170 378178 154226
rect 378246 154170 378302 154226
rect 377874 154046 377930 154102
rect 377998 154046 378054 154102
rect 378122 154046 378178 154102
rect 378246 154046 378302 154102
rect 377874 153922 377930 153978
rect 377998 153922 378054 153978
rect 378122 153922 378178 153978
rect 378246 153922 378302 153978
rect 377874 136294 377930 136350
rect 377998 136294 378054 136350
rect 378122 136294 378178 136350
rect 378246 136294 378302 136350
rect 377874 136170 377930 136226
rect 377998 136170 378054 136226
rect 378122 136170 378178 136226
rect 378246 136170 378302 136226
rect 377874 136046 377930 136102
rect 377998 136046 378054 136102
rect 378122 136046 378178 136102
rect 378246 136046 378302 136102
rect 377874 135922 377930 135978
rect 377998 135922 378054 135978
rect 378122 135922 378178 135978
rect 378246 135922 378302 135978
rect 404874 166294 404930 166350
rect 404998 166294 405054 166350
rect 405122 166294 405178 166350
rect 405246 166294 405302 166350
rect 404874 166170 404930 166226
rect 404998 166170 405054 166226
rect 405122 166170 405178 166226
rect 405246 166170 405302 166226
rect 404874 166046 404930 166102
rect 404998 166046 405054 166102
rect 405122 166046 405178 166102
rect 405246 166046 405302 166102
rect 404874 165922 404930 165978
rect 404998 165922 405054 165978
rect 405122 165922 405178 165978
rect 405246 165922 405302 165978
rect 404874 148294 404930 148350
rect 404998 148294 405054 148350
rect 405122 148294 405178 148350
rect 405246 148294 405302 148350
rect 404874 148170 404930 148226
rect 404998 148170 405054 148226
rect 405122 148170 405178 148226
rect 405246 148170 405302 148226
rect 404874 148046 404930 148102
rect 404998 148046 405054 148102
rect 405122 148046 405178 148102
rect 405246 148046 405302 148102
rect 404874 147922 404930 147978
rect 404998 147922 405054 147978
rect 405122 147922 405178 147978
rect 405246 147922 405302 147978
rect 404874 130294 404930 130350
rect 404998 130294 405054 130350
rect 405122 130294 405178 130350
rect 405246 130294 405302 130350
rect 404874 130170 404930 130226
rect 404998 130170 405054 130226
rect 405122 130170 405178 130226
rect 405246 130170 405302 130226
rect 404874 130046 404930 130102
rect 404998 130046 405054 130102
rect 405122 130046 405178 130102
rect 405246 130046 405302 130102
rect 404874 129922 404930 129978
rect 404998 129922 405054 129978
rect 405122 129922 405178 129978
rect 405246 129922 405302 129978
rect 394940 124262 394996 124318
rect 388892 124082 388948 124138
rect 386876 123722 386932 123778
rect 384860 123542 384916 123598
rect 390908 123902 390964 123958
rect 377874 118294 377930 118350
rect 377998 118294 378054 118350
rect 378122 118294 378178 118350
rect 378246 118294 378302 118350
rect 377874 118170 377930 118226
rect 377998 118170 378054 118226
rect 378122 118170 378178 118226
rect 378246 118170 378302 118226
rect 377874 118046 377930 118102
rect 377998 118046 378054 118102
rect 378122 118046 378178 118102
rect 378246 118046 378302 118102
rect 377874 117922 377930 117978
rect 377998 117922 378054 117978
rect 378122 117922 378178 117978
rect 378246 117922 378302 117978
rect 408594 172294 408650 172350
rect 408718 172294 408774 172350
rect 408842 172294 408898 172350
rect 408966 172294 409022 172350
rect 408594 172170 408650 172226
rect 408718 172170 408774 172226
rect 408842 172170 408898 172226
rect 408966 172170 409022 172226
rect 408594 172046 408650 172102
rect 408718 172046 408774 172102
rect 408842 172046 408898 172102
rect 408966 172046 409022 172102
rect 408594 171922 408650 171978
rect 408718 171922 408774 171978
rect 408842 171922 408898 171978
rect 408966 171922 409022 171978
rect 408594 154294 408650 154350
rect 408718 154294 408774 154350
rect 408842 154294 408898 154350
rect 408966 154294 409022 154350
rect 408594 154170 408650 154226
rect 408718 154170 408774 154226
rect 408842 154170 408898 154226
rect 408966 154170 409022 154226
rect 408594 154046 408650 154102
rect 408718 154046 408774 154102
rect 408842 154046 408898 154102
rect 408966 154046 409022 154102
rect 408594 153922 408650 153978
rect 408718 153922 408774 153978
rect 408842 153922 408898 153978
rect 408966 153922 409022 153978
rect 435594 166294 435650 166350
rect 435718 166294 435774 166350
rect 435842 166294 435898 166350
rect 435966 166294 436022 166350
rect 435594 166170 435650 166226
rect 435718 166170 435774 166226
rect 435842 166170 435898 166226
rect 435966 166170 436022 166226
rect 435594 166046 435650 166102
rect 435718 166046 435774 166102
rect 435842 166046 435898 166102
rect 435966 166046 436022 166102
rect 435594 165922 435650 165978
rect 435718 165922 435774 165978
rect 435842 165922 435898 165978
rect 435966 165922 436022 165978
rect 435594 148294 435650 148350
rect 435718 148294 435774 148350
rect 435842 148294 435898 148350
rect 435966 148294 436022 148350
rect 435594 148170 435650 148226
rect 435718 148170 435774 148226
rect 435842 148170 435898 148226
rect 435966 148170 436022 148226
rect 435594 148046 435650 148102
rect 435718 148046 435774 148102
rect 435842 148046 435898 148102
rect 435966 148046 436022 148102
rect 435594 147922 435650 147978
rect 435718 147922 435774 147978
rect 435842 147922 435898 147978
rect 435966 147922 436022 147978
rect 408594 136294 408650 136350
rect 408718 136294 408774 136350
rect 408842 136294 408898 136350
rect 408966 136294 409022 136350
rect 408594 136170 408650 136226
rect 408718 136170 408774 136226
rect 408842 136170 408898 136226
rect 408966 136170 409022 136226
rect 408594 136046 408650 136102
rect 408718 136046 408774 136102
rect 408842 136046 408898 136102
rect 408966 136046 409022 136102
rect 408594 135922 408650 135978
rect 408718 135922 408774 135978
rect 408842 135922 408898 135978
rect 408966 135922 409022 135978
rect 414988 136862 415044 136918
rect 411628 133442 411684 133498
rect 435594 130294 435650 130350
rect 435718 130294 435774 130350
rect 435842 130294 435898 130350
rect 435966 130294 436022 130350
rect 435594 130170 435650 130226
rect 435718 130170 435774 130226
rect 435842 130170 435898 130226
rect 435966 130170 436022 130226
rect 435594 130046 435650 130102
rect 435718 130046 435774 130102
rect 435842 130046 435898 130102
rect 435966 130046 436022 130102
rect 435594 129922 435650 129978
rect 435718 129922 435774 129978
rect 435842 129922 435898 129978
rect 435966 129922 436022 129978
rect 408594 118294 408650 118350
rect 408718 118294 408774 118350
rect 408842 118294 408898 118350
rect 408966 118294 409022 118350
rect 408594 118170 408650 118226
rect 408718 118170 408774 118226
rect 408842 118170 408898 118226
rect 408966 118170 409022 118226
rect 408594 118046 408650 118102
rect 408718 118046 408774 118102
rect 408842 118046 408898 118102
rect 408966 118046 409022 118102
rect 408594 117922 408650 117978
rect 408718 117922 408774 117978
rect 408842 117922 408898 117978
rect 408966 117922 409022 117978
rect 364518 112294 364574 112350
rect 364642 112294 364698 112350
rect 364518 112170 364574 112226
rect 364642 112170 364698 112226
rect 364518 112046 364574 112102
rect 364642 112046 364698 112102
rect 364518 111922 364574 111978
rect 364642 111922 364698 111978
rect 395238 112294 395294 112350
rect 395362 112294 395418 112350
rect 395238 112170 395294 112226
rect 395362 112170 395418 112226
rect 395238 112046 395294 112102
rect 395362 112046 395418 112102
rect 395238 111922 395294 111978
rect 395362 111922 395418 111978
rect 379878 100294 379934 100350
rect 380002 100294 380058 100350
rect 379878 100170 379934 100226
rect 380002 100170 380058 100226
rect 379878 100046 379934 100102
rect 380002 100046 380058 100102
rect 379878 99922 379934 99978
rect 380002 99922 380058 99978
rect 410598 100294 410654 100350
rect 410722 100294 410778 100350
rect 410598 100170 410654 100226
rect 410722 100170 410778 100226
rect 410598 100046 410654 100102
rect 410722 100046 410778 100102
rect 410598 99922 410654 99978
rect 410722 99922 410778 99978
rect 364518 94294 364574 94350
rect 364642 94294 364698 94350
rect 364518 94170 364574 94226
rect 364642 94170 364698 94226
rect 364518 94046 364574 94102
rect 364642 94046 364698 94102
rect 364518 93922 364574 93978
rect 364642 93922 364698 93978
rect 395238 94294 395294 94350
rect 395362 94294 395418 94350
rect 395238 94170 395294 94226
rect 395362 94170 395418 94226
rect 395238 94046 395294 94102
rect 395362 94046 395418 94102
rect 395238 93922 395294 93978
rect 395362 93922 395418 93978
rect 379878 82294 379934 82350
rect 380002 82294 380058 82350
rect 379878 82170 379934 82226
rect 380002 82170 380058 82226
rect 379878 82046 379934 82102
rect 380002 82046 380058 82102
rect 379878 81922 379934 81978
rect 380002 81922 380058 81978
rect 410598 82294 410654 82350
rect 410722 82294 410778 82350
rect 410598 82170 410654 82226
rect 410722 82170 410778 82226
rect 410598 82046 410654 82102
rect 410722 82046 410778 82102
rect 410598 81922 410654 81978
rect 410722 81922 410778 81978
rect 364518 76294 364574 76350
rect 364642 76294 364698 76350
rect 364518 76170 364574 76226
rect 364642 76170 364698 76226
rect 364518 76046 364574 76102
rect 364642 76046 364698 76102
rect 364518 75922 364574 75978
rect 364642 75922 364698 75978
rect 395238 76294 395294 76350
rect 395362 76294 395418 76350
rect 395238 76170 395294 76226
rect 395362 76170 395418 76226
rect 395238 76046 395294 76102
rect 395362 76046 395418 76102
rect 395238 75922 395294 75978
rect 395362 75922 395418 75978
rect 379878 64294 379934 64350
rect 380002 64294 380058 64350
rect 379878 64170 379934 64226
rect 380002 64170 380058 64226
rect 379878 64046 379934 64102
rect 380002 64046 380058 64102
rect 379878 63922 379934 63978
rect 380002 63922 380058 63978
rect 410598 64294 410654 64350
rect 410722 64294 410778 64350
rect 410598 64170 410654 64226
rect 410722 64170 410778 64226
rect 410598 64046 410654 64102
rect 410722 64046 410778 64102
rect 410598 63922 410654 63978
rect 410722 63922 410778 63978
rect 435594 112294 435650 112350
rect 435718 112294 435774 112350
rect 435842 112294 435898 112350
rect 435966 112294 436022 112350
rect 435594 112170 435650 112226
rect 435718 112170 435774 112226
rect 435842 112170 435898 112226
rect 435966 112170 436022 112226
rect 435594 112046 435650 112102
rect 435718 112046 435774 112102
rect 435842 112046 435898 112102
rect 435966 112046 436022 112102
rect 435594 111922 435650 111978
rect 435718 111922 435774 111978
rect 435842 111922 435898 111978
rect 435966 111922 436022 111978
rect 435594 94294 435650 94350
rect 435718 94294 435774 94350
rect 435842 94294 435898 94350
rect 435966 94294 436022 94350
rect 435594 94170 435650 94226
rect 435718 94170 435774 94226
rect 435842 94170 435898 94226
rect 435966 94170 436022 94226
rect 435594 94046 435650 94102
rect 435718 94046 435774 94102
rect 435842 94046 435898 94102
rect 435966 94046 436022 94102
rect 435594 93922 435650 93978
rect 435718 93922 435774 93978
rect 435842 93922 435898 93978
rect 435966 93922 436022 93978
rect 435594 76294 435650 76350
rect 435718 76294 435774 76350
rect 435842 76294 435898 76350
rect 435966 76294 436022 76350
rect 435594 76170 435650 76226
rect 435718 76170 435774 76226
rect 435842 76170 435898 76226
rect 435966 76170 436022 76226
rect 435594 76046 435650 76102
rect 435718 76046 435774 76102
rect 435842 76046 435898 76102
rect 435966 76046 436022 76102
rect 435594 75922 435650 75978
rect 435718 75922 435774 75978
rect 435842 75922 435898 75978
rect 435966 75922 436022 75978
rect 364518 58294 364574 58350
rect 364642 58294 364698 58350
rect 364518 58170 364574 58226
rect 364642 58170 364698 58226
rect 364518 58046 364574 58102
rect 364642 58046 364698 58102
rect 364518 57922 364574 57978
rect 364642 57922 364698 57978
rect 395238 58294 395294 58350
rect 395362 58294 395418 58350
rect 395238 58170 395294 58226
rect 395362 58170 395418 58226
rect 395238 58046 395294 58102
rect 395362 58046 395418 58102
rect 395238 57922 395294 57978
rect 395362 57922 395418 57978
rect 435594 58294 435650 58350
rect 435718 58294 435774 58350
rect 435842 58294 435898 58350
rect 435966 58294 436022 58350
rect 435594 58170 435650 58226
rect 435718 58170 435774 58226
rect 435842 58170 435898 58226
rect 435966 58170 436022 58226
rect 435594 58046 435650 58102
rect 435718 58046 435774 58102
rect 435842 58046 435898 58102
rect 435966 58046 436022 58102
rect 435594 57922 435650 57978
rect 435718 57922 435774 57978
rect 435842 57922 435898 57978
rect 435966 57922 436022 57978
rect 347154 28294 347210 28350
rect 347278 28294 347334 28350
rect 347402 28294 347458 28350
rect 347526 28294 347582 28350
rect 347154 28170 347210 28226
rect 347278 28170 347334 28226
rect 347402 28170 347458 28226
rect 347526 28170 347582 28226
rect 347154 28046 347210 28102
rect 347278 28046 347334 28102
rect 347402 28046 347458 28102
rect 347526 28046 347582 28102
rect 347154 27922 347210 27978
rect 347278 27922 347334 27978
rect 347402 27922 347458 27978
rect 347526 27922 347582 27978
rect 347154 10294 347210 10350
rect 347278 10294 347334 10350
rect 347402 10294 347458 10350
rect 347526 10294 347582 10350
rect 347154 10170 347210 10226
rect 347278 10170 347334 10226
rect 347402 10170 347458 10226
rect 347526 10170 347582 10226
rect 347154 10046 347210 10102
rect 347278 10046 347334 10102
rect 347402 10046 347458 10102
rect 347526 10046 347582 10102
rect 347154 9922 347210 9978
rect 347278 9922 347334 9978
rect 347402 9922 347458 9978
rect 347526 9922 347582 9978
rect 347154 -1176 347210 -1120
rect 347278 -1176 347334 -1120
rect 347402 -1176 347458 -1120
rect 347526 -1176 347582 -1120
rect 347154 -1300 347210 -1244
rect 347278 -1300 347334 -1244
rect 347402 -1300 347458 -1244
rect 347526 -1300 347582 -1244
rect 347154 -1424 347210 -1368
rect 347278 -1424 347334 -1368
rect 347402 -1424 347458 -1368
rect 347526 -1424 347582 -1368
rect 347154 -1548 347210 -1492
rect 347278 -1548 347334 -1492
rect 347402 -1548 347458 -1492
rect 347526 -1548 347582 -1492
rect 374154 40294 374210 40350
rect 374278 40294 374334 40350
rect 374402 40294 374458 40350
rect 374526 40294 374582 40350
rect 374154 40170 374210 40226
rect 374278 40170 374334 40226
rect 374402 40170 374458 40226
rect 374526 40170 374582 40226
rect 374154 40046 374210 40102
rect 374278 40046 374334 40102
rect 374402 40046 374458 40102
rect 374526 40046 374582 40102
rect 374154 39922 374210 39978
rect 374278 39922 374334 39978
rect 374402 39922 374458 39978
rect 374526 39922 374582 39978
rect 374154 22294 374210 22350
rect 374278 22294 374334 22350
rect 374402 22294 374458 22350
rect 374526 22294 374582 22350
rect 374154 22170 374210 22226
rect 374278 22170 374334 22226
rect 374402 22170 374458 22226
rect 374526 22170 374582 22226
rect 374154 22046 374210 22102
rect 374278 22046 374334 22102
rect 374402 22046 374458 22102
rect 374526 22046 374582 22102
rect 374154 21922 374210 21978
rect 374278 21922 374334 21978
rect 374402 21922 374458 21978
rect 374526 21922 374582 21978
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 377874 46294 377930 46350
rect 377998 46294 378054 46350
rect 378122 46294 378178 46350
rect 378246 46294 378302 46350
rect 377874 46170 377930 46226
rect 377998 46170 378054 46226
rect 378122 46170 378178 46226
rect 378246 46170 378302 46226
rect 377874 46046 377930 46102
rect 377998 46046 378054 46102
rect 378122 46046 378178 46102
rect 378246 46046 378302 46102
rect 377874 45922 377930 45978
rect 377998 45922 378054 45978
rect 378122 45922 378178 45978
rect 378246 45922 378302 45978
rect 377874 28294 377930 28350
rect 377998 28294 378054 28350
rect 378122 28294 378178 28350
rect 378246 28294 378302 28350
rect 377874 28170 377930 28226
rect 377998 28170 378054 28226
rect 378122 28170 378178 28226
rect 378246 28170 378302 28226
rect 377874 28046 377930 28102
rect 377998 28046 378054 28102
rect 378122 28046 378178 28102
rect 378246 28046 378302 28102
rect 377874 27922 377930 27978
rect 377998 27922 378054 27978
rect 378122 27922 378178 27978
rect 378246 27922 378302 27978
rect 377874 10294 377930 10350
rect 377998 10294 378054 10350
rect 378122 10294 378178 10350
rect 378246 10294 378302 10350
rect 377874 10170 377930 10226
rect 377998 10170 378054 10226
rect 378122 10170 378178 10226
rect 378246 10170 378302 10226
rect 377874 10046 377930 10102
rect 377998 10046 378054 10102
rect 378122 10046 378178 10102
rect 378246 10046 378302 10102
rect 377874 9922 377930 9978
rect 377998 9922 378054 9978
rect 378122 9922 378178 9978
rect 378246 9922 378302 9978
rect 377874 -1176 377930 -1120
rect 377998 -1176 378054 -1120
rect 378122 -1176 378178 -1120
rect 378246 -1176 378302 -1120
rect 377874 -1300 377930 -1244
rect 377998 -1300 378054 -1244
rect 378122 -1300 378178 -1244
rect 378246 -1300 378302 -1244
rect 377874 -1424 377930 -1368
rect 377998 -1424 378054 -1368
rect 378122 -1424 378178 -1368
rect 378246 -1424 378302 -1368
rect 377874 -1548 377930 -1492
rect 377998 -1548 378054 -1492
rect 378122 -1548 378178 -1492
rect 378246 -1548 378302 -1492
rect 404874 40294 404930 40350
rect 404998 40294 405054 40350
rect 405122 40294 405178 40350
rect 405246 40294 405302 40350
rect 404874 40170 404930 40226
rect 404998 40170 405054 40226
rect 405122 40170 405178 40226
rect 405246 40170 405302 40226
rect 404874 40046 404930 40102
rect 404998 40046 405054 40102
rect 405122 40046 405178 40102
rect 405246 40046 405302 40102
rect 404874 39922 404930 39978
rect 404998 39922 405054 39978
rect 405122 39922 405178 39978
rect 405246 39922 405302 39978
rect 404874 22294 404930 22350
rect 404998 22294 405054 22350
rect 405122 22294 405178 22350
rect 405246 22294 405302 22350
rect 404874 22170 404930 22226
rect 404998 22170 405054 22226
rect 405122 22170 405178 22226
rect 405246 22170 405302 22226
rect 404874 22046 404930 22102
rect 404998 22046 405054 22102
rect 405122 22046 405178 22102
rect 405246 22046 405302 22102
rect 404874 21922 404930 21978
rect 404998 21922 405054 21978
rect 405122 21922 405178 21978
rect 405246 21922 405302 21978
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 408594 46294 408650 46350
rect 408718 46294 408774 46350
rect 408842 46294 408898 46350
rect 408966 46294 409022 46350
rect 408594 46170 408650 46226
rect 408718 46170 408774 46226
rect 408842 46170 408898 46226
rect 408966 46170 409022 46226
rect 408594 46046 408650 46102
rect 408718 46046 408774 46102
rect 408842 46046 408898 46102
rect 408966 46046 409022 46102
rect 408594 45922 408650 45978
rect 408718 45922 408774 45978
rect 408842 45922 408898 45978
rect 408966 45922 409022 45978
rect 408594 28294 408650 28350
rect 408718 28294 408774 28350
rect 408842 28294 408898 28350
rect 408966 28294 409022 28350
rect 408594 28170 408650 28226
rect 408718 28170 408774 28226
rect 408842 28170 408898 28226
rect 408966 28170 409022 28226
rect 408594 28046 408650 28102
rect 408718 28046 408774 28102
rect 408842 28046 408898 28102
rect 408966 28046 409022 28102
rect 408594 27922 408650 27978
rect 408718 27922 408774 27978
rect 408842 27922 408898 27978
rect 408966 27922 409022 27978
rect 408594 10294 408650 10350
rect 408718 10294 408774 10350
rect 408842 10294 408898 10350
rect 408966 10294 409022 10350
rect 408594 10170 408650 10226
rect 408718 10170 408774 10226
rect 408842 10170 408898 10226
rect 408966 10170 409022 10226
rect 408594 10046 408650 10102
rect 408718 10046 408774 10102
rect 408842 10046 408898 10102
rect 408966 10046 409022 10102
rect 408594 9922 408650 9978
rect 408718 9922 408774 9978
rect 408842 9922 408898 9978
rect 408966 9922 409022 9978
rect 408594 -1176 408650 -1120
rect 408718 -1176 408774 -1120
rect 408842 -1176 408898 -1120
rect 408966 -1176 409022 -1120
rect 408594 -1300 408650 -1244
rect 408718 -1300 408774 -1244
rect 408842 -1300 408898 -1244
rect 408966 -1300 409022 -1244
rect 408594 -1424 408650 -1368
rect 408718 -1424 408774 -1368
rect 408842 -1424 408898 -1368
rect 408966 -1424 409022 -1368
rect 408594 -1548 408650 -1492
rect 408718 -1548 408774 -1492
rect 408842 -1548 408898 -1492
rect 408966 -1548 409022 -1492
rect 435594 40294 435650 40350
rect 435718 40294 435774 40350
rect 435842 40294 435898 40350
rect 435966 40294 436022 40350
rect 435594 40170 435650 40226
rect 435718 40170 435774 40226
rect 435842 40170 435898 40226
rect 435966 40170 436022 40226
rect 435594 40046 435650 40102
rect 435718 40046 435774 40102
rect 435842 40046 435898 40102
rect 435966 40046 436022 40102
rect 435594 39922 435650 39978
rect 435718 39922 435774 39978
rect 435842 39922 435898 39978
rect 435966 39922 436022 39978
rect 435594 22294 435650 22350
rect 435718 22294 435774 22350
rect 435842 22294 435898 22350
rect 435966 22294 436022 22350
rect 435594 22170 435650 22226
rect 435718 22170 435774 22226
rect 435842 22170 435898 22226
rect 435966 22170 436022 22226
rect 435594 22046 435650 22102
rect 435718 22046 435774 22102
rect 435842 22046 435898 22102
rect 435966 22046 436022 22102
rect 435594 21922 435650 21978
rect 435718 21922 435774 21978
rect 435842 21922 435898 21978
rect 435966 21922 436022 21978
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 439314 172294 439370 172350
rect 439438 172294 439494 172350
rect 439562 172294 439618 172350
rect 439686 172294 439742 172350
rect 439314 172170 439370 172226
rect 439438 172170 439494 172226
rect 439562 172170 439618 172226
rect 439686 172170 439742 172226
rect 439314 172046 439370 172102
rect 439438 172046 439494 172102
rect 439562 172046 439618 172102
rect 439686 172046 439742 172102
rect 439314 171922 439370 171978
rect 439438 171922 439494 171978
rect 439562 171922 439618 171978
rect 439686 171922 439742 171978
rect 470034 172294 470090 172350
rect 470158 172294 470214 172350
rect 470282 172294 470338 172350
rect 470406 172294 470462 172350
rect 470034 172170 470090 172226
rect 470158 172170 470214 172226
rect 470282 172170 470338 172226
rect 470406 172170 470462 172226
rect 470034 172046 470090 172102
rect 470158 172046 470214 172102
rect 470282 172046 470338 172102
rect 470406 172046 470462 172102
rect 470034 171922 470090 171978
rect 470158 171922 470214 171978
rect 470282 171922 470338 171978
rect 470406 171922 470462 171978
rect 439314 154294 439370 154350
rect 439438 154294 439494 154350
rect 439562 154294 439618 154350
rect 439686 154294 439742 154350
rect 439314 154170 439370 154226
rect 439438 154170 439494 154226
rect 439562 154170 439618 154226
rect 439686 154170 439742 154226
rect 439314 154046 439370 154102
rect 439438 154046 439494 154102
rect 439562 154046 439618 154102
rect 439686 154046 439742 154102
rect 439314 153922 439370 153978
rect 439438 153922 439494 153978
rect 439562 153922 439618 153978
rect 439686 153922 439742 153978
rect 439314 136294 439370 136350
rect 439438 136294 439494 136350
rect 439562 136294 439618 136350
rect 439686 136294 439742 136350
rect 439314 136170 439370 136226
rect 439438 136170 439494 136226
rect 439562 136170 439618 136226
rect 439686 136170 439742 136226
rect 439314 136046 439370 136102
rect 439438 136046 439494 136102
rect 439562 136046 439618 136102
rect 439686 136046 439742 136102
rect 439314 135922 439370 135978
rect 439438 135922 439494 135978
rect 439562 135922 439618 135978
rect 439686 135922 439742 135978
rect 439314 118294 439370 118350
rect 439438 118294 439494 118350
rect 439562 118294 439618 118350
rect 439686 118294 439742 118350
rect 439314 118170 439370 118226
rect 439438 118170 439494 118226
rect 439562 118170 439618 118226
rect 439686 118170 439742 118226
rect 439314 118046 439370 118102
rect 439438 118046 439494 118102
rect 439562 118046 439618 118102
rect 439686 118046 439742 118102
rect 439314 117922 439370 117978
rect 439438 117922 439494 117978
rect 439562 117922 439618 117978
rect 439686 117922 439742 117978
rect 457660 115836 457716 115858
rect 457660 115802 457716 115836
rect 439314 100294 439370 100350
rect 439438 100294 439494 100350
rect 439562 100294 439618 100350
rect 439686 100294 439742 100350
rect 439314 100170 439370 100226
rect 439438 100170 439494 100226
rect 439562 100170 439618 100226
rect 439686 100170 439742 100226
rect 439314 100046 439370 100102
rect 439438 100046 439494 100102
rect 439562 100046 439618 100102
rect 439686 100046 439742 100102
rect 439314 99922 439370 99978
rect 439438 99922 439494 99978
rect 439562 99922 439618 99978
rect 439686 99922 439742 99978
rect 439314 82294 439370 82350
rect 439438 82294 439494 82350
rect 439562 82294 439618 82350
rect 439686 82294 439742 82350
rect 439314 82170 439370 82226
rect 439438 82170 439494 82226
rect 439562 82170 439618 82226
rect 439686 82170 439742 82226
rect 439314 82046 439370 82102
rect 439438 82046 439494 82102
rect 439562 82046 439618 82102
rect 439686 82046 439742 82102
rect 439314 81922 439370 81978
rect 439438 81922 439494 81978
rect 439562 81922 439618 81978
rect 439686 81922 439742 81978
rect 490588 173042 490644 173098
rect 470034 154294 470090 154350
rect 470158 154294 470214 154350
rect 470282 154294 470338 154350
rect 470406 154294 470462 154350
rect 470034 154170 470090 154226
rect 470158 154170 470214 154226
rect 470282 154170 470338 154226
rect 470406 154170 470462 154226
rect 470034 154046 470090 154102
rect 470158 154046 470214 154102
rect 470282 154046 470338 154102
rect 470406 154046 470462 154102
rect 488908 168722 488964 168778
rect 500754 172294 500810 172350
rect 500878 172294 500934 172350
rect 501002 172294 501058 172350
rect 501126 172294 501182 172350
rect 500754 172170 500810 172226
rect 500878 172170 500934 172226
rect 501002 172170 501058 172226
rect 501126 172170 501182 172226
rect 500754 172046 500810 172102
rect 500878 172046 500934 172102
rect 501002 172046 501058 172102
rect 501126 172046 501182 172102
rect 500754 171922 500810 171978
rect 500878 171922 500934 171978
rect 501002 171922 501058 171978
rect 501126 171922 501182 171978
rect 493164 157022 493220 157078
rect 470034 153922 470090 153978
rect 470158 153922 470214 153978
rect 470282 153922 470338 153978
rect 470406 153922 470462 153978
rect 500754 154294 500810 154350
rect 500878 154294 500934 154350
rect 501002 154294 501058 154350
rect 501126 154294 501182 154350
rect 500754 154170 500810 154226
rect 500878 154170 500934 154226
rect 501002 154170 501058 154226
rect 501126 154170 501182 154226
rect 500754 154046 500810 154102
rect 500878 154046 500934 154102
rect 501002 154046 501058 154102
rect 501126 154046 501182 154102
rect 500754 153922 500810 153978
rect 500878 153922 500934 153978
rect 501002 153922 501058 153978
rect 501126 153922 501182 153978
rect 482076 150542 482132 150598
rect 559580 395342 559636 395398
rect 568652 411002 568708 411058
rect 566972 408122 567028 408178
rect 565292 404342 565348 404398
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 584668 409382 584724 409438
rect 585452 409022 585508 409078
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 570332 404162 570388 404218
rect 572012 402002 572068 402058
rect 562194 388294 562250 388350
rect 562318 388294 562374 388350
rect 562442 388294 562498 388350
rect 562566 388294 562622 388350
rect 562194 388170 562250 388226
rect 562318 388170 562374 388226
rect 562442 388170 562498 388226
rect 562566 388170 562622 388226
rect 562194 388046 562250 388102
rect 562318 388046 562374 388102
rect 562442 388046 562498 388102
rect 562566 388046 562622 388102
rect 562194 387922 562250 387978
rect 562318 387922 562374 387978
rect 562442 387922 562498 387978
rect 562566 387922 562622 387978
rect 562194 370294 562250 370350
rect 562318 370294 562374 370350
rect 562442 370294 562498 370350
rect 562566 370294 562622 370350
rect 562194 370170 562250 370226
rect 562318 370170 562374 370226
rect 562442 370170 562498 370226
rect 562566 370170 562622 370226
rect 562194 370046 562250 370102
rect 562318 370046 562374 370102
rect 562442 370046 562498 370102
rect 562566 370046 562622 370102
rect 562194 369922 562250 369978
rect 562318 369922 562374 369978
rect 562442 369922 562498 369978
rect 562566 369922 562622 369978
rect 562194 352294 562250 352350
rect 562318 352294 562374 352350
rect 562442 352294 562498 352350
rect 562566 352294 562622 352350
rect 562194 352170 562250 352226
rect 562318 352170 562374 352226
rect 562442 352170 562498 352226
rect 562566 352170 562622 352226
rect 562194 352046 562250 352102
rect 562318 352046 562374 352102
rect 562442 352046 562498 352102
rect 562566 352046 562622 352102
rect 562194 351922 562250 351978
rect 562318 351922 562374 351978
rect 562442 351922 562498 351978
rect 562566 351922 562622 351978
rect 562194 334294 562250 334350
rect 562318 334294 562374 334350
rect 562442 334294 562498 334350
rect 562566 334294 562622 334350
rect 562194 334170 562250 334226
rect 562318 334170 562374 334226
rect 562442 334170 562498 334226
rect 562566 334170 562622 334226
rect 562194 334046 562250 334102
rect 562318 334046 562374 334102
rect 562442 334046 562498 334102
rect 562566 334046 562622 334102
rect 562194 333922 562250 333978
rect 562318 333922 562374 333978
rect 562442 333922 562498 333978
rect 562566 333922 562622 333978
rect 562194 316294 562250 316350
rect 562318 316294 562374 316350
rect 562442 316294 562498 316350
rect 562566 316294 562622 316350
rect 562194 316170 562250 316226
rect 562318 316170 562374 316226
rect 562442 316170 562498 316226
rect 562566 316170 562622 316226
rect 562194 316046 562250 316102
rect 562318 316046 562374 316102
rect 562442 316046 562498 316102
rect 562566 316046 562622 316102
rect 562194 315922 562250 315978
rect 562318 315922 562374 315978
rect 562442 315922 562498 315978
rect 562566 315922 562622 315978
rect 562194 298294 562250 298350
rect 562318 298294 562374 298350
rect 562442 298294 562498 298350
rect 562566 298294 562622 298350
rect 562194 298170 562250 298226
rect 562318 298170 562374 298226
rect 562442 298170 562498 298226
rect 562566 298170 562622 298226
rect 562194 298046 562250 298102
rect 562318 298046 562374 298102
rect 562442 298046 562498 298102
rect 562566 298046 562622 298102
rect 562194 297922 562250 297978
rect 562318 297922 562374 297978
rect 562442 297922 562498 297978
rect 562566 297922 562622 297978
rect 562194 280294 562250 280350
rect 562318 280294 562374 280350
rect 562442 280294 562498 280350
rect 562566 280294 562622 280350
rect 562194 280170 562250 280226
rect 562318 280170 562374 280226
rect 562442 280170 562498 280226
rect 562566 280170 562622 280226
rect 562194 280046 562250 280102
rect 562318 280046 562374 280102
rect 562442 280046 562498 280102
rect 562566 280046 562622 280102
rect 562194 279922 562250 279978
rect 562318 279922 562374 279978
rect 562442 279922 562498 279978
rect 562566 279922 562622 279978
rect 562194 262294 562250 262350
rect 562318 262294 562374 262350
rect 562442 262294 562498 262350
rect 562566 262294 562622 262350
rect 562194 262170 562250 262226
rect 562318 262170 562374 262226
rect 562442 262170 562498 262226
rect 562566 262170 562622 262226
rect 562194 262046 562250 262102
rect 562318 262046 562374 262102
rect 562442 262046 562498 262102
rect 562566 262046 562622 262102
rect 562194 261922 562250 261978
rect 562318 261922 562374 261978
rect 562442 261922 562498 261978
rect 562566 261922 562622 261978
rect 562194 244294 562250 244350
rect 562318 244294 562374 244350
rect 562442 244294 562498 244350
rect 562566 244294 562622 244350
rect 562194 244170 562250 244226
rect 562318 244170 562374 244226
rect 562442 244170 562498 244226
rect 562566 244170 562622 244226
rect 562194 244046 562250 244102
rect 562318 244046 562374 244102
rect 562442 244046 562498 244102
rect 562566 244046 562622 244102
rect 562194 243922 562250 243978
rect 562318 243922 562374 243978
rect 562442 243922 562498 243978
rect 562566 243922 562622 243978
rect 562194 226294 562250 226350
rect 562318 226294 562374 226350
rect 562442 226294 562498 226350
rect 562566 226294 562622 226350
rect 562194 226170 562250 226226
rect 562318 226170 562374 226226
rect 562442 226170 562498 226226
rect 562566 226170 562622 226226
rect 562194 226046 562250 226102
rect 562318 226046 562374 226102
rect 562442 226046 562498 226102
rect 562566 226046 562622 226102
rect 562194 225922 562250 225978
rect 562318 225922 562374 225978
rect 562442 225922 562498 225978
rect 562566 225922 562622 225978
rect 562194 208294 562250 208350
rect 562318 208294 562374 208350
rect 562442 208294 562498 208350
rect 562566 208294 562622 208350
rect 562194 208170 562250 208226
rect 562318 208170 562374 208226
rect 562442 208170 562498 208226
rect 562566 208170 562622 208226
rect 562194 208046 562250 208102
rect 562318 208046 562374 208102
rect 562442 208046 562498 208102
rect 562566 208046 562622 208102
rect 562194 207922 562250 207978
rect 562318 207922 562374 207978
rect 562442 207922 562498 207978
rect 562566 207922 562622 207978
rect 562194 190294 562250 190350
rect 562318 190294 562374 190350
rect 562442 190294 562498 190350
rect 562566 190294 562622 190350
rect 562194 190170 562250 190226
rect 562318 190170 562374 190226
rect 562442 190170 562498 190226
rect 562566 190170 562622 190226
rect 562194 190046 562250 190102
rect 562318 190046 562374 190102
rect 562442 190046 562498 190102
rect 562566 190046 562622 190102
rect 562194 189922 562250 189978
rect 562318 189922 562374 189978
rect 562442 189922 562498 189978
rect 562566 189922 562622 189978
rect 561148 173762 561204 173818
rect 531474 172294 531530 172350
rect 531598 172294 531654 172350
rect 531722 172294 531778 172350
rect 531846 172294 531902 172350
rect 531474 172170 531530 172226
rect 531598 172170 531654 172226
rect 531722 172170 531778 172226
rect 531846 172170 531902 172226
rect 531474 172046 531530 172102
rect 531598 172046 531654 172102
rect 531722 172046 531778 172102
rect 531846 172046 531902 172102
rect 531474 171922 531530 171978
rect 531598 171922 531654 171978
rect 531722 171922 531778 171978
rect 531846 171922 531902 171978
rect 531474 154294 531530 154350
rect 531598 154294 531654 154350
rect 531722 154294 531778 154350
rect 531846 154294 531902 154350
rect 531474 154170 531530 154226
rect 531598 154170 531654 154226
rect 531722 154170 531778 154226
rect 531846 154170 531902 154226
rect 531474 154046 531530 154102
rect 531598 154046 531654 154102
rect 531722 154046 531778 154102
rect 531846 154046 531902 154102
rect 531474 153922 531530 153978
rect 531598 153922 531654 153978
rect 531722 153922 531778 153978
rect 531846 153922 531902 153978
rect 502572 153602 502628 153658
rect 503132 153422 503188 153478
rect 463372 147662 463428 147718
rect 462028 146042 462084 146098
rect 479878 136294 479934 136350
rect 480002 136294 480058 136350
rect 479878 136170 479934 136226
rect 480002 136170 480058 136226
rect 479878 136046 479934 136102
rect 480002 136046 480058 136102
rect 479878 135922 479934 135978
rect 480002 135922 480058 135978
rect 510598 136294 510654 136350
rect 510722 136294 510778 136350
rect 510598 136170 510654 136226
rect 510722 136170 510778 136226
rect 510598 136046 510654 136102
rect 510722 136046 510778 136102
rect 510598 135922 510654 135978
rect 510722 135922 510778 135978
rect 541318 136294 541374 136350
rect 541442 136294 541498 136350
rect 541318 136170 541374 136226
rect 541442 136170 541498 136226
rect 541318 136046 541374 136102
rect 541442 136046 541498 136102
rect 541318 135922 541374 135978
rect 541442 135922 541498 135978
rect 464518 130294 464574 130350
rect 464642 130294 464698 130350
rect 464518 130170 464574 130226
rect 464642 130170 464698 130226
rect 464518 130046 464574 130102
rect 464642 130046 464698 130102
rect 464518 129922 464574 129978
rect 464642 129922 464698 129978
rect 495238 130294 495294 130350
rect 495362 130294 495418 130350
rect 495238 130170 495294 130226
rect 495362 130170 495418 130226
rect 495238 130046 495294 130102
rect 495362 130046 495418 130102
rect 495238 129922 495294 129978
rect 495362 129922 495418 129978
rect 525958 130294 526014 130350
rect 526082 130294 526138 130350
rect 525958 130170 526014 130226
rect 526082 130170 526138 130226
rect 525958 130046 526014 130102
rect 526082 130046 526138 130102
rect 525958 129922 526014 129978
rect 526082 129922 526138 129978
rect 556678 130294 556734 130350
rect 556802 130294 556858 130350
rect 556678 130170 556734 130226
rect 556802 130170 556858 130226
rect 556678 130046 556734 130102
rect 556802 130046 556858 130102
rect 556678 129922 556734 129978
rect 556802 129922 556858 129978
rect 479878 118294 479934 118350
rect 480002 118294 480058 118350
rect 479878 118170 479934 118226
rect 480002 118170 480058 118226
rect 479878 118046 479934 118102
rect 480002 118046 480058 118102
rect 479878 117922 479934 117978
rect 480002 117922 480058 117978
rect 510598 118294 510654 118350
rect 510722 118294 510778 118350
rect 510598 118170 510654 118226
rect 510722 118170 510778 118226
rect 510598 118046 510654 118102
rect 510722 118046 510778 118102
rect 510598 117922 510654 117978
rect 510722 117922 510778 117978
rect 541318 118294 541374 118350
rect 541442 118294 541498 118350
rect 541318 118170 541374 118226
rect 541442 118170 541498 118226
rect 541318 118046 541374 118102
rect 541442 118046 541498 118102
rect 541318 117922 541374 117978
rect 541442 117922 541498 117978
rect 464518 112294 464574 112350
rect 464642 112294 464698 112350
rect 464518 112170 464574 112226
rect 464642 112170 464698 112226
rect 464518 112046 464574 112102
rect 464642 112046 464698 112102
rect 464518 111922 464574 111978
rect 464642 111922 464698 111978
rect 495238 112294 495294 112350
rect 495362 112294 495418 112350
rect 495238 112170 495294 112226
rect 495362 112170 495418 112226
rect 495238 112046 495294 112102
rect 495362 112046 495418 112102
rect 495238 111922 495294 111978
rect 495362 111922 495418 111978
rect 525958 112294 526014 112350
rect 526082 112294 526138 112350
rect 525958 112170 526014 112226
rect 526082 112170 526138 112226
rect 525958 112046 526014 112102
rect 526082 112046 526138 112102
rect 525958 111922 526014 111978
rect 526082 111922 526138 111978
rect 556678 112294 556734 112350
rect 556802 112294 556858 112350
rect 556678 112170 556734 112226
rect 556802 112170 556858 112226
rect 556678 112046 556734 112102
rect 556802 112046 556858 112102
rect 556678 111922 556734 111978
rect 556802 111922 556858 111978
rect 479878 100294 479934 100350
rect 480002 100294 480058 100350
rect 479878 100170 479934 100226
rect 480002 100170 480058 100226
rect 479878 100046 479934 100102
rect 480002 100046 480058 100102
rect 479878 99922 479934 99978
rect 480002 99922 480058 99978
rect 510598 100294 510654 100350
rect 510722 100294 510778 100350
rect 510598 100170 510654 100226
rect 510722 100170 510778 100226
rect 510598 100046 510654 100102
rect 510722 100046 510778 100102
rect 510598 99922 510654 99978
rect 510722 99922 510778 99978
rect 541318 100294 541374 100350
rect 541442 100294 541498 100350
rect 541318 100170 541374 100226
rect 541442 100170 541498 100226
rect 541318 100046 541374 100102
rect 541442 100046 541498 100102
rect 541318 99922 541374 99978
rect 541442 99922 541498 99978
rect 464518 94294 464574 94350
rect 464642 94294 464698 94350
rect 464518 94170 464574 94226
rect 464642 94170 464698 94226
rect 464518 94046 464574 94102
rect 464642 94046 464698 94102
rect 464518 93922 464574 93978
rect 464642 93922 464698 93978
rect 495238 94294 495294 94350
rect 495362 94294 495418 94350
rect 495238 94170 495294 94226
rect 495362 94170 495418 94226
rect 495238 94046 495294 94102
rect 495362 94046 495418 94102
rect 495238 93922 495294 93978
rect 495362 93922 495418 93978
rect 525958 94294 526014 94350
rect 526082 94294 526138 94350
rect 525958 94170 526014 94226
rect 526082 94170 526138 94226
rect 525958 94046 526014 94102
rect 526082 94046 526138 94102
rect 525958 93922 526014 93978
rect 526082 93922 526138 93978
rect 556678 94294 556734 94350
rect 556802 94294 556858 94350
rect 556678 94170 556734 94226
rect 556802 94170 556858 94226
rect 556678 94046 556734 94102
rect 556802 94046 556858 94102
rect 556678 93922 556734 93978
rect 556802 93922 556858 93978
rect 479878 82294 479934 82350
rect 480002 82294 480058 82350
rect 479878 82170 479934 82226
rect 480002 82170 480058 82226
rect 479878 82046 479934 82102
rect 480002 82046 480058 82102
rect 479878 81922 479934 81978
rect 480002 81922 480058 81978
rect 510598 82294 510654 82350
rect 510722 82294 510778 82350
rect 510598 82170 510654 82226
rect 510722 82170 510778 82226
rect 510598 82046 510654 82102
rect 510722 82046 510778 82102
rect 510598 81922 510654 81978
rect 510722 81922 510778 81978
rect 541318 82294 541374 82350
rect 541442 82294 541498 82350
rect 541318 82170 541374 82226
rect 541442 82170 541498 82226
rect 541318 82046 541374 82102
rect 541442 82046 541498 82102
rect 541318 81922 541374 81978
rect 541442 81922 541498 81978
rect 464518 76294 464574 76350
rect 464642 76294 464698 76350
rect 464518 76170 464574 76226
rect 464642 76170 464698 76226
rect 464518 76046 464574 76102
rect 464642 76046 464698 76102
rect 464518 75922 464574 75978
rect 464642 75922 464698 75978
rect 495238 76294 495294 76350
rect 495362 76294 495418 76350
rect 495238 76170 495294 76226
rect 495362 76170 495418 76226
rect 495238 76046 495294 76102
rect 495362 76046 495418 76102
rect 495238 75922 495294 75978
rect 495362 75922 495418 75978
rect 525958 76294 526014 76350
rect 526082 76294 526138 76350
rect 525958 76170 526014 76226
rect 526082 76170 526138 76226
rect 525958 76046 526014 76102
rect 526082 76046 526138 76102
rect 525958 75922 526014 75978
rect 526082 75922 526138 75978
rect 556678 76294 556734 76350
rect 556802 76294 556858 76350
rect 556678 76170 556734 76226
rect 556802 76170 556858 76226
rect 556678 76046 556734 76102
rect 556802 76046 556858 76102
rect 556678 75922 556734 75978
rect 556802 75922 556858 75978
rect 559580 170522 559636 170578
rect 570332 393542 570388 393598
rect 562194 172294 562250 172350
rect 562318 172294 562374 172350
rect 562442 172294 562498 172350
rect 562566 172294 562622 172350
rect 562194 172170 562250 172226
rect 562318 172170 562374 172226
rect 562442 172170 562498 172226
rect 562566 172170 562622 172226
rect 562194 172046 562250 172102
rect 562318 172046 562374 172102
rect 562442 172046 562498 172102
rect 562566 172046 562622 172102
rect 562194 171922 562250 171978
rect 562318 171922 562374 171978
rect 562442 171922 562498 171978
rect 562566 171922 562622 171978
rect 561260 158822 561316 158878
rect 562194 154294 562250 154350
rect 562318 154294 562374 154350
rect 562442 154294 562498 154350
rect 562566 154294 562622 154350
rect 562194 154170 562250 154226
rect 562318 154170 562374 154226
rect 562442 154170 562498 154226
rect 562566 154170 562622 154226
rect 562194 154046 562250 154102
rect 562318 154046 562374 154102
rect 562442 154046 562498 154102
rect 562566 154046 562622 154102
rect 562194 153922 562250 153978
rect 562318 153922 562374 153978
rect 562442 153922 562498 153978
rect 562566 153922 562622 153978
rect 562194 136294 562250 136350
rect 562318 136294 562374 136350
rect 562442 136294 562498 136350
rect 562566 136294 562622 136350
rect 562194 136170 562250 136226
rect 562318 136170 562374 136226
rect 562442 136170 562498 136226
rect 562566 136170 562622 136226
rect 562194 136046 562250 136102
rect 562318 136046 562374 136102
rect 562442 136046 562498 136102
rect 562566 136046 562622 136102
rect 562194 135922 562250 135978
rect 562318 135922 562374 135978
rect 562442 135922 562498 135978
rect 562566 135922 562622 135978
rect 562194 118294 562250 118350
rect 562318 118294 562374 118350
rect 562442 118294 562498 118350
rect 562566 118294 562622 118350
rect 562194 118170 562250 118226
rect 562318 118170 562374 118226
rect 562442 118170 562498 118226
rect 562566 118170 562622 118226
rect 562194 118046 562250 118102
rect 562318 118046 562374 118102
rect 562442 118046 562498 118102
rect 562566 118046 562622 118102
rect 562194 117922 562250 117978
rect 562318 117922 562374 117978
rect 562442 117922 562498 117978
rect 562566 117922 562622 117978
rect 562194 100294 562250 100350
rect 562318 100294 562374 100350
rect 562442 100294 562498 100350
rect 562566 100294 562622 100350
rect 562194 100170 562250 100226
rect 562318 100170 562374 100226
rect 562442 100170 562498 100226
rect 562566 100170 562622 100226
rect 562194 100046 562250 100102
rect 562318 100046 562374 100102
rect 562442 100046 562498 100102
rect 562566 100046 562622 100102
rect 562194 99922 562250 99978
rect 562318 99922 562374 99978
rect 562442 99922 562498 99978
rect 562566 99922 562622 99978
rect 439314 64294 439370 64350
rect 439438 64294 439494 64350
rect 439562 64294 439618 64350
rect 439686 64294 439742 64350
rect 439314 64170 439370 64226
rect 439438 64170 439494 64226
rect 439562 64170 439618 64226
rect 439686 64170 439742 64226
rect 439314 64046 439370 64102
rect 439438 64046 439494 64102
rect 439562 64046 439618 64102
rect 439686 64046 439742 64102
rect 439314 63922 439370 63978
rect 439438 63922 439494 63978
rect 439562 63922 439618 63978
rect 439686 63922 439742 63978
rect 479878 64294 479934 64350
rect 480002 64294 480058 64350
rect 479878 64170 479934 64226
rect 480002 64170 480058 64226
rect 479878 64046 479934 64102
rect 480002 64046 480058 64102
rect 479878 63922 479934 63978
rect 480002 63922 480058 63978
rect 510598 64294 510654 64350
rect 510722 64294 510778 64350
rect 510598 64170 510654 64226
rect 510722 64170 510778 64226
rect 510598 64046 510654 64102
rect 510722 64046 510778 64102
rect 510598 63922 510654 63978
rect 510722 63922 510778 63978
rect 541318 64294 541374 64350
rect 541442 64294 541498 64350
rect 541318 64170 541374 64226
rect 541442 64170 541498 64226
rect 541318 64046 541374 64102
rect 541442 64046 541498 64102
rect 541318 63922 541374 63978
rect 541442 63922 541498 63978
rect 464518 58294 464574 58350
rect 464642 58294 464698 58350
rect 464518 58170 464574 58226
rect 464642 58170 464698 58226
rect 464518 58046 464574 58102
rect 464642 58046 464698 58102
rect 464518 57922 464574 57978
rect 464642 57922 464698 57978
rect 495238 58294 495294 58350
rect 495362 58294 495418 58350
rect 495238 58170 495294 58226
rect 495362 58170 495418 58226
rect 495238 58046 495294 58102
rect 495362 58046 495418 58102
rect 495238 57922 495294 57978
rect 495362 57922 495418 57978
rect 525958 58294 526014 58350
rect 526082 58294 526138 58350
rect 525958 58170 526014 58226
rect 526082 58170 526138 58226
rect 525958 58046 526014 58102
rect 526082 58046 526138 58102
rect 525958 57922 526014 57978
rect 526082 57922 526138 57978
rect 556678 58294 556734 58350
rect 556802 58294 556858 58350
rect 556678 58170 556734 58226
rect 556802 58170 556858 58226
rect 556678 58046 556734 58102
rect 556802 58046 556858 58102
rect 556678 57922 556734 57978
rect 556802 57922 556858 57978
rect 439314 46294 439370 46350
rect 439438 46294 439494 46350
rect 439562 46294 439618 46350
rect 439686 46294 439742 46350
rect 439314 46170 439370 46226
rect 439438 46170 439494 46226
rect 439562 46170 439618 46226
rect 439686 46170 439742 46226
rect 439314 46046 439370 46102
rect 439438 46046 439494 46102
rect 439562 46046 439618 46102
rect 439686 46046 439742 46102
rect 439314 45922 439370 45978
rect 439438 45922 439494 45978
rect 439562 45922 439618 45978
rect 439686 45922 439742 45978
rect 439314 28294 439370 28350
rect 439438 28294 439494 28350
rect 439562 28294 439618 28350
rect 439686 28294 439742 28350
rect 439314 28170 439370 28226
rect 439438 28170 439494 28226
rect 439562 28170 439618 28226
rect 439686 28170 439742 28226
rect 439314 28046 439370 28102
rect 439438 28046 439494 28102
rect 439562 28046 439618 28102
rect 439686 28046 439742 28102
rect 439314 27922 439370 27978
rect 439438 27922 439494 27978
rect 439562 27922 439618 27978
rect 439686 27922 439742 27978
rect 439314 10294 439370 10350
rect 439438 10294 439494 10350
rect 439562 10294 439618 10350
rect 439686 10294 439742 10350
rect 439314 10170 439370 10226
rect 439438 10170 439494 10226
rect 439562 10170 439618 10226
rect 439686 10170 439742 10226
rect 439314 10046 439370 10102
rect 439438 10046 439494 10102
rect 439562 10046 439618 10102
rect 439686 10046 439742 10102
rect 439314 9922 439370 9978
rect 439438 9922 439494 9978
rect 439562 9922 439618 9978
rect 439686 9922 439742 9978
rect 439314 -1176 439370 -1120
rect 439438 -1176 439494 -1120
rect 439562 -1176 439618 -1120
rect 439686 -1176 439742 -1120
rect 439314 -1300 439370 -1244
rect 439438 -1300 439494 -1244
rect 439562 -1300 439618 -1244
rect 439686 -1300 439742 -1244
rect 439314 -1424 439370 -1368
rect 439438 -1424 439494 -1368
rect 439562 -1424 439618 -1368
rect 439686 -1424 439742 -1368
rect 439314 -1548 439370 -1492
rect 439438 -1548 439494 -1492
rect 439562 -1548 439618 -1492
rect 439686 -1548 439742 -1492
rect 466314 40294 466370 40350
rect 466438 40294 466494 40350
rect 466562 40294 466618 40350
rect 466686 40294 466742 40350
rect 466314 40170 466370 40226
rect 466438 40170 466494 40226
rect 466562 40170 466618 40226
rect 466686 40170 466742 40226
rect 466314 40046 466370 40102
rect 466438 40046 466494 40102
rect 466562 40046 466618 40102
rect 466686 40046 466742 40102
rect 466314 39922 466370 39978
rect 466438 39922 466494 39978
rect 466562 39922 466618 39978
rect 466686 39922 466742 39978
rect 466314 22294 466370 22350
rect 466438 22294 466494 22350
rect 466562 22294 466618 22350
rect 466686 22294 466742 22350
rect 466314 22170 466370 22226
rect 466438 22170 466494 22226
rect 466562 22170 466618 22226
rect 466686 22170 466742 22226
rect 466314 22046 466370 22102
rect 466438 22046 466494 22102
rect 466562 22046 466618 22102
rect 466686 22046 466742 22102
rect 466314 21922 466370 21978
rect 466438 21922 466494 21978
rect 466562 21922 466618 21978
rect 466686 21922 466742 21978
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 470034 46294 470090 46350
rect 470158 46294 470214 46350
rect 470282 46294 470338 46350
rect 470406 46294 470462 46350
rect 470034 46170 470090 46226
rect 470158 46170 470214 46226
rect 470282 46170 470338 46226
rect 470406 46170 470462 46226
rect 470034 46046 470090 46102
rect 470158 46046 470214 46102
rect 470282 46046 470338 46102
rect 470406 46046 470462 46102
rect 470034 45922 470090 45978
rect 470158 45922 470214 45978
rect 470282 45922 470338 45978
rect 470406 45922 470462 45978
rect 470034 28294 470090 28350
rect 470158 28294 470214 28350
rect 470282 28294 470338 28350
rect 470406 28294 470462 28350
rect 470034 28170 470090 28226
rect 470158 28170 470214 28226
rect 470282 28170 470338 28226
rect 470406 28170 470462 28226
rect 470034 28046 470090 28102
rect 470158 28046 470214 28102
rect 470282 28046 470338 28102
rect 470406 28046 470462 28102
rect 470034 27922 470090 27978
rect 470158 27922 470214 27978
rect 470282 27922 470338 27978
rect 470406 27922 470462 27978
rect 470034 10294 470090 10350
rect 470158 10294 470214 10350
rect 470282 10294 470338 10350
rect 470406 10294 470462 10350
rect 470034 10170 470090 10226
rect 470158 10170 470214 10226
rect 470282 10170 470338 10226
rect 470406 10170 470462 10226
rect 470034 10046 470090 10102
rect 470158 10046 470214 10102
rect 470282 10046 470338 10102
rect 470406 10046 470462 10102
rect 470034 9922 470090 9978
rect 470158 9922 470214 9978
rect 470282 9922 470338 9978
rect 470406 9922 470462 9978
rect 470034 -1176 470090 -1120
rect 470158 -1176 470214 -1120
rect 470282 -1176 470338 -1120
rect 470406 -1176 470462 -1120
rect 470034 -1300 470090 -1244
rect 470158 -1300 470214 -1244
rect 470282 -1300 470338 -1244
rect 470406 -1300 470462 -1244
rect 470034 -1424 470090 -1368
rect 470158 -1424 470214 -1368
rect 470282 -1424 470338 -1368
rect 470406 -1424 470462 -1368
rect 470034 -1548 470090 -1492
rect 470158 -1548 470214 -1492
rect 470282 -1548 470338 -1492
rect 470406 -1548 470462 -1492
rect 497034 40294 497090 40350
rect 497158 40294 497214 40350
rect 497282 40294 497338 40350
rect 497406 40294 497462 40350
rect 497034 40170 497090 40226
rect 497158 40170 497214 40226
rect 497282 40170 497338 40226
rect 497406 40170 497462 40226
rect 497034 40046 497090 40102
rect 497158 40046 497214 40102
rect 497282 40046 497338 40102
rect 497406 40046 497462 40102
rect 497034 39922 497090 39978
rect 497158 39922 497214 39978
rect 497282 39922 497338 39978
rect 497406 39922 497462 39978
rect 497034 22294 497090 22350
rect 497158 22294 497214 22350
rect 497282 22294 497338 22350
rect 497406 22294 497462 22350
rect 497034 22170 497090 22226
rect 497158 22170 497214 22226
rect 497282 22170 497338 22226
rect 497406 22170 497462 22226
rect 497034 22046 497090 22102
rect 497158 22046 497214 22102
rect 497282 22046 497338 22102
rect 497406 22046 497462 22102
rect 497034 21922 497090 21978
rect 497158 21922 497214 21978
rect 497282 21922 497338 21978
rect 497406 21922 497462 21978
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 500754 46294 500810 46350
rect 500878 46294 500934 46350
rect 501002 46294 501058 46350
rect 501126 46294 501182 46350
rect 500754 46170 500810 46226
rect 500878 46170 500934 46226
rect 501002 46170 501058 46226
rect 501126 46170 501182 46226
rect 500754 46046 500810 46102
rect 500878 46046 500934 46102
rect 501002 46046 501058 46102
rect 501126 46046 501182 46102
rect 500754 45922 500810 45978
rect 500878 45922 500934 45978
rect 501002 45922 501058 45978
rect 501126 45922 501182 45978
rect 500754 28294 500810 28350
rect 500878 28294 500934 28350
rect 501002 28294 501058 28350
rect 501126 28294 501182 28350
rect 500754 28170 500810 28226
rect 500878 28170 500934 28226
rect 501002 28170 501058 28226
rect 501126 28170 501182 28226
rect 500754 28046 500810 28102
rect 500878 28046 500934 28102
rect 501002 28046 501058 28102
rect 501126 28046 501182 28102
rect 500754 27922 500810 27978
rect 500878 27922 500934 27978
rect 501002 27922 501058 27978
rect 501126 27922 501182 27978
rect 500754 10294 500810 10350
rect 500878 10294 500934 10350
rect 501002 10294 501058 10350
rect 501126 10294 501182 10350
rect 500754 10170 500810 10226
rect 500878 10170 500934 10226
rect 501002 10170 501058 10226
rect 501126 10170 501182 10226
rect 500754 10046 500810 10102
rect 500878 10046 500934 10102
rect 501002 10046 501058 10102
rect 501126 10046 501182 10102
rect 500754 9922 500810 9978
rect 500878 9922 500934 9978
rect 501002 9922 501058 9978
rect 501126 9922 501182 9978
rect 500754 -1176 500810 -1120
rect 500878 -1176 500934 -1120
rect 501002 -1176 501058 -1120
rect 501126 -1176 501182 -1120
rect 500754 -1300 500810 -1244
rect 500878 -1300 500934 -1244
rect 501002 -1300 501058 -1244
rect 501126 -1300 501182 -1244
rect 500754 -1424 500810 -1368
rect 500878 -1424 500934 -1368
rect 501002 -1424 501058 -1368
rect 501126 -1424 501182 -1368
rect 500754 -1548 500810 -1492
rect 500878 -1548 500934 -1492
rect 501002 -1548 501058 -1492
rect 501126 -1548 501182 -1492
rect 527754 40294 527810 40350
rect 527878 40294 527934 40350
rect 528002 40294 528058 40350
rect 528126 40294 528182 40350
rect 527754 40170 527810 40226
rect 527878 40170 527934 40226
rect 528002 40170 528058 40226
rect 528126 40170 528182 40226
rect 527754 40046 527810 40102
rect 527878 40046 527934 40102
rect 528002 40046 528058 40102
rect 528126 40046 528182 40102
rect 527754 39922 527810 39978
rect 527878 39922 527934 39978
rect 528002 39922 528058 39978
rect 528126 39922 528182 39978
rect 527754 22294 527810 22350
rect 527878 22294 527934 22350
rect 528002 22294 528058 22350
rect 528126 22294 528182 22350
rect 527754 22170 527810 22226
rect 527878 22170 527934 22226
rect 528002 22170 528058 22226
rect 528126 22170 528182 22226
rect 527754 22046 527810 22102
rect 527878 22046 527934 22102
rect 528002 22046 528058 22102
rect 528126 22046 528182 22102
rect 527754 21922 527810 21978
rect 527878 21922 527934 21978
rect 528002 21922 528058 21978
rect 528126 21922 528182 21978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 531474 46294 531530 46350
rect 531598 46294 531654 46350
rect 531722 46294 531778 46350
rect 531846 46294 531902 46350
rect 531474 46170 531530 46226
rect 531598 46170 531654 46226
rect 531722 46170 531778 46226
rect 531846 46170 531902 46226
rect 531474 46046 531530 46102
rect 531598 46046 531654 46102
rect 531722 46046 531778 46102
rect 531846 46046 531902 46102
rect 531474 45922 531530 45978
rect 531598 45922 531654 45978
rect 531722 45922 531778 45978
rect 531846 45922 531902 45978
rect 531474 28294 531530 28350
rect 531598 28294 531654 28350
rect 531722 28294 531778 28350
rect 531846 28294 531902 28350
rect 531474 28170 531530 28226
rect 531598 28170 531654 28226
rect 531722 28170 531778 28226
rect 531846 28170 531902 28226
rect 531474 28046 531530 28102
rect 531598 28046 531654 28102
rect 531722 28046 531778 28102
rect 531846 28046 531902 28102
rect 531474 27922 531530 27978
rect 531598 27922 531654 27978
rect 531722 27922 531778 27978
rect 531846 27922 531902 27978
rect 531474 10294 531530 10350
rect 531598 10294 531654 10350
rect 531722 10294 531778 10350
rect 531846 10294 531902 10350
rect 531474 10170 531530 10226
rect 531598 10170 531654 10226
rect 531722 10170 531778 10226
rect 531846 10170 531902 10226
rect 531474 10046 531530 10102
rect 531598 10046 531654 10102
rect 531722 10046 531778 10102
rect 531846 10046 531902 10102
rect 531474 9922 531530 9978
rect 531598 9922 531654 9978
rect 531722 9922 531778 9978
rect 531846 9922 531902 9978
rect 531474 -1176 531530 -1120
rect 531598 -1176 531654 -1120
rect 531722 -1176 531778 -1120
rect 531846 -1176 531902 -1120
rect 531474 -1300 531530 -1244
rect 531598 -1300 531654 -1244
rect 531722 -1300 531778 -1244
rect 531846 -1300 531902 -1244
rect 531474 -1424 531530 -1368
rect 531598 -1424 531654 -1368
rect 531722 -1424 531778 -1368
rect 531846 -1424 531902 -1368
rect 531474 -1548 531530 -1492
rect 531598 -1548 531654 -1492
rect 531722 -1548 531778 -1492
rect 531846 -1548 531902 -1492
rect 566188 160622 566244 160678
rect 564620 160442 564676 160498
rect 564508 158642 564564 158698
rect 564732 155402 564788 155458
rect 562194 82294 562250 82350
rect 562318 82294 562374 82350
rect 562442 82294 562498 82350
rect 562566 82294 562622 82350
rect 562194 82170 562250 82226
rect 562318 82170 562374 82226
rect 562442 82170 562498 82226
rect 562566 82170 562622 82226
rect 562194 82046 562250 82102
rect 562318 82046 562374 82102
rect 562442 82046 562498 82102
rect 562566 82046 562622 82102
rect 562194 81922 562250 81978
rect 562318 81922 562374 81978
rect 562442 81922 562498 81978
rect 562566 81922 562622 81978
rect 562194 64294 562250 64350
rect 562318 64294 562374 64350
rect 562442 64294 562498 64350
rect 562566 64294 562622 64350
rect 562194 64170 562250 64226
rect 562318 64170 562374 64226
rect 562442 64170 562498 64226
rect 562566 64170 562622 64226
rect 562194 64046 562250 64102
rect 562318 64046 562374 64102
rect 562442 64046 562498 64102
rect 562566 64046 562622 64102
rect 562194 63922 562250 63978
rect 562318 63922 562374 63978
rect 562442 63922 562498 63978
rect 562566 63922 562622 63978
rect 562194 46294 562250 46350
rect 562318 46294 562374 46350
rect 562442 46294 562498 46350
rect 562566 46294 562622 46350
rect 562194 46170 562250 46226
rect 562318 46170 562374 46226
rect 562442 46170 562498 46226
rect 562566 46170 562622 46226
rect 562194 46046 562250 46102
rect 562318 46046 562374 46102
rect 562442 46046 562498 46102
rect 562566 46046 562622 46102
rect 562194 45922 562250 45978
rect 562318 45922 562374 45978
rect 562442 45922 562498 45978
rect 562566 45922 562622 45978
rect 558474 40294 558530 40350
rect 558598 40294 558654 40350
rect 558722 40294 558778 40350
rect 558846 40294 558902 40350
rect 558474 40170 558530 40226
rect 558598 40170 558654 40226
rect 558722 40170 558778 40226
rect 558846 40170 558902 40226
rect 558474 40046 558530 40102
rect 558598 40046 558654 40102
rect 558722 40046 558778 40102
rect 558846 40046 558902 40102
rect 558474 39922 558530 39978
rect 558598 39922 558654 39978
rect 558722 39922 558778 39978
rect 558846 39922 558902 39978
rect 558474 22294 558530 22350
rect 558598 22294 558654 22350
rect 558722 22294 558778 22350
rect 558846 22294 558902 22350
rect 558474 22170 558530 22226
rect 558598 22170 558654 22226
rect 558722 22170 558778 22226
rect 558846 22170 558902 22226
rect 558474 22046 558530 22102
rect 558598 22046 558654 22102
rect 558722 22046 558778 22102
rect 558846 22046 558902 22102
rect 558474 21922 558530 21978
rect 558598 21922 558654 21978
rect 558722 21922 558778 21978
rect 558846 21922 558902 21978
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 562194 28294 562250 28350
rect 562318 28294 562374 28350
rect 562442 28294 562498 28350
rect 562566 28294 562622 28350
rect 562194 28170 562250 28226
rect 562318 28170 562374 28226
rect 562442 28170 562498 28226
rect 562566 28170 562622 28226
rect 562194 28046 562250 28102
rect 562318 28046 562374 28102
rect 562442 28046 562498 28102
rect 562566 28046 562622 28102
rect 562194 27922 562250 27978
rect 562318 27922 562374 27978
rect 562442 27922 562498 27978
rect 562566 27922 562622 27978
rect 573692 401822 573748 401878
rect 575372 401642 575428 401698
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 590492 403982 590548 404038
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 590604 402362 590660 402418
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 581308 395162 581364 395218
rect 579628 393722 579684 393778
rect 577052 393362 577108 393418
rect 562194 10294 562250 10350
rect 562318 10294 562374 10350
rect 562442 10294 562498 10350
rect 562566 10294 562622 10350
rect 562194 10170 562250 10226
rect 562318 10170 562374 10226
rect 562442 10170 562498 10226
rect 562566 10170 562622 10226
rect 562194 10046 562250 10102
rect 562318 10046 562374 10102
rect 562442 10046 562498 10102
rect 562566 10046 562622 10102
rect 562194 9922 562250 9978
rect 562318 9922 562374 9978
rect 562442 9922 562498 9978
rect 562566 9922 562622 9978
rect 582988 394982 583044 395038
rect 585452 393182 585508 393238
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 590492 392102 590548 392158
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 590492 150362 590548 150418
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 562194 -1176 562250 -1120
rect 562318 -1176 562374 -1120
rect 562442 -1176 562498 -1120
rect 562566 -1176 562622 -1120
rect 562194 -1300 562250 -1244
rect 562318 -1300 562374 -1244
rect 562442 -1300 562498 -1244
rect 562566 -1300 562622 -1244
rect 562194 -1424 562250 -1368
rect 562318 -1424 562374 -1368
rect 562442 -1424 562498 -1368
rect 562566 -1424 562622 -1368
rect 562194 -1548 562250 -1492
rect 562318 -1548 562374 -1492
rect 562442 -1548 562498 -1492
rect 562566 -1548 562622 -1492
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 39954 568350
rect 40010 568294 40078 568350
rect 40134 568294 40202 568350
rect 40258 568294 40326 568350
rect 40382 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 101394 568350
rect 101450 568294 101518 568350
rect 101574 568294 101642 568350
rect 101698 568294 101766 568350
rect 101822 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 39954 568226
rect 40010 568170 40078 568226
rect 40134 568170 40202 568226
rect 40258 568170 40326 568226
rect 40382 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 101394 568226
rect 101450 568170 101518 568226
rect 101574 568170 101642 568226
rect 101698 568170 101766 568226
rect 101822 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 39954 568102
rect 40010 568046 40078 568102
rect 40134 568046 40202 568102
rect 40258 568046 40326 568102
rect 40382 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 101394 568102
rect 101450 568046 101518 568102
rect 101574 568046 101642 568102
rect 101698 568046 101766 568102
rect 101822 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 39954 567978
rect 40010 567922 40078 567978
rect 40134 567922 40202 567978
rect 40258 567922 40326 567978
rect 40382 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 101394 567978
rect 101450 567922 101518 567978
rect 101574 567922 101642 567978
rect 101698 567922 101766 567978
rect 101822 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 194518 562350
rect 194574 562294 194642 562350
rect 194698 562294 225238 562350
rect 225294 562294 225362 562350
rect 225418 562294 255958 562350
rect 256014 562294 256082 562350
rect 256138 562294 286678 562350
rect 286734 562294 286802 562350
rect 286858 562294 317398 562350
rect 317454 562294 317522 562350
rect 317578 562294 348118 562350
rect 348174 562294 348242 562350
rect 348298 562294 378838 562350
rect 378894 562294 378962 562350
rect 379018 562294 409558 562350
rect 409614 562294 409682 562350
rect 409738 562294 440278 562350
rect 440334 562294 440402 562350
rect 440458 562294 470998 562350
rect 471054 562294 471122 562350
rect 471178 562294 501718 562350
rect 501774 562294 501842 562350
rect 501898 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 532438 562350
rect 532494 562294 532562 562350
rect 532618 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 194518 562226
rect 194574 562170 194642 562226
rect 194698 562170 225238 562226
rect 225294 562170 225362 562226
rect 225418 562170 255958 562226
rect 256014 562170 256082 562226
rect 256138 562170 286678 562226
rect 286734 562170 286802 562226
rect 286858 562170 317398 562226
rect 317454 562170 317522 562226
rect 317578 562170 348118 562226
rect 348174 562170 348242 562226
rect 348298 562170 378838 562226
rect 378894 562170 378962 562226
rect 379018 562170 409558 562226
rect 409614 562170 409682 562226
rect 409738 562170 440278 562226
rect 440334 562170 440402 562226
rect 440458 562170 470998 562226
rect 471054 562170 471122 562226
rect 471178 562170 501718 562226
rect 501774 562170 501842 562226
rect 501898 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 532438 562226
rect 532494 562170 532562 562226
rect 532618 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 194518 562102
rect 194574 562046 194642 562102
rect 194698 562046 225238 562102
rect 225294 562046 225362 562102
rect 225418 562046 255958 562102
rect 256014 562046 256082 562102
rect 256138 562046 286678 562102
rect 286734 562046 286802 562102
rect 286858 562046 317398 562102
rect 317454 562046 317522 562102
rect 317578 562046 348118 562102
rect 348174 562046 348242 562102
rect 348298 562046 378838 562102
rect 378894 562046 378962 562102
rect 379018 562046 409558 562102
rect 409614 562046 409682 562102
rect 409738 562046 440278 562102
rect 440334 562046 440402 562102
rect 440458 562046 470998 562102
rect 471054 562046 471122 562102
rect 471178 562046 501718 562102
rect 501774 562046 501842 562102
rect 501898 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 532438 562102
rect 532494 562046 532562 562102
rect 532618 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561988 597980 562046
rect -1916 561978 117336 561988
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561932 117336 561978
rect 117392 561932 117460 561988
rect 117516 561932 117584 561988
rect 117640 561932 117708 561988
rect 117764 561932 117832 561988
rect 117888 561932 117956 561988
rect 118012 561932 118080 561988
rect 118136 561932 118204 561988
rect 118260 561932 118328 561988
rect 118384 561932 118452 561988
rect 118508 561932 118576 561988
rect 118632 561932 118700 561988
rect 118756 561932 118824 561988
rect 118880 561932 118948 561988
rect 119004 561932 119072 561988
rect 119128 561932 119196 561988
rect 119252 561932 119320 561988
rect 119376 561932 119444 561988
rect 119500 561932 119568 561988
rect 119624 561932 119692 561988
rect 119748 561932 119816 561988
rect 119872 561932 119940 561988
rect 119996 561932 120064 561988
rect 120120 561932 120188 561988
rect 120244 561932 120312 561988
rect 120368 561932 120436 561988
rect 120492 561932 120560 561988
rect 120616 561932 120684 561988
rect 120740 561932 120808 561988
rect 120864 561932 120932 561988
rect 120988 561932 121056 561988
rect 121112 561932 121180 561988
rect 121236 561932 121304 561988
rect 121360 561932 121428 561988
rect 121484 561932 121552 561988
rect 121608 561932 121676 561988
rect 121732 561932 121800 561988
rect 121856 561932 121924 561988
rect 121980 561932 122048 561988
rect 122104 561932 122172 561988
rect 122228 561932 122296 561988
rect 122352 561932 122420 561988
rect 122476 561932 122544 561988
rect 122600 561932 122668 561988
rect 122724 561932 122792 561988
rect 122848 561932 122916 561988
rect 122972 561932 123040 561988
rect 123096 561932 123164 561988
rect 123220 561932 123288 561988
rect 123344 561932 123412 561988
rect 123468 561932 123536 561988
rect 123592 561932 123660 561988
rect 123716 561932 123784 561988
rect 123840 561932 123908 561988
rect 123964 561932 124032 561988
rect 124088 561932 124156 561988
rect 124212 561932 124280 561988
rect 124336 561932 124404 561988
rect 124460 561932 124528 561988
rect 124584 561978 597980 561988
rect 124584 561932 128394 561978
rect 98102 561922 128394 561932
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 194518 561978
rect 194574 561922 194642 561978
rect 194698 561922 225238 561978
rect 225294 561922 225362 561978
rect 225418 561922 255958 561978
rect 256014 561922 256082 561978
rect 256138 561922 286678 561978
rect 286734 561922 286802 561978
rect 286858 561922 317398 561978
rect 317454 561922 317522 561978
rect 317578 561922 348118 561978
rect 348174 561922 348242 561978
rect 348298 561922 378838 561978
rect 378894 561922 378962 561978
rect 379018 561922 409558 561978
rect 409614 561922 409682 561978
rect 409738 561922 440278 561978
rect 440334 561922 440402 561978
rect 440458 561922 470998 561978
rect 471054 561922 471122 561978
rect 471178 561922 501718 561978
rect 501774 561922 501842 561978
rect 501898 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 532438 561978
rect 532494 561922 532562 561978
rect 532618 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 39954 550350
rect 40010 550294 40078 550350
rect 40134 550294 40202 550350
rect 40258 550294 40326 550350
rect 40382 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 101394 550350
rect 101450 550294 101518 550350
rect 101574 550294 101642 550350
rect 101698 550294 101766 550350
rect 101822 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 162834 550350
rect 162890 550294 162958 550350
rect 163014 550294 163082 550350
rect 163138 550294 163206 550350
rect 163262 550294 209878 550350
rect 209934 550294 210002 550350
rect 210058 550294 240598 550350
rect 240654 550294 240722 550350
rect 240778 550294 271318 550350
rect 271374 550294 271442 550350
rect 271498 550294 302038 550350
rect 302094 550294 302162 550350
rect 302218 550294 332758 550350
rect 332814 550294 332882 550350
rect 332938 550294 363478 550350
rect 363534 550294 363602 550350
rect 363658 550294 394198 550350
rect 394254 550294 394322 550350
rect 394378 550294 424918 550350
rect 424974 550294 425042 550350
rect 425098 550294 455638 550350
rect 455694 550294 455762 550350
rect 455818 550294 486358 550350
rect 486414 550294 486482 550350
rect 486538 550294 517078 550350
rect 517134 550294 517202 550350
rect 517258 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 547798 550350
rect 547854 550294 547922 550350
rect 547978 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 39954 550226
rect 40010 550170 40078 550226
rect 40134 550170 40202 550226
rect 40258 550170 40326 550226
rect 40382 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 101394 550226
rect 101450 550170 101518 550226
rect 101574 550170 101642 550226
rect 101698 550170 101766 550226
rect 101822 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 162834 550226
rect 162890 550170 162958 550226
rect 163014 550170 163082 550226
rect 163138 550170 163206 550226
rect 163262 550170 209878 550226
rect 209934 550170 210002 550226
rect 210058 550170 240598 550226
rect 240654 550170 240722 550226
rect 240778 550170 271318 550226
rect 271374 550170 271442 550226
rect 271498 550170 302038 550226
rect 302094 550170 302162 550226
rect 302218 550170 332758 550226
rect 332814 550170 332882 550226
rect 332938 550170 363478 550226
rect 363534 550170 363602 550226
rect 363658 550170 394198 550226
rect 394254 550170 394322 550226
rect 394378 550170 424918 550226
rect 424974 550170 425042 550226
rect 425098 550170 455638 550226
rect 455694 550170 455762 550226
rect 455818 550170 486358 550226
rect 486414 550170 486482 550226
rect 486538 550170 517078 550226
rect 517134 550170 517202 550226
rect 517258 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 547798 550226
rect 547854 550170 547922 550226
rect 547978 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 39954 550102
rect 40010 550046 40078 550102
rect 40134 550046 40202 550102
rect 40258 550046 40326 550102
rect 40382 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 101394 550102
rect 101450 550046 101518 550102
rect 101574 550046 101642 550102
rect 101698 550046 101766 550102
rect 101822 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 162834 550102
rect 162890 550046 162958 550102
rect 163014 550046 163082 550102
rect 163138 550046 163206 550102
rect 163262 550046 209878 550102
rect 209934 550046 210002 550102
rect 210058 550046 240598 550102
rect 240654 550046 240722 550102
rect 240778 550046 271318 550102
rect 271374 550046 271442 550102
rect 271498 550046 302038 550102
rect 302094 550046 302162 550102
rect 302218 550046 332758 550102
rect 332814 550046 332882 550102
rect 332938 550046 363478 550102
rect 363534 550046 363602 550102
rect 363658 550046 394198 550102
rect 394254 550046 394322 550102
rect 394378 550046 424918 550102
rect 424974 550046 425042 550102
rect 425098 550046 455638 550102
rect 455694 550046 455762 550102
rect 455818 550046 486358 550102
rect 486414 550046 486482 550102
rect 486538 550046 517078 550102
rect 517134 550046 517202 550102
rect 517258 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 547798 550102
rect 547854 550046 547922 550102
rect 547978 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 39954 549978
rect 40010 549922 40078 549978
rect 40134 549922 40202 549978
rect 40258 549922 40326 549978
rect 40382 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 101394 549978
rect 101450 549922 101518 549978
rect 101574 549922 101642 549978
rect 101698 549922 101766 549978
rect 101822 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 162834 549978
rect 162890 549922 162958 549978
rect 163014 549922 163082 549978
rect 163138 549922 163206 549978
rect 163262 549922 209878 549978
rect 209934 549922 210002 549978
rect 210058 549922 240598 549978
rect 240654 549922 240722 549978
rect 240778 549922 271318 549978
rect 271374 549922 271442 549978
rect 271498 549922 302038 549978
rect 302094 549922 302162 549978
rect 302218 549922 332758 549978
rect 332814 549922 332882 549978
rect 332938 549922 363478 549978
rect 363534 549922 363602 549978
rect 363658 549922 394198 549978
rect 394254 549922 394322 549978
rect 394378 549922 424918 549978
rect 424974 549922 425042 549978
rect 425098 549922 455638 549978
rect 455694 549922 455762 549978
rect 455818 549922 486358 549978
rect 486414 549922 486482 549978
rect 486538 549922 517078 549978
rect 517134 549922 517202 549978
rect 517258 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 547798 549978
rect 547854 549922 547922 549978
rect 547978 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 97674 544350
rect 97730 544294 97798 544350
rect 97854 544294 97922 544350
rect 97978 544294 98046 544350
rect 98102 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 194518 544350
rect 194574 544294 194642 544350
rect 194698 544294 225238 544350
rect 225294 544294 225362 544350
rect 225418 544294 255958 544350
rect 256014 544294 256082 544350
rect 256138 544294 286678 544350
rect 286734 544294 286802 544350
rect 286858 544294 317398 544350
rect 317454 544294 317522 544350
rect 317578 544294 348118 544350
rect 348174 544294 348242 544350
rect 348298 544294 378838 544350
rect 378894 544294 378962 544350
rect 379018 544294 409558 544350
rect 409614 544294 409682 544350
rect 409738 544294 440278 544350
rect 440334 544294 440402 544350
rect 440458 544294 470998 544350
rect 471054 544294 471122 544350
rect 471178 544294 501718 544350
rect 501774 544294 501842 544350
rect 501898 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 532438 544350
rect 532494 544294 532562 544350
rect 532618 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 97674 544226
rect 97730 544170 97798 544226
rect 97854 544170 97922 544226
rect 97978 544170 98046 544226
rect 98102 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 194518 544226
rect 194574 544170 194642 544226
rect 194698 544170 225238 544226
rect 225294 544170 225362 544226
rect 225418 544170 255958 544226
rect 256014 544170 256082 544226
rect 256138 544170 286678 544226
rect 286734 544170 286802 544226
rect 286858 544170 317398 544226
rect 317454 544170 317522 544226
rect 317578 544170 348118 544226
rect 348174 544170 348242 544226
rect 348298 544170 378838 544226
rect 378894 544170 378962 544226
rect 379018 544170 409558 544226
rect 409614 544170 409682 544226
rect 409738 544170 440278 544226
rect 440334 544170 440402 544226
rect 440458 544170 470998 544226
rect 471054 544170 471122 544226
rect 471178 544170 501718 544226
rect 501774 544170 501842 544226
rect 501898 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 532438 544226
rect 532494 544170 532562 544226
rect 532618 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 97674 544102
rect 97730 544046 97798 544102
rect 97854 544046 97922 544102
rect 97978 544046 98046 544102
rect 98102 544063 128394 544102
rect 98102 544046 104066 544063
rect -1916 544007 104066 544046
rect 104122 544007 104190 544063
rect 104246 544007 104314 544063
rect 104370 544007 104438 544063
rect 104494 544007 104562 544063
rect 104618 544007 104686 544063
rect 104742 544007 104810 544063
rect 104866 544007 104934 544063
rect 104990 544007 105058 544063
rect 105114 544007 105182 544063
rect 105238 544007 105306 544063
rect 105362 544007 105430 544063
rect 105486 544007 105554 544063
rect 105610 544007 105678 544063
rect 105734 544007 105802 544063
rect 105858 544007 105926 544063
rect 105982 544007 106050 544063
rect 106106 544007 106174 544063
rect 106230 544007 106298 544063
rect 106354 544007 106422 544063
rect 106478 544007 106546 544063
rect 106602 544007 106670 544063
rect 106726 544007 106794 544063
rect 106850 544007 106918 544063
rect 106974 544007 107042 544063
rect 107098 544007 107166 544063
rect 107222 544007 107290 544063
rect 107346 544007 107414 544063
rect 107470 544007 107538 544063
rect 107594 544007 107662 544063
rect 107718 544007 107786 544063
rect 107842 544007 107910 544063
rect 107966 544007 108034 544063
rect 108090 544007 108158 544063
rect 108214 544007 108282 544063
rect 108338 544007 108406 544063
rect 108462 544007 108530 544063
rect 108586 544007 108654 544063
rect 108710 544007 108778 544063
rect 108834 544007 108902 544063
rect 108958 544007 109026 544063
rect 109082 544007 109150 544063
rect 109206 544007 109274 544063
rect 109330 544007 109398 544063
rect 109454 544007 109522 544063
rect 109578 544007 109646 544063
rect 109702 544007 109770 544063
rect 109826 544007 109894 544063
rect 109950 544007 110018 544063
rect 110074 544007 110142 544063
rect 110198 544007 110266 544063
rect 110322 544007 110390 544063
rect 110446 544007 110514 544063
rect 110570 544007 110638 544063
rect 110694 544007 110762 544063
rect 110818 544007 110886 544063
rect 110942 544007 111010 544063
rect 111066 544007 111134 544063
rect 111190 544007 111258 544063
rect 111314 544007 111382 544063
rect 111438 544007 111506 544063
rect 111562 544007 111630 544063
rect 111686 544007 111754 544063
rect 111810 544007 111878 544063
rect 111934 544007 112002 544063
rect 112058 544007 112126 544063
rect 112182 544007 112250 544063
rect 112306 544007 112374 544063
rect 112430 544007 112498 544063
rect 112554 544007 112622 544063
rect 112678 544007 112746 544063
rect 112802 544007 112870 544063
rect 112926 544007 112994 544063
rect 113050 544007 113118 544063
rect 113174 544007 113242 544063
rect 113298 544007 113366 544063
rect 113422 544007 113490 544063
rect 113546 544007 113614 544063
rect 113670 544007 113738 544063
rect 113794 544007 113862 544063
rect 113918 544007 113986 544063
rect 114042 544007 114110 544063
rect 114166 544007 114234 544063
rect 114290 544007 114358 544063
rect 114414 544007 114482 544063
rect 114538 544007 114606 544063
rect 114662 544007 114730 544063
rect 114786 544007 114854 544063
rect 114910 544007 114978 544063
rect 115034 544007 115102 544063
rect 115158 544007 115226 544063
rect 115282 544007 115350 544063
rect 115406 544007 115474 544063
rect 115530 544007 115598 544063
rect 115654 544007 115722 544063
rect 115778 544007 115846 544063
rect 115902 544007 115970 544063
rect 116026 544007 116094 544063
rect 116150 544007 116218 544063
rect 116274 544007 116342 544063
rect 116398 544007 116466 544063
rect 116522 544007 116590 544063
rect 116646 544007 116714 544063
rect 116770 544007 116838 544063
rect 116894 544007 116962 544063
rect 117018 544007 117086 544063
rect 117142 544007 117210 544063
rect 117266 544007 117334 544063
rect 117390 544007 117458 544063
rect 117514 544007 117582 544063
rect 117638 544007 117706 544063
rect 117762 544007 117830 544063
rect 117886 544007 117954 544063
rect 118010 544007 118078 544063
rect 118134 544007 118202 544063
rect 118258 544007 118326 544063
rect 118382 544007 118450 544063
rect 118506 544007 118574 544063
rect 118630 544007 118698 544063
rect 118754 544007 118822 544063
rect 118878 544007 118946 544063
rect 119002 544007 119070 544063
rect 119126 544007 119194 544063
rect 119250 544007 119318 544063
rect 119374 544007 119442 544063
rect 119498 544007 119566 544063
rect 119622 544007 119690 544063
rect 119746 544007 119814 544063
rect 119870 544007 119938 544063
rect 119994 544007 120062 544063
rect 120118 544007 120186 544063
rect 120242 544007 120310 544063
rect 120366 544007 120434 544063
rect 120490 544007 120558 544063
rect 120614 544007 120682 544063
rect 120738 544007 120806 544063
rect 120862 544007 120930 544063
rect 120986 544007 121054 544063
rect 121110 544007 121178 544063
rect 121234 544007 121302 544063
rect 121358 544007 121426 544063
rect 121482 544007 121550 544063
rect 121606 544007 121674 544063
rect 121730 544007 121798 544063
rect 121854 544046 128394 544063
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 194518 544102
rect 194574 544046 194642 544102
rect 194698 544046 225238 544102
rect 225294 544046 225362 544102
rect 225418 544046 255958 544102
rect 256014 544046 256082 544102
rect 256138 544046 286678 544102
rect 286734 544046 286802 544102
rect 286858 544046 317398 544102
rect 317454 544046 317522 544102
rect 317578 544046 348118 544102
rect 348174 544046 348242 544102
rect 348298 544046 378838 544102
rect 378894 544046 378962 544102
rect 379018 544046 409558 544102
rect 409614 544046 409682 544102
rect 409738 544046 440278 544102
rect 440334 544046 440402 544102
rect 440458 544046 470998 544102
rect 471054 544046 471122 544102
rect 471178 544046 501718 544102
rect 501774 544046 501842 544102
rect 501898 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 532438 544102
rect 532494 544046 532562 544102
rect 532618 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect 121854 544007 597980 544046
rect -1916 543978 597980 544007
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 97674 543978
rect 97730 543922 97798 543978
rect 97854 543922 97922 543978
rect 97978 543922 98046 543978
rect 98102 543939 128394 543978
rect 98102 543922 104066 543939
rect -1916 543883 104066 543922
rect 104122 543883 104190 543939
rect 104246 543883 104314 543939
rect 104370 543883 104438 543939
rect 104494 543883 104562 543939
rect 104618 543883 104686 543939
rect 104742 543883 104810 543939
rect 104866 543883 104934 543939
rect 104990 543883 105058 543939
rect 105114 543883 105182 543939
rect 105238 543883 105306 543939
rect 105362 543883 105430 543939
rect 105486 543883 105554 543939
rect 105610 543883 105678 543939
rect 105734 543883 105802 543939
rect 105858 543883 105926 543939
rect 105982 543883 106050 543939
rect 106106 543883 106174 543939
rect 106230 543883 106298 543939
rect 106354 543883 106422 543939
rect 106478 543883 106546 543939
rect 106602 543883 106670 543939
rect 106726 543883 106794 543939
rect 106850 543883 106918 543939
rect 106974 543883 107042 543939
rect 107098 543883 107166 543939
rect 107222 543883 107290 543939
rect 107346 543883 107414 543939
rect 107470 543883 107538 543939
rect 107594 543883 107662 543939
rect 107718 543883 107786 543939
rect 107842 543883 107910 543939
rect 107966 543883 108034 543939
rect 108090 543883 108158 543939
rect 108214 543883 108282 543939
rect 108338 543883 108406 543939
rect 108462 543883 108530 543939
rect 108586 543883 108654 543939
rect 108710 543883 108778 543939
rect 108834 543883 108902 543939
rect 108958 543883 109026 543939
rect 109082 543883 109150 543939
rect 109206 543883 109274 543939
rect 109330 543883 109398 543939
rect 109454 543883 109522 543939
rect 109578 543883 109646 543939
rect 109702 543883 109770 543939
rect 109826 543883 109894 543939
rect 109950 543883 110018 543939
rect 110074 543883 110142 543939
rect 110198 543883 110266 543939
rect 110322 543883 110390 543939
rect 110446 543883 110514 543939
rect 110570 543883 110638 543939
rect 110694 543883 110762 543939
rect 110818 543883 110886 543939
rect 110942 543883 111010 543939
rect 111066 543883 111134 543939
rect 111190 543883 111258 543939
rect 111314 543883 111382 543939
rect 111438 543883 111506 543939
rect 111562 543883 111630 543939
rect 111686 543883 111754 543939
rect 111810 543883 111878 543939
rect 111934 543883 112002 543939
rect 112058 543883 112126 543939
rect 112182 543883 112250 543939
rect 112306 543883 112374 543939
rect 112430 543883 112498 543939
rect 112554 543883 112622 543939
rect 112678 543883 112746 543939
rect 112802 543883 112870 543939
rect 112926 543883 112994 543939
rect 113050 543883 113118 543939
rect 113174 543883 113242 543939
rect 113298 543883 113366 543939
rect 113422 543883 113490 543939
rect 113546 543883 113614 543939
rect 113670 543883 113738 543939
rect 113794 543883 113862 543939
rect 113918 543883 113986 543939
rect 114042 543883 114110 543939
rect 114166 543883 114234 543939
rect 114290 543883 114358 543939
rect 114414 543883 114482 543939
rect 114538 543883 114606 543939
rect 114662 543883 114730 543939
rect 114786 543883 114854 543939
rect 114910 543883 114978 543939
rect 115034 543883 115102 543939
rect 115158 543883 115226 543939
rect 115282 543883 115350 543939
rect 115406 543883 115474 543939
rect 115530 543883 115598 543939
rect 115654 543883 115722 543939
rect 115778 543883 115846 543939
rect 115902 543883 115970 543939
rect 116026 543883 116094 543939
rect 116150 543883 116218 543939
rect 116274 543883 116342 543939
rect 116398 543883 116466 543939
rect 116522 543883 116590 543939
rect 116646 543883 116714 543939
rect 116770 543883 116838 543939
rect 116894 543883 116962 543939
rect 117018 543883 117086 543939
rect 117142 543883 117210 543939
rect 117266 543883 117334 543939
rect 117390 543883 117458 543939
rect 117514 543883 117582 543939
rect 117638 543883 117706 543939
rect 117762 543883 117830 543939
rect 117886 543883 117954 543939
rect 118010 543883 118078 543939
rect 118134 543883 118202 543939
rect 118258 543883 118326 543939
rect 118382 543883 118450 543939
rect 118506 543883 118574 543939
rect 118630 543883 118698 543939
rect 118754 543883 118822 543939
rect 118878 543883 118946 543939
rect 119002 543883 119070 543939
rect 119126 543883 119194 543939
rect 119250 543883 119318 543939
rect 119374 543883 119442 543939
rect 119498 543883 119566 543939
rect 119622 543883 119690 543939
rect 119746 543883 119814 543939
rect 119870 543883 119938 543939
rect 119994 543883 120062 543939
rect 120118 543883 120186 543939
rect 120242 543883 120310 543939
rect 120366 543883 120434 543939
rect 120490 543883 120558 543939
rect 120614 543883 120682 543939
rect 120738 543883 120806 543939
rect 120862 543883 120930 543939
rect 120986 543883 121054 543939
rect 121110 543883 121178 543939
rect 121234 543883 121302 543939
rect 121358 543883 121426 543939
rect 121482 543883 121550 543939
rect 121606 543883 121674 543939
rect 121730 543883 121798 543939
rect 121854 543922 128394 543939
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 194518 543978
rect 194574 543922 194642 543978
rect 194698 543922 225238 543978
rect 225294 543922 225362 543978
rect 225418 543922 255958 543978
rect 256014 543922 256082 543978
rect 256138 543922 286678 543978
rect 286734 543922 286802 543978
rect 286858 543922 317398 543978
rect 317454 543922 317522 543978
rect 317578 543922 348118 543978
rect 348174 543922 348242 543978
rect 348298 543922 378838 543978
rect 378894 543922 378962 543978
rect 379018 543922 409558 543978
rect 409614 543922 409682 543978
rect 409738 543922 440278 543978
rect 440334 543922 440402 543978
rect 440458 543922 470998 543978
rect 471054 543922 471122 543978
rect 471178 543922 501718 543978
rect 501774 543922 501842 543978
rect 501898 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 532438 543978
rect 532494 543922 532562 543978
rect 532618 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect 121854 543883 597980 543922
rect -1916 543826 597980 543883
rect -1916 532388 597980 532446
rect -1916 532350 71876 532388
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 39954 532350
rect 40010 532294 40078 532350
rect 40134 532294 40202 532350
rect 40258 532294 40326 532350
rect 40382 532332 71876 532350
rect 71932 532332 72000 532388
rect 72056 532332 72124 532388
rect 72180 532332 72248 532388
rect 72304 532332 72372 532388
rect 72428 532332 72496 532388
rect 72552 532332 72620 532388
rect 72676 532332 72744 532388
rect 72800 532332 72868 532388
rect 72924 532332 72992 532388
rect 73048 532332 73116 532388
rect 73172 532332 73240 532388
rect 73296 532332 73364 532388
rect 73420 532332 73488 532388
rect 73544 532332 73612 532388
rect 73668 532332 73736 532388
rect 73792 532332 73860 532388
rect 73916 532332 73984 532388
rect 74040 532332 74108 532388
rect 74164 532332 74232 532388
rect 74288 532332 74356 532388
rect 74412 532332 74480 532388
rect 74536 532332 74604 532388
rect 74660 532332 74728 532388
rect 74784 532332 74852 532388
rect 74908 532332 74976 532388
rect 75032 532332 75100 532388
rect 75156 532332 75224 532388
rect 75280 532332 75348 532388
rect 75404 532332 75472 532388
rect 75528 532332 75596 532388
rect 75652 532332 75720 532388
rect 75776 532332 75844 532388
rect 75900 532332 75968 532388
rect 76024 532332 76092 532388
rect 76148 532332 76216 532388
rect 76272 532332 76340 532388
rect 76396 532332 76464 532388
rect 76520 532332 76588 532388
rect 76644 532332 76712 532388
rect 76768 532332 76836 532388
rect 76892 532332 76960 532388
rect 77016 532332 77084 532388
rect 77140 532332 77208 532388
rect 77264 532332 77332 532388
rect 77388 532332 77456 532388
rect 77512 532332 77580 532388
rect 77636 532332 77704 532388
rect 77760 532332 77828 532388
rect 77884 532332 77952 532388
rect 78008 532332 78076 532388
rect 78132 532332 78200 532388
rect 78256 532332 78324 532388
rect 78380 532332 78448 532388
rect 78504 532332 78572 532388
rect 78628 532332 78696 532388
rect 78752 532332 78820 532388
rect 78876 532332 78944 532388
rect 79000 532332 79068 532388
rect 79124 532332 79192 532388
rect 79248 532332 79316 532388
rect 79372 532332 79440 532388
rect 79496 532332 79564 532388
rect 79620 532332 79688 532388
rect 79744 532332 79812 532388
rect 79868 532332 79936 532388
rect 79992 532332 80060 532388
rect 80116 532332 80184 532388
rect 80240 532332 80308 532388
rect 80364 532332 80432 532388
rect 80488 532332 80556 532388
rect 80612 532332 80680 532388
rect 80736 532332 80804 532388
rect 80860 532332 80928 532388
rect 80984 532332 81052 532388
rect 81108 532332 81176 532388
rect 81232 532332 81300 532388
rect 81356 532332 81424 532388
rect 81480 532332 81548 532388
rect 81604 532332 81672 532388
rect 81728 532332 81796 532388
rect 81852 532332 81920 532388
rect 81976 532332 82044 532388
rect 82100 532332 82168 532388
rect 82224 532332 82292 532388
rect 82348 532332 82416 532388
rect 82472 532332 82540 532388
rect 82596 532332 82664 532388
rect 82720 532332 82788 532388
rect 82844 532350 597980 532388
rect 82844 532332 162834 532350
rect 40382 532294 162834 532332
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 209878 532350
rect 209934 532294 210002 532350
rect 210058 532294 240598 532350
rect 240654 532294 240722 532350
rect 240778 532294 271318 532350
rect 271374 532294 271442 532350
rect 271498 532294 302038 532350
rect 302094 532294 302162 532350
rect 302218 532294 332758 532350
rect 332814 532294 332882 532350
rect 332938 532294 363478 532350
rect 363534 532294 363602 532350
rect 363658 532294 394198 532350
rect 394254 532294 394322 532350
rect 394378 532294 424918 532350
rect 424974 532294 425042 532350
rect 425098 532294 455638 532350
rect 455694 532294 455762 532350
rect 455818 532294 486358 532350
rect 486414 532294 486482 532350
rect 486538 532294 517078 532350
rect 517134 532294 517202 532350
rect 517258 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 547798 532350
rect 547854 532294 547922 532350
rect 547978 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 39954 532226
rect 40010 532170 40078 532226
rect 40134 532170 40202 532226
rect 40258 532170 40326 532226
rect 40382 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 209878 532226
rect 209934 532170 210002 532226
rect 210058 532170 240598 532226
rect 240654 532170 240722 532226
rect 240778 532170 271318 532226
rect 271374 532170 271442 532226
rect 271498 532170 302038 532226
rect 302094 532170 302162 532226
rect 302218 532170 332758 532226
rect 332814 532170 332882 532226
rect 332938 532170 363478 532226
rect 363534 532170 363602 532226
rect 363658 532170 394198 532226
rect 394254 532170 394322 532226
rect 394378 532170 424918 532226
rect 424974 532170 425042 532226
rect 425098 532170 455638 532226
rect 455694 532170 455762 532226
rect 455818 532170 486358 532226
rect 486414 532170 486482 532226
rect 486538 532170 517078 532226
rect 517134 532170 517202 532226
rect 517258 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 547798 532226
rect 547854 532170 547922 532226
rect 547978 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 39954 532102
rect 40010 532046 40078 532102
rect 40134 532046 40202 532102
rect 40258 532046 40326 532102
rect 40382 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 209878 532102
rect 209934 532046 210002 532102
rect 210058 532046 240598 532102
rect 240654 532046 240722 532102
rect 240778 532046 271318 532102
rect 271374 532046 271442 532102
rect 271498 532046 302038 532102
rect 302094 532046 302162 532102
rect 302218 532046 332758 532102
rect 332814 532046 332882 532102
rect 332938 532046 363478 532102
rect 363534 532046 363602 532102
rect 363658 532046 394198 532102
rect 394254 532046 394322 532102
rect 394378 532046 424918 532102
rect 424974 532046 425042 532102
rect 425098 532046 455638 532102
rect 455694 532046 455762 532102
rect 455818 532046 486358 532102
rect 486414 532046 486482 532102
rect 486538 532046 517078 532102
rect 517134 532046 517202 532102
rect 517258 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 547798 532102
rect 547854 532046 547922 532102
rect 547978 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 39954 531978
rect 40010 531922 40078 531978
rect 40134 531922 40202 531978
rect 40258 531922 40326 531978
rect 40382 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 209878 531978
rect 209934 531922 210002 531978
rect 210058 531922 240598 531978
rect 240654 531922 240722 531978
rect 240778 531922 271318 531978
rect 271374 531922 271442 531978
rect 271498 531922 302038 531978
rect 302094 531922 302162 531978
rect 302218 531922 332758 531978
rect 332814 531922 332882 531978
rect 332938 531922 363478 531978
rect 363534 531922 363602 531978
rect 363658 531922 394198 531978
rect 394254 531922 394322 531978
rect 394378 531922 424918 531978
rect 424974 531922 425042 531978
rect 425098 531922 455638 531978
rect 455694 531922 455762 531978
rect 455818 531922 486358 531978
rect 486414 531922 486482 531978
rect 486538 531922 517078 531978
rect 517134 531922 517202 531978
rect 517258 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 547798 531978
rect 547854 531922 547922 531978
rect 547978 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 194518 526350
rect 194574 526294 194642 526350
rect 194698 526294 225238 526350
rect 225294 526294 225362 526350
rect 225418 526294 255958 526350
rect 256014 526294 256082 526350
rect 256138 526294 286678 526350
rect 286734 526294 286802 526350
rect 286858 526294 317398 526350
rect 317454 526294 317522 526350
rect 317578 526294 348118 526350
rect 348174 526294 348242 526350
rect 348298 526294 378838 526350
rect 378894 526294 378962 526350
rect 379018 526294 409558 526350
rect 409614 526294 409682 526350
rect 409738 526294 440278 526350
rect 440334 526294 440402 526350
rect 440458 526294 470998 526350
rect 471054 526294 471122 526350
rect 471178 526294 501718 526350
rect 501774 526294 501842 526350
rect 501898 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 532438 526350
rect 532494 526294 532562 526350
rect 532618 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 194518 526226
rect 194574 526170 194642 526226
rect 194698 526170 225238 526226
rect 225294 526170 225362 526226
rect 225418 526170 255958 526226
rect 256014 526170 256082 526226
rect 256138 526170 286678 526226
rect 286734 526170 286802 526226
rect 286858 526170 317398 526226
rect 317454 526170 317522 526226
rect 317578 526170 348118 526226
rect 348174 526170 348242 526226
rect 348298 526170 378838 526226
rect 378894 526170 378962 526226
rect 379018 526170 409558 526226
rect 409614 526170 409682 526226
rect 409738 526170 440278 526226
rect 440334 526170 440402 526226
rect 440458 526170 470998 526226
rect 471054 526170 471122 526226
rect 471178 526170 501718 526226
rect 501774 526170 501842 526226
rect 501898 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 532438 526226
rect 532494 526170 532562 526226
rect 532618 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526148 597980 526170
rect -1916 526102 94310 526148
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526092 94310 526102
rect 94366 526092 94434 526148
rect 94490 526092 94558 526148
rect 94614 526092 94682 526148
rect 94738 526092 94806 526148
rect 94862 526092 94930 526148
rect 94986 526092 95054 526148
rect 95110 526092 95178 526148
rect 95234 526092 95302 526148
rect 95358 526092 95426 526148
rect 95482 526092 95550 526148
rect 95606 526092 95674 526148
rect 95730 526092 95798 526148
rect 95854 526092 95922 526148
rect 95978 526092 96046 526148
rect 96102 526092 96170 526148
rect 96226 526092 96294 526148
rect 96350 526092 96418 526148
rect 96474 526092 96542 526148
rect 96598 526092 96666 526148
rect 96722 526092 96790 526148
rect 96846 526092 96914 526148
rect 96970 526092 97038 526148
rect 97094 526092 97162 526148
rect 97218 526092 97286 526148
rect 97342 526092 97410 526148
rect 97466 526092 97534 526148
rect 97590 526092 97658 526148
rect 97714 526092 97782 526148
rect 97838 526092 97906 526148
rect 97962 526092 98030 526148
rect 98086 526092 98154 526148
rect 98210 526092 98278 526148
rect 98334 526092 98402 526148
rect 98458 526092 98526 526148
rect 98582 526092 98650 526148
rect 98706 526092 98774 526148
rect 98830 526092 98898 526148
rect 98954 526092 99022 526148
rect 99078 526092 99146 526148
rect 99202 526092 99270 526148
rect 99326 526092 99394 526148
rect 99450 526092 99518 526148
rect 99574 526092 99642 526148
rect 99698 526092 99766 526148
rect 99822 526092 99890 526148
rect 99946 526092 100014 526148
rect 100070 526092 100138 526148
rect 100194 526092 100262 526148
rect 100318 526092 100386 526148
rect 100442 526092 100510 526148
rect 100566 526092 100634 526148
rect 100690 526092 100758 526148
rect 100814 526092 100882 526148
rect 100938 526092 101006 526148
rect 101062 526092 101130 526148
rect 101186 526092 101254 526148
rect 101310 526092 101378 526148
rect 101434 526092 101502 526148
rect 101558 526092 101626 526148
rect 101682 526092 101750 526148
rect 101806 526092 101874 526148
rect 101930 526092 101998 526148
rect 102054 526092 102122 526148
rect 102178 526092 102246 526148
rect 102302 526092 102370 526148
rect 102426 526092 102494 526148
rect 102550 526092 102618 526148
rect 102674 526092 102742 526148
rect 102798 526092 102866 526148
rect 102922 526092 102990 526148
rect 103046 526092 103114 526148
rect 103170 526092 103238 526148
rect 103294 526092 103362 526148
rect 103418 526092 103486 526148
rect 103542 526092 103610 526148
rect 103666 526092 103734 526148
rect 103790 526092 103858 526148
rect 103914 526092 103982 526148
rect 104038 526092 104106 526148
rect 104162 526092 104230 526148
rect 104286 526092 104354 526148
rect 104410 526092 104478 526148
rect 104534 526092 104602 526148
rect 104658 526092 104726 526148
rect 104782 526092 104850 526148
rect 104906 526092 104974 526148
rect 105030 526092 105098 526148
rect 105154 526092 105222 526148
rect 105278 526092 105346 526148
rect 105402 526092 105470 526148
rect 105526 526092 105594 526148
rect 105650 526092 105718 526148
rect 105774 526092 105842 526148
rect 105898 526092 105966 526148
rect 106022 526092 106090 526148
rect 106146 526092 106214 526148
rect 106270 526092 106338 526148
rect 106394 526092 106462 526148
rect 106518 526092 106586 526148
rect 106642 526092 106710 526148
rect 106766 526092 106834 526148
rect 106890 526092 106958 526148
rect 107014 526092 107082 526148
rect 107138 526092 107206 526148
rect 107262 526092 107330 526148
rect 107386 526092 107454 526148
rect 107510 526092 107578 526148
rect 107634 526092 107702 526148
rect 107758 526092 107826 526148
rect 107882 526092 107950 526148
rect 108006 526092 108074 526148
rect 108130 526092 108198 526148
rect 108254 526092 108322 526148
rect 108378 526092 108446 526148
rect 108502 526092 108570 526148
rect 108626 526092 108694 526148
rect 108750 526092 108818 526148
rect 108874 526092 108942 526148
rect 108998 526092 109066 526148
rect 109122 526092 109190 526148
rect 109246 526092 109314 526148
rect 109370 526092 109438 526148
rect 109494 526092 109562 526148
rect 109618 526092 109686 526148
rect 109742 526092 109810 526148
rect 109866 526092 109934 526148
rect 109990 526092 110058 526148
rect 110114 526092 110182 526148
rect 110238 526092 110306 526148
rect 110362 526092 110430 526148
rect 110486 526092 110554 526148
rect 110610 526092 110678 526148
rect 110734 526092 110802 526148
rect 110858 526092 110926 526148
rect 110982 526092 111050 526148
rect 111106 526092 111174 526148
rect 111230 526092 111298 526148
rect 111354 526092 111422 526148
rect 111478 526092 111546 526148
rect 111602 526092 111670 526148
rect 111726 526092 111794 526148
rect 111850 526092 111918 526148
rect 111974 526092 112042 526148
rect 112098 526092 112166 526148
rect 112222 526092 112290 526148
rect 112346 526092 112414 526148
rect 112470 526092 112538 526148
rect 112594 526092 112662 526148
rect 112718 526092 112786 526148
rect 112842 526092 112910 526148
rect 112966 526092 113034 526148
rect 113090 526092 113158 526148
rect 113214 526092 113282 526148
rect 113338 526092 113406 526148
rect 113462 526092 113530 526148
rect 113586 526092 113654 526148
rect 113710 526092 113778 526148
rect 113834 526092 113902 526148
rect 113958 526092 114026 526148
rect 114082 526092 114150 526148
rect 114206 526092 114274 526148
rect 114330 526102 597980 526148
rect 114330 526092 159114 526102
rect 36662 526046 159114 526092
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 194518 526102
rect 194574 526046 194642 526102
rect 194698 526046 225238 526102
rect 225294 526046 225362 526102
rect 225418 526046 255958 526102
rect 256014 526046 256082 526102
rect 256138 526046 286678 526102
rect 286734 526046 286802 526102
rect 286858 526046 317398 526102
rect 317454 526046 317522 526102
rect 317578 526046 348118 526102
rect 348174 526046 348242 526102
rect 348298 526046 378838 526102
rect 378894 526046 378962 526102
rect 379018 526046 409558 526102
rect 409614 526046 409682 526102
rect 409738 526046 440278 526102
rect 440334 526046 440402 526102
rect 440458 526046 470998 526102
rect 471054 526046 471122 526102
rect 471178 526046 501718 526102
rect 501774 526046 501842 526102
rect 501898 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 532438 526102
rect 532494 526046 532562 526102
rect 532618 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 194518 525978
rect 194574 525922 194642 525978
rect 194698 525922 225238 525978
rect 225294 525922 225362 525978
rect 225418 525922 255958 525978
rect 256014 525922 256082 525978
rect 256138 525922 286678 525978
rect 286734 525922 286802 525978
rect 286858 525922 317398 525978
rect 317454 525922 317522 525978
rect 317578 525922 348118 525978
rect 348174 525922 348242 525978
rect 348298 525922 378838 525978
rect 378894 525922 378962 525978
rect 379018 525922 409558 525978
rect 409614 525922 409682 525978
rect 409738 525922 440278 525978
rect 440334 525922 440402 525978
rect 440458 525922 470998 525978
rect 471054 525922 471122 525978
rect 471178 525922 501718 525978
rect 501774 525922 501842 525978
rect 501898 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 532438 525978
rect 532494 525922 532562 525978
rect 532618 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 39954 514350
rect 40010 514294 40078 514350
rect 40134 514294 40202 514350
rect 40258 514294 40326 514350
rect 40382 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 209878 514350
rect 209934 514294 210002 514350
rect 210058 514294 240598 514350
rect 240654 514294 240722 514350
rect 240778 514294 271318 514350
rect 271374 514294 271442 514350
rect 271498 514294 302038 514350
rect 302094 514294 302162 514350
rect 302218 514294 332758 514350
rect 332814 514294 332882 514350
rect 332938 514294 363478 514350
rect 363534 514294 363602 514350
rect 363658 514294 394198 514350
rect 394254 514294 394322 514350
rect 394378 514294 424918 514350
rect 424974 514294 425042 514350
rect 425098 514294 455638 514350
rect 455694 514294 455762 514350
rect 455818 514294 486358 514350
rect 486414 514294 486482 514350
rect 486538 514294 517078 514350
rect 517134 514294 517202 514350
rect 517258 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 547798 514350
rect 547854 514294 547922 514350
rect 547978 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 39954 514226
rect 40010 514170 40078 514226
rect 40134 514170 40202 514226
rect 40258 514170 40326 514226
rect 40382 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 209878 514226
rect 209934 514170 210002 514226
rect 210058 514170 240598 514226
rect 240654 514170 240722 514226
rect 240778 514170 271318 514226
rect 271374 514170 271442 514226
rect 271498 514170 302038 514226
rect 302094 514170 302162 514226
rect 302218 514170 332758 514226
rect 332814 514170 332882 514226
rect 332938 514170 363478 514226
rect 363534 514170 363602 514226
rect 363658 514170 394198 514226
rect 394254 514170 394322 514226
rect 394378 514170 424918 514226
rect 424974 514170 425042 514226
rect 425098 514170 455638 514226
rect 455694 514170 455762 514226
rect 455818 514170 486358 514226
rect 486414 514170 486482 514226
rect 486538 514170 517078 514226
rect 517134 514170 517202 514226
rect 517258 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 547798 514226
rect 547854 514170 547922 514226
rect 547978 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514130 597980 514170
rect -1916 514102 60844 514130
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 39954 514102
rect 40010 514046 40078 514102
rect 40134 514046 40202 514102
rect 40258 514046 40326 514102
rect 40382 514074 60844 514102
rect 60900 514074 60968 514130
rect 61024 514074 61092 514130
rect 61148 514074 61216 514130
rect 61272 514074 61340 514130
rect 61396 514074 61464 514130
rect 61520 514074 61588 514130
rect 61644 514074 61712 514130
rect 61768 514074 61836 514130
rect 61892 514074 61960 514130
rect 62016 514074 62084 514130
rect 62140 514074 62208 514130
rect 62264 514074 62332 514130
rect 62388 514074 62456 514130
rect 62512 514074 62580 514130
rect 62636 514074 62704 514130
rect 62760 514074 62828 514130
rect 62884 514074 62952 514130
rect 63008 514074 63076 514130
rect 63132 514074 63200 514130
rect 63256 514074 63324 514130
rect 63380 514074 63448 514130
rect 63504 514074 63572 514130
rect 63628 514074 63696 514130
rect 63752 514074 63820 514130
rect 63876 514074 63944 514130
rect 64000 514074 64068 514130
rect 64124 514074 64192 514130
rect 64248 514074 64316 514130
rect 64372 514074 64440 514130
rect 64496 514074 64564 514130
rect 64620 514074 64688 514130
rect 64744 514074 64812 514130
rect 64868 514074 64936 514130
rect 64992 514074 65060 514130
rect 65116 514074 65184 514130
rect 65240 514074 65308 514130
rect 65364 514074 65432 514130
rect 65488 514074 65556 514130
rect 65612 514074 65680 514130
rect 65736 514074 65804 514130
rect 65860 514074 65928 514130
rect 65984 514074 66052 514130
rect 66108 514074 66176 514130
rect 66232 514074 66300 514130
rect 66356 514102 597980 514130
rect 66356 514074 162834 514102
rect 40382 514046 162834 514074
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 209878 514102
rect 209934 514046 210002 514102
rect 210058 514046 240598 514102
rect 240654 514046 240722 514102
rect 240778 514046 271318 514102
rect 271374 514046 271442 514102
rect 271498 514046 302038 514102
rect 302094 514046 302162 514102
rect 302218 514046 332758 514102
rect 332814 514046 332882 514102
rect 332938 514046 363478 514102
rect 363534 514046 363602 514102
rect 363658 514046 394198 514102
rect 394254 514046 394322 514102
rect 394378 514046 424918 514102
rect 424974 514046 425042 514102
rect 425098 514046 455638 514102
rect 455694 514046 455762 514102
rect 455818 514046 486358 514102
rect 486414 514046 486482 514102
rect 486538 514046 517078 514102
rect 517134 514046 517202 514102
rect 517258 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 547798 514102
rect 547854 514046 547922 514102
rect 547978 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 514006 597980 514046
rect -1916 513978 60844 514006
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 39954 513978
rect 40010 513922 40078 513978
rect 40134 513922 40202 513978
rect 40258 513922 40326 513978
rect 40382 513950 60844 513978
rect 60900 513950 60968 514006
rect 61024 513950 61092 514006
rect 61148 513950 61216 514006
rect 61272 513950 61340 514006
rect 61396 513950 61464 514006
rect 61520 513950 61588 514006
rect 61644 513950 61712 514006
rect 61768 513950 61836 514006
rect 61892 513950 61960 514006
rect 62016 513950 62084 514006
rect 62140 513950 62208 514006
rect 62264 513950 62332 514006
rect 62388 513950 62456 514006
rect 62512 513950 62580 514006
rect 62636 513950 62704 514006
rect 62760 513950 62828 514006
rect 62884 513950 62952 514006
rect 63008 513950 63076 514006
rect 63132 513950 63200 514006
rect 63256 513950 63324 514006
rect 63380 513950 63448 514006
rect 63504 513950 63572 514006
rect 63628 513950 63696 514006
rect 63752 513950 63820 514006
rect 63876 513950 63944 514006
rect 64000 513950 64068 514006
rect 64124 513950 64192 514006
rect 64248 513950 64316 514006
rect 64372 513950 64440 514006
rect 64496 513950 64564 514006
rect 64620 513950 64688 514006
rect 64744 513950 64812 514006
rect 64868 513950 64936 514006
rect 64992 513950 65060 514006
rect 65116 513950 65184 514006
rect 65240 513950 65308 514006
rect 65364 513950 65432 514006
rect 65488 513950 65556 514006
rect 65612 513950 65680 514006
rect 65736 513950 65804 514006
rect 65860 513950 65928 514006
rect 65984 513950 66052 514006
rect 66108 513950 66176 514006
rect 66232 513950 66300 514006
rect 66356 513978 597980 514006
rect 66356 513950 162834 513978
rect 40382 513922 162834 513950
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 209878 513978
rect 209934 513922 210002 513978
rect 210058 513922 240598 513978
rect 240654 513922 240722 513978
rect 240778 513922 271318 513978
rect 271374 513922 271442 513978
rect 271498 513922 302038 513978
rect 302094 513922 302162 513978
rect 302218 513922 332758 513978
rect 332814 513922 332882 513978
rect 332938 513922 363478 513978
rect 363534 513922 363602 513978
rect 363658 513922 394198 513978
rect 394254 513922 394322 513978
rect 394378 513922 424918 513978
rect 424974 513922 425042 513978
rect 425098 513922 455638 513978
rect 455694 513922 455762 513978
rect 455818 513922 486358 513978
rect 486414 513922 486482 513978
rect 486538 513922 517078 513978
rect 517134 513922 517202 513978
rect 517258 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 547798 513978
rect 547854 513922 547922 513978
rect 547978 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508388 597980 508446
rect -1916 508350 87884 508388
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508332 87884 508350
rect 87940 508332 88008 508388
rect 88064 508332 88132 508388
rect 88188 508332 88256 508388
rect 88312 508332 88380 508388
rect 88436 508332 88504 508388
rect 88560 508332 88628 508388
rect 88684 508332 88752 508388
rect 88808 508332 88876 508388
rect 88932 508332 89000 508388
rect 89056 508332 89124 508388
rect 89180 508332 89248 508388
rect 89304 508332 89372 508388
rect 89428 508332 89496 508388
rect 89552 508332 89620 508388
rect 89676 508332 89744 508388
rect 89800 508332 89868 508388
rect 89924 508332 89992 508388
rect 90048 508332 90116 508388
rect 90172 508332 90240 508388
rect 90296 508332 90364 508388
rect 90420 508332 90488 508388
rect 90544 508332 90612 508388
rect 90668 508332 90736 508388
rect 90792 508332 90860 508388
rect 90916 508332 90984 508388
rect 91040 508332 91108 508388
rect 91164 508332 91232 508388
rect 91288 508332 91356 508388
rect 91412 508332 91480 508388
rect 91536 508332 91604 508388
rect 91660 508332 91728 508388
rect 91784 508332 91852 508388
rect 91908 508332 91976 508388
rect 92032 508332 92100 508388
rect 92156 508332 92224 508388
rect 92280 508332 92348 508388
rect 92404 508332 92472 508388
rect 92528 508332 92596 508388
rect 92652 508332 92720 508388
rect 92776 508332 92844 508388
rect 92900 508332 92968 508388
rect 93024 508332 93092 508388
rect 93148 508332 93216 508388
rect 93272 508332 93340 508388
rect 93396 508332 93464 508388
rect 93520 508332 93588 508388
rect 93644 508332 93712 508388
rect 93768 508332 93836 508388
rect 93892 508332 93960 508388
rect 94016 508332 94084 508388
rect 94140 508332 94208 508388
rect 94264 508332 94332 508388
rect 94388 508332 94456 508388
rect 94512 508332 94580 508388
rect 94636 508332 94704 508388
rect 94760 508332 94828 508388
rect 94884 508332 94952 508388
rect 95008 508332 95076 508388
rect 95132 508332 95200 508388
rect 95256 508332 95324 508388
rect 95380 508332 95448 508388
rect 95504 508332 95572 508388
rect 95628 508332 95696 508388
rect 95752 508332 95820 508388
rect 95876 508332 95944 508388
rect 96000 508332 96068 508388
rect 96124 508332 96192 508388
rect 96248 508332 96316 508388
rect 96372 508332 96440 508388
rect 96496 508332 96564 508388
rect 96620 508332 96688 508388
rect 96744 508332 96812 508388
rect 96868 508332 96936 508388
rect 96992 508332 97060 508388
rect 97116 508332 97184 508388
rect 97240 508332 97308 508388
rect 97364 508332 97432 508388
rect 97488 508332 97556 508388
rect 97612 508332 97680 508388
rect 97736 508332 97804 508388
rect 97860 508332 97928 508388
rect 97984 508332 98052 508388
rect 98108 508332 98176 508388
rect 98232 508332 98300 508388
rect 98356 508350 597980 508388
rect 98356 508332 159114 508350
rect 36662 508294 159114 508332
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 194518 508350
rect 194574 508294 194642 508350
rect 194698 508294 225238 508350
rect 225294 508294 225362 508350
rect 225418 508294 255958 508350
rect 256014 508294 256082 508350
rect 256138 508294 286678 508350
rect 286734 508294 286802 508350
rect 286858 508294 317398 508350
rect 317454 508294 317522 508350
rect 317578 508294 348118 508350
rect 348174 508294 348242 508350
rect 348298 508294 378838 508350
rect 378894 508294 378962 508350
rect 379018 508294 409558 508350
rect 409614 508294 409682 508350
rect 409738 508294 440278 508350
rect 440334 508294 440402 508350
rect 440458 508294 470998 508350
rect 471054 508294 471122 508350
rect 471178 508294 501718 508350
rect 501774 508294 501842 508350
rect 501898 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 532438 508350
rect 532494 508294 532562 508350
rect 532618 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 194518 508226
rect 194574 508170 194642 508226
rect 194698 508170 225238 508226
rect 225294 508170 225362 508226
rect 225418 508170 255958 508226
rect 256014 508170 256082 508226
rect 256138 508170 286678 508226
rect 286734 508170 286802 508226
rect 286858 508170 317398 508226
rect 317454 508170 317522 508226
rect 317578 508170 348118 508226
rect 348174 508170 348242 508226
rect 348298 508170 378838 508226
rect 378894 508170 378962 508226
rect 379018 508170 409558 508226
rect 409614 508170 409682 508226
rect 409738 508170 440278 508226
rect 440334 508170 440402 508226
rect 440458 508170 470998 508226
rect 471054 508170 471122 508226
rect 471178 508170 501718 508226
rect 501774 508170 501842 508226
rect 501898 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 532438 508226
rect 532494 508170 532562 508226
rect 532618 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508068 159114 508102
rect 36662 508046 87724 508068
rect -1916 508012 87724 508046
rect 87780 508012 87848 508068
rect 87904 508012 87972 508068
rect 88028 508012 88096 508068
rect 88152 508012 88220 508068
rect 88276 508012 88344 508068
rect 88400 508012 88468 508068
rect 88524 508012 88592 508068
rect 88648 508012 88716 508068
rect 88772 508012 88840 508068
rect 88896 508012 88964 508068
rect 89020 508012 89088 508068
rect 89144 508012 89212 508068
rect 89268 508012 89336 508068
rect 89392 508012 89460 508068
rect 89516 508012 89584 508068
rect 89640 508012 89708 508068
rect 89764 508012 89832 508068
rect 89888 508012 89956 508068
rect 90012 508012 90080 508068
rect 90136 508012 90204 508068
rect 90260 508012 90328 508068
rect 90384 508012 90452 508068
rect 90508 508012 90576 508068
rect 90632 508012 90700 508068
rect 90756 508012 90824 508068
rect 90880 508012 90948 508068
rect 91004 508012 91072 508068
rect 91128 508012 91196 508068
rect 91252 508012 91320 508068
rect 91376 508012 91444 508068
rect 91500 508012 91568 508068
rect 91624 508012 91692 508068
rect 91748 508012 91816 508068
rect 91872 508012 91940 508068
rect 91996 508012 92064 508068
rect 92120 508012 92188 508068
rect 92244 508012 92312 508068
rect 92368 508012 92436 508068
rect 92492 508012 92560 508068
rect 92616 508012 92684 508068
rect 92740 508012 92808 508068
rect 92864 508012 92932 508068
rect 92988 508012 93056 508068
rect 93112 508012 93180 508068
rect 93236 508012 93304 508068
rect 93360 508012 93428 508068
rect 93484 508012 93552 508068
rect 93608 508012 93676 508068
rect 93732 508012 93800 508068
rect 93856 508012 93924 508068
rect 93980 508012 94048 508068
rect 94104 508012 94172 508068
rect 94228 508012 94296 508068
rect 94352 508012 94420 508068
rect 94476 508012 94544 508068
rect 94600 508012 94668 508068
rect 94724 508012 94792 508068
rect 94848 508012 94916 508068
rect 94972 508012 95040 508068
rect 95096 508012 95164 508068
rect 95220 508012 95288 508068
rect 95344 508012 95412 508068
rect 95468 508012 95536 508068
rect 95592 508012 95660 508068
rect 95716 508012 95784 508068
rect 95840 508012 95908 508068
rect 95964 508012 96032 508068
rect 96088 508012 96156 508068
rect 96212 508012 96280 508068
rect 96336 508012 96404 508068
rect 96460 508012 96528 508068
rect 96584 508012 96652 508068
rect 96708 508012 96776 508068
rect 96832 508012 96900 508068
rect 96956 508012 97024 508068
rect 97080 508012 97148 508068
rect 97204 508012 97272 508068
rect 97328 508012 97396 508068
rect 97452 508012 97520 508068
rect 97576 508012 97644 508068
rect 97700 508012 97768 508068
rect 97824 508012 97892 508068
rect 97948 508012 98016 508068
rect 98072 508012 98140 508068
rect 98196 508046 159114 508068
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 194518 508102
rect 194574 508046 194642 508102
rect 194698 508046 225238 508102
rect 225294 508046 225362 508102
rect 225418 508046 255958 508102
rect 256014 508046 256082 508102
rect 256138 508046 286678 508102
rect 286734 508046 286802 508102
rect 286858 508046 317398 508102
rect 317454 508046 317522 508102
rect 317578 508046 348118 508102
rect 348174 508046 348242 508102
rect 348298 508046 378838 508102
rect 378894 508046 378962 508102
rect 379018 508046 409558 508102
rect 409614 508046 409682 508102
rect 409738 508046 440278 508102
rect 440334 508046 440402 508102
rect 440458 508046 470998 508102
rect 471054 508046 471122 508102
rect 471178 508046 501718 508102
rect 501774 508046 501842 508102
rect 501898 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 532438 508102
rect 532494 508046 532562 508102
rect 532618 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect 98196 508012 597980 508046
rect -1916 507978 597980 508012
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 194518 507978
rect 194574 507922 194642 507978
rect 194698 507922 225238 507978
rect 225294 507922 225362 507978
rect 225418 507922 255958 507978
rect 256014 507922 256082 507978
rect 256138 507922 286678 507978
rect 286734 507922 286802 507978
rect 286858 507922 317398 507978
rect 317454 507922 317522 507978
rect 317578 507922 348118 507978
rect 348174 507922 348242 507978
rect 348298 507922 378838 507978
rect 378894 507922 378962 507978
rect 379018 507922 409558 507978
rect 409614 507922 409682 507978
rect 409738 507922 440278 507978
rect 440334 507922 440402 507978
rect 440458 507922 470998 507978
rect 471054 507922 471122 507978
rect 471178 507922 501718 507978
rect 501774 507922 501842 507978
rect 501898 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 532438 507978
rect 532494 507922 532562 507978
rect 532618 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496388 597980 496446
rect -1916 496350 61956 496388
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 39954 496350
rect 40010 496294 40078 496350
rect 40134 496294 40202 496350
rect 40258 496294 40326 496350
rect 40382 496332 61956 496350
rect 62012 496332 62080 496388
rect 62136 496332 62204 496388
rect 62260 496332 62328 496388
rect 62384 496332 62452 496388
rect 62508 496332 62576 496388
rect 62632 496332 62700 496388
rect 62756 496332 62824 496388
rect 62880 496332 62948 496388
rect 63004 496332 63072 496388
rect 63128 496332 63196 496388
rect 63252 496332 63320 496388
rect 63376 496332 63444 496388
rect 63500 496332 63568 496388
rect 63624 496332 63692 496388
rect 63748 496332 63816 496388
rect 63872 496332 63940 496388
rect 63996 496332 64064 496388
rect 64120 496332 64188 496388
rect 64244 496332 64312 496388
rect 64368 496332 64436 496388
rect 64492 496332 64560 496388
rect 64616 496332 64684 496388
rect 64740 496332 64808 496388
rect 64864 496332 64932 496388
rect 64988 496332 65056 496388
rect 65112 496332 65180 496388
rect 65236 496332 65304 496388
rect 65360 496332 65428 496388
rect 65484 496332 65552 496388
rect 65608 496332 65676 496388
rect 65732 496332 65800 496388
rect 65856 496332 65924 496388
rect 65980 496332 66048 496388
rect 66104 496332 66172 496388
rect 66228 496332 66296 496388
rect 66352 496332 66420 496388
rect 66476 496332 66544 496388
rect 66600 496332 66668 496388
rect 66724 496332 66792 496388
rect 66848 496332 66916 496388
rect 66972 496332 67040 496388
rect 67096 496332 67164 496388
rect 67220 496332 67288 496388
rect 67344 496332 67412 496388
rect 67468 496332 67536 496388
rect 67592 496332 67660 496388
rect 67716 496332 67784 496388
rect 67840 496332 67908 496388
rect 67964 496350 597980 496388
rect 67964 496332 162834 496350
rect 40382 496294 162834 496332
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 209878 496350
rect 209934 496294 210002 496350
rect 210058 496294 240598 496350
rect 240654 496294 240722 496350
rect 240778 496294 271318 496350
rect 271374 496294 271442 496350
rect 271498 496294 302038 496350
rect 302094 496294 302162 496350
rect 302218 496294 332758 496350
rect 332814 496294 332882 496350
rect 332938 496294 363478 496350
rect 363534 496294 363602 496350
rect 363658 496294 394198 496350
rect 394254 496294 394322 496350
rect 394378 496294 424918 496350
rect 424974 496294 425042 496350
rect 425098 496294 455638 496350
rect 455694 496294 455762 496350
rect 455818 496294 486358 496350
rect 486414 496294 486482 496350
rect 486538 496294 517078 496350
rect 517134 496294 517202 496350
rect 517258 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 547798 496350
rect 547854 496294 547922 496350
rect 547978 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 39954 496226
rect 40010 496170 40078 496226
rect 40134 496170 40202 496226
rect 40258 496170 40326 496226
rect 40382 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 209878 496226
rect 209934 496170 210002 496226
rect 210058 496170 240598 496226
rect 240654 496170 240722 496226
rect 240778 496170 271318 496226
rect 271374 496170 271442 496226
rect 271498 496170 302038 496226
rect 302094 496170 302162 496226
rect 302218 496170 332758 496226
rect 332814 496170 332882 496226
rect 332938 496170 363478 496226
rect 363534 496170 363602 496226
rect 363658 496170 394198 496226
rect 394254 496170 394322 496226
rect 394378 496170 424918 496226
rect 424974 496170 425042 496226
rect 425098 496170 455638 496226
rect 455694 496170 455762 496226
rect 455818 496170 486358 496226
rect 486414 496170 486482 496226
rect 486538 496170 517078 496226
rect 517134 496170 517202 496226
rect 517258 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 547798 496226
rect 547854 496170 547922 496226
rect 547978 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 39954 496102
rect 40010 496046 40078 496102
rect 40134 496046 40202 496102
rect 40258 496046 40326 496102
rect 40382 496063 162834 496102
rect 40382 496046 62116 496063
rect -1916 496007 62116 496046
rect 62172 496007 62240 496063
rect 62296 496007 62364 496063
rect 62420 496007 62488 496063
rect 62544 496007 62612 496063
rect 62668 496007 62736 496063
rect 62792 496007 62860 496063
rect 62916 496007 62984 496063
rect 63040 496007 63108 496063
rect 63164 496007 63232 496063
rect 63288 496007 63356 496063
rect 63412 496007 63480 496063
rect 63536 496007 63604 496063
rect 63660 496007 63728 496063
rect 63784 496007 63852 496063
rect 63908 496007 63976 496063
rect 64032 496007 64100 496063
rect 64156 496007 64224 496063
rect 64280 496007 64348 496063
rect 64404 496007 64472 496063
rect 64528 496007 64596 496063
rect 64652 496007 64720 496063
rect 64776 496007 64844 496063
rect 64900 496007 64968 496063
rect 65024 496007 65092 496063
rect 65148 496007 65216 496063
rect 65272 496007 65340 496063
rect 65396 496007 65464 496063
rect 65520 496007 65588 496063
rect 65644 496007 65712 496063
rect 65768 496007 65836 496063
rect 65892 496007 65960 496063
rect 66016 496007 66084 496063
rect 66140 496007 66208 496063
rect 66264 496007 66332 496063
rect 66388 496007 66456 496063
rect 66512 496007 66580 496063
rect 66636 496007 66704 496063
rect 66760 496007 66828 496063
rect 66884 496007 66952 496063
rect 67008 496007 67076 496063
rect 67132 496007 67200 496063
rect 67256 496007 67324 496063
rect 67380 496007 67448 496063
rect 67504 496007 67572 496063
rect 67628 496007 67696 496063
rect 67752 496007 67820 496063
rect 67876 496007 67944 496063
rect 68000 496007 68068 496063
rect 68124 496046 162834 496063
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 209878 496102
rect 209934 496046 210002 496102
rect 210058 496046 240598 496102
rect 240654 496046 240722 496102
rect 240778 496046 271318 496102
rect 271374 496046 271442 496102
rect 271498 496046 302038 496102
rect 302094 496046 302162 496102
rect 302218 496046 332758 496102
rect 332814 496046 332882 496102
rect 332938 496046 363478 496102
rect 363534 496046 363602 496102
rect 363658 496046 394198 496102
rect 394254 496046 394322 496102
rect 394378 496046 424918 496102
rect 424974 496046 425042 496102
rect 425098 496046 455638 496102
rect 455694 496046 455762 496102
rect 455818 496046 486358 496102
rect 486414 496046 486482 496102
rect 486538 496046 517078 496102
rect 517134 496046 517202 496102
rect 517258 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 547798 496102
rect 547854 496046 547922 496102
rect 547978 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 68124 496007 597980 496046
rect -1916 495978 597980 496007
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 39954 495978
rect 40010 495922 40078 495978
rect 40134 495922 40202 495978
rect 40258 495922 40326 495978
rect 40382 495939 162834 495978
rect 40382 495922 62116 495939
rect -1916 495883 62116 495922
rect 62172 495883 62240 495939
rect 62296 495883 62364 495939
rect 62420 495883 62488 495939
rect 62544 495883 62612 495939
rect 62668 495883 62736 495939
rect 62792 495883 62860 495939
rect 62916 495883 62984 495939
rect 63040 495883 63108 495939
rect 63164 495883 63232 495939
rect 63288 495883 63356 495939
rect 63412 495883 63480 495939
rect 63536 495883 63604 495939
rect 63660 495883 63728 495939
rect 63784 495883 63852 495939
rect 63908 495883 63976 495939
rect 64032 495883 64100 495939
rect 64156 495883 64224 495939
rect 64280 495883 64348 495939
rect 64404 495883 64472 495939
rect 64528 495883 64596 495939
rect 64652 495883 64720 495939
rect 64776 495883 64844 495939
rect 64900 495883 64968 495939
rect 65024 495883 65092 495939
rect 65148 495883 65216 495939
rect 65272 495883 65340 495939
rect 65396 495883 65464 495939
rect 65520 495883 65588 495939
rect 65644 495883 65712 495939
rect 65768 495883 65836 495939
rect 65892 495883 65960 495939
rect 66016 495883 66084 495939
rect 66140 495883 66208 495939
rect 66264 495883 66332 495939
rect 66388 495883 66456 495939
rect 66512 495883 66580 495939
rect 66636 495883 66704 495939
rect 66760 495883 66828 495939
rect 66884 495883 66952 495939
rect 67008 495883 67076 495939
rect 67132 495883 67200 495939
rect 67256 495883 67324 495939
rect 67380 495883 67448 495939
rect 67504 495883 67572 495939
rect 67628 495883 67696 495939
rect 67752 495883 67820 495939
rect 67876 495883 67944 495939
rect 68000 495883 68068 495939
rect 68124 495922 162834 495939
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 209878 495978
rect 209934 495922 210002 495978
rect 210058 495922 240598 495978
rect 240654 495922 240722 495978
rect 240778 495922 271318 495978
rect 271374 495922 271442 495978
rect 271498 495922 302038 495978
rect 302094 495922 302162 495978
rect 302218 495922 332758 495978
rect 332814 495922 332882 495978
rect 332938 495922 363478 495978
rect 363534 495922 363602 495978
rect 363658 495922 394198 495978
rect 394254 495922 394322 495978
rect 394378 495922 424918 495978
rect 424974 495922 425042 495978
rect 425098 495922 455638 495978
rect 455694 495922 455762 495978
rect 455818 495922 486358 495978
rect 486414 495922 486482 495978
rect 486538 495922 517078 495978
rect 517134 495922 517202 495978
rect 517258 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 547798 495978
rect 547854 495922 547922 495978
rect 547978 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 68124 495883 597980 495922
rect -1916 495826 597980 495883
rect -1916 490413 597980 490446
rect -1916 490357 82894 490413
rect 82950 490357 83018 490413
rect 83074 490357 83142 490413
rect 83198 490357 83266 490413
rect 83322 490357 83390 490413
rect 83446 490357 83514 490413
rect 83570 490357 83638 490413
rect 83694 490357 83762 490413
rect 83818 490357 83886 490413
rect 83942 490357 84010 490413
rect 84066 490357 84134 490413
rect 84190 490357 84258 490413
rect 84314 490357 84382 490413
rect 84438 490357 84506 490413
rect 84562 490357 84630 490413
rect 84686 490357 84754 490413
rect 84810 490357 84878 490413
rect 84934 490357 85002 490413
rect 85058 490357 85126 490413
rect 85182 490357 85250 490413
rect 85306 490357 85374 490413
rect 85430 490357 85498 490413
rect 85554 490357 85622 490413
rect 85678 490357 85746 490413
rect 85802 490357 85870 490413
rect 85926 490357 85994 490413
rect 86050 490357 86118 490413
rect 86174 490357 86242 490413
rect 86298 490357 86366 490413
rect 86422 490357 86490 490413
rect 86546 490357 597980 490413
rect -1916 490350 597980 490357
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 194518 490350
rect 194574 490294 194642 490350
rect 194698 490294 225238 490350
rect 225294 490294 225362 490350
rect 225418 490294 255958 490350
rect 256014 490294 256082 490350
rect 256138 490294 286678 490350
rect 286734 490294 286802 490350
rect 286858 490294 317398 490350
rect 317454 490294 317522 490350
rect 317578 490294 348118 490350
rect 348174 490294 348242 490350
rect 348298 490294 378838 490350
rect 378894 490294 378962 490350
rect 379018 490294 409558 490350
rect 409614 490294 409682 490350
rect 409738 490294 440278 490350
rect 440334 490294 440402 490350
rect 440458 490294 470998 490350
rect 471054 490294 471122 490350
rect 471178 490294 501718 490350
rect 501774 490294 501842 490350
rect 501898 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 532438 490350
rect 532494 490294 532562 490350
rect 532618 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490289 597980 490294
rect -1916 490233 82894 490289
rect 82950 490233 83018 490289
rect 83074 490233 83142 490289
rect 83198 490233 83266 490289
rect 83322 490233 83390 490289
rect 83446 490233 83514 490289
rect 83570 490233 83638 490289
rect 83694 490233 83762 490289
rect 83818 490233 83886 490289
rect 83942 490233 84010 490289
rect 84066 490233 84134 490289
rect 84190 490233 84258 490289
rect 84314 490233 84382 490289
rect 84438 490233 84506 490289
rect 84562 490233 84630 490289
rect 84686 490233 84754 490289
rect 84810 490233 84878 490289
rect 84934 490233 85002 490289
rect 85058 490233 85126 490289
rect 85182 490233 85250 490289
rect 85306 490233 85374 490289
rect 85430 490233 85498 490289
rect 85554 490233 85622 490289
rect 85678 490233 85746 490289
rect 85802 490233 85870 490289
rect 85926 490233 85994 490289
rect 86050 490233 86118 490289
rect 86174 490233 86242 490289
rect 86298 490233 86366 490289
rect 86422 490233 86490 490289
rect 86546 490233 597980 490289
rect -1916 490226 597980 490233
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 194518 490226
rect 194574 490170 194642 490226
rect 194698 490170 225238 490226
rect 225294 490170 225362 490226
rect 225418 490170 255958 490226
rect 256014 490170 256082 490226
rect 256138 490170 286678 490226
rect 286734 490170 286802 490226
rect 286858 490170 317398 490226
rect 317454 490170 317522 490226
rect 317578 490170 348118 490226
rect 348174 490170 348242 490226
rect 348298 490170 378838 490226
rect 378894 490170 378962 490226
rect 379018 490170 409558 490226
rect 409614 490170 409682 490226
rect 409738 490170 440278 490226
rect 440334 490170 440402 490226
rect 440458 490170 470998 490226
rect 471054 490170 471122 490226
rect 471178 490170 501718 490226
rect 501774 490170 501842 490226
rect 501898 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 532438 490226
rect 532494 490170 532562 490226
rect 532618 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 194518 490102
rect 194574 490046 194642 490102
rect 194698 490046 225238 490102
rect 225294 490046 225362 490102
rect 225418 490046 255958 490102
rect 256014 490046 256082 490102
rect 256138 490046 286678 490102
rect 286734 490046 286802 490102
rect 286858 490046 317398 490102
rect 317454 490046 317522 490102
rect 317578 490046 348118 490102
rect 348174 490046 348242 490102
rect 348298 490046 378838 490102
rect 378894 490046 378962 490102
rect 379018 490046 409558 490102
rect 409614 490046 409682 490102
rect 409738 490046 440278 490102
rect 440334 490046 440402 490102
rect 440458 490046 470998 490102
rect 471054 490046 471122 490102
rect 471178 490046 501718 490102
rect 501774 490046 501842 490102
rect 501898 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 532438 490102
rect 532494 490046 532562 490102
rect 532618 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489988 597980 490046
rect -1916 489978 82734 489988
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489932 82734 489978
rect 82790 489932 82858 489988
rect 82914 489932 82982 489988
rect 83038 489932 83106 489988
rect 83162 489932 83230 489988
rect 83286 489932 83354 489988
rect 83410 489932 83478 489988
rect 83534 489932 83602 489988
rect 83658 489932 83726 489988
rect 83782 489932 83850 489988
rect 83906 489932 83974 489988
rect 84030 489932 84098 489988
rect 84154 489932 84222 489988
rect 84278 489932 84346 489988
rect 84402 489932 84470 489988
rect 84526 489932 84594 489988
rect 84650 489932 84718 489988
rect 84774 489932 84842 489988
rect 84898 489932 84966 489988
rect 85022 489932 85090 489988
rect 85146 489932 85214 489988
rect 85270 489932 85338 489988
rect 85394 489932 85462 489988
rect 85518 489932 85586 489988
rect 85642 489932 85710 489988
rect 85766 489932 85834 489988
rect 85890 489932 85958 489988
rect 86014 489932 86082 489988
rect 86138 489932 86206 489988
rect 86262 489932 86330 489988
rect 86386 489978 597980 489988
rect 86386 489932 128394 489978
rect 36662 489922 128394 489932
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 194518 489978
rect 194574 489922 194642 489978
rect 194698 489922 225238 489978
rect 225294 489922 225362 489978
rect 225418 489922 255958 489978
rect 256014 489922 256082 489978
rect 256138 489922 286678 489978
rect 286734 489922 286802 489978
rect 286858 489922 317398 489978
rect 317454 489922 317522 489978
rect 317578 489922 348118 489978
rect 348174 489922 348242 489978
rect 348298 489922 378838 489978
rect 378894 489922 378962 489978
rect 379018 489922 409558 489978
rect 409614 489922 409682 489978
rect 409738 489922 440278 489978
rect 440334 489922 440402 489978
rect 440458 489922 470998 489978
rect 471054 489922 471122 489978
rect 471178 489922 501718 489978
rect 501774 489922 501842 489978
rect 501898 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 532438 489978
rect 532494 489922 532562 489978
rect 532618 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 39954 478350
rect 40010 478294 40078 478350
rect 40134 478294 40202 478350
rect 40258 478294 40326 478350
rect 40382 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478308 132114 478350
rect 71102 478294 77956 478308
rect -1916 478252 77956 478294
rect 78012 478252 78080 478308
rect 78136 478252 78204 478308
rect 78260 478252 78328 478308
rect 78384 478252 78452 478308
rect 78508 478252 78576 478308
rect 78632 478252 78700 478308
rect 78756 478252 78824 478308
rect 78880 478252 78948 478308
rect 79004 478294 132114 478308
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 209878 478350
rect 209934 478294 210002 478350
rect 210058 478294 240598 478350
rect 240654 478294 240722 478350
rect 240778 478294 271318 478350
rect 271374 478294 271442 478350
rect 271498 478294 302038 478350
rect 302094 478294 302162 478350
rect 302218 478294 332758 478350
rect 332814 478294 332882 478350
rect 332938 478294 363478 478350
rect 363534 478294 363602 478350
rect 363658 478294 394198 478350
rect 394254 478294 394322 478350
rect 394378 478294 424918 478350
rect 424974 478294 425042 478350
rect 425098 478294 455638 478350
rect 455694 478294 455762 478350
rect 455818 478294 486358 478350
rect 486414 478294 486482 478350
rect 486538 478294 517078 478350
rect 517134 478294 517202 478350
rect 517258 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 547798 478350
rect 547854 478294 547922 478350
rect 547978 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 79004 478252 597980 478294
rect -1916 478226 597980 478252
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 39954 478226
rect 40010 478170 40078 478226
rect 40134 478170 40202 478226
rect 40258 478170 40326 478226
rect 40382 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 209878 478226
rect 209934 478170 210002 478226
rect 210058 478170 240598 478226
rect 240654 478170 240722 478226
rect 240778 478170 271318 478226
rect 271374 478170 271442 478226
rect 271498 478170 302038 478226
rect 302094 478170 302162 478226
rect 302218 478170 332758 478226
rect 332814 478170 332882 478226
rect 332938 478170 363478 478226
rect 363534 478170 363602 478226
rect 363658 478170 394198 478226
rect 394254 478170 394322 478226
rect 394378 478170 424918 478226
rect 424974 478170 425042 478226
rect 425098 478170 455638 478226
rect 455694 478170 455762 478226
rect 455818 478170 486358 478226
rect 486414 478170 486482 478226
rect 486538 478170 517078 478226
rect 517134 478170 517202 478226
rect 517258 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 547798 478226
rect 547854 478170 547922 478226
rect 547978 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 39954 478102
rect 40010 478046 40078 478102
rect 40134 478046 40202 478102
rect 40258 478046 40326 478102
rect 40382 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 209878 478102
rect 209934 478046 210002 478102
rect 210058 478046 240598 478102
rect 240654 478046 240722 478102
rect 240778 478046 271318 478102
rect 271374 478046 271442 478102
rect 271498 478046 302038 478102
rect 302094 478046 302162 478102
rect 302218 478046 332758 478102
rect 332814 478046 332882 478102
rect 332938 478046 363478 478102
rect 363534 478046 363602 478102
rect 363658 478046 394198 478102
rect 394254 478046 394322 478102
rect 394378 478046 424918 478102
rect 424974 478046 425042 478102
rect 425098 478046 455638 478102
rect 455694 478046 455762 478102
rect 455818 478046 486358 478102
rect 486414 478046 486482 478102
rect 486538 478046 517078 478102
rect 517134 478046 517202 478102
rect 517258 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 547798 478102
rect 547854 478046 547922 478102
rect 547978 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477988 597980 478046
rect -1916 477978 78586 477988
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 39954 477978
rect 40010 477922 40078 477978
rect 40134 477922 40202 477978
rect 40258 477922 40326 477978
rect 40382 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477932 78586 477978
rect 78642 477932 78710 477988
rect 78766 477932 78834 477988
rect 78890 477932 78958 477988
rect 79014 477978 597980 477988
rect 79014 477932 132114 477978
rect 71102 477922 132114 477932
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 209878 477978
rect 209934 477922 210002 477978
rect 210058 477922 240598 477978
rect 240654 477922 240722 477978
rect 240778 477922 271318 477978
rect 271374 477922 271442 477978
rect 271498 477922 302038 477978
rect 302094 477922 302162 477978
rect 302218 477922 332758 477978
rect 332814 477922 332882 477978
rect 332938 477922 363478 477978
rect 363534 477922 363602 477978
rect 363658 477922 394198 477978
rect 394254 477922 394322 477978
rect 394378 477922 424918 477978
rect 424974 477922 425042 477978
rect 425098 477922 455638 477978
rect 455694 477922 455762 477978
rect 455818 477922 486358 477978
rect 486414 477922 486482 477978
rect 486538 477922 517078 477978
rect 517134 477922 517202 477978
rect 517258 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 547798 477978
rect 547854 477922 547922 477978
rect 547978 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 194518 472350
rect 194574 472294 194642 472350
rect 194698 472294 225238 472350
rect 225294 472294 225362 472350
rect 225418 472294 255958 472350
rect 256014 472294 256082 472350
rect 256138 472294 286678 472350
rect 286734 472294 286802 472350
rect 286858 472294 317398 472350
rect 317454 472294 317522 472350
rect 317578 472294 348118 472350
rect 348174 472294 348242 472350
rect 348298 472294 378838 472350
rect 378894 472294 378962 472350
rect 379018 472294 409558 472350
rect 409614 472294 409682 472350
rect 409738 472294 440278 472350
rect 440334 472294 440402 472350
rect 440458 472294 470998 472350
rect 471054 472294 471122 472350
rect 471178 472294 501718 472350
rect 501774 472294 501842 472350
rect 501898 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 532438 472350
rect 532494 472294 532562 472350
rect 532618 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 194518 472226
rect 194574 472170 194642 472226
rect 194698 472170 225238 472226
rect 225294 472170 225362 472226
rect 225418 472170 255958 472226
rect 256014 472170 256082 472226
rect 256138 472170 286678 472226
rect 286734 472170 286802 472226
rect 286858 472170 317398 472226
rect 317454 472170 317522 472226
rect 317578 472170 348118 472226
rect 348174 472170 348242 472226
rect 348298 472170 378838 472226
rect 378894 472170 378962 472226
rect 379018 472170 409558 472226
rect 409614 472170 409682 472226
rect 409738 472170 440278 472226
rect 440334 472170 440402 472226
rect 440458 472170 470998 472226
rect 471054 472170 471122 472226
rect 471178 472170 501718 472226
rect 501774 472170 501842 472226
rect 501898 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 532438 472226
rect 532494 472170 532562 472226
rect 532618 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 194518 472102
rect 194574 472046 194642 472102
rect 194698 472046 225238 472102
rect 225294 472046 225362 472102
rect 225418 472046 255958 472102
rect 256014 472046 256082 472102
rect 256138 472046 286678 472102
rect 286734 472046 286802 472102
rect 286858 472046 317398 472102
rect 317454 472046 317522 472102
rect 317578 472046 348118 472102
rect 348174 472046 348242 472102
rect 348298 472046 378838 472102
rect 378894 472046 378962 472102
rect 379018 472046 409558 472102
rect 409614 472046 409682 472102
rect 409738 472046 440278 472102
rect 440334 472046 440402 472102
rect 440458 472046 470998 472102
rect 471054 472046 471122 472102
rect 471178 472046 501718 472102
rect 501774 472046 501842 472102
rect 501898 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 532438 472102
rect 532494 472046 532562 472102
rect 532618 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 194518 471978
rect 194574 471922 194642 471978
rect 194698 471922 225238 471978
rect 225294 471922 225362 471978
rect 225418 471922 255958 471978
rect 256014 471922 256082 471978
rect 256138 471922 286678 471978
rect 286734 471922 286802 471978
rect 286858 471922 317398 471978
rect 317454 471922 317522 471978
rect 317578 471922 348118 471978
rect 348174 471922 348242 471978
rect 348298 471922 378838 471978
rect 378894 471922 378962 471978
rect 379018 471922 409558 471978
rect 409614 471922 409682 471978
rect 409738 471922 440278 471978
rect 440334 471922 440402 471978
rect 440458 471922 470998 471978
rect 471054 471922 471122 471978
rect 471178 471922 501718 471978
rect 501774 471922 501842 471978
rect 501898 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 532438 471978
rect 532494 471922 532562 471978
rect 532618 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 39954 460350
rect 40010 460294 40078 460350
rect 40134 460294 40202 460350
rect 40258 460294 40326 460350
rect 40382 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 101394 460350
rect 101450 460294 101518 460350
rect 101574 460294 101642 460350
rect 101698 460294 101766 460350
rect 101822 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 209878 460350
rect 209934 460294 210002 460350
rect 210058 460294 240598 460350
rect 240654 460294 240722 460350
rect 240778 460294 271318 460350
rect 271374 460294 271442 460350
rect 271498 460294 302038 460350
rect 302094 460294 302162 460350
rect 302218 460294 332758 460350
rect 332814 460294 332882 460350
rect 332938 460294 363478 460350
rect 363534 460294 363602 460350
rect 363658 460294 394198 460350
rect 394254 460294 394322 460350
rect 394378 460294 424918 460350
rect 424974 460294 425042 460350
rect 425098 460294 455638 460350
rect 455694 460294 455762 460350
rect 455818 460294 486358 460350
rect 486414 460294 486482 460350
rect 486538 460294 517078 460350
rect 517134 460294 517202 460350
rect 517258 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 547798 460350
rect 547854 460294 547922 460350
rect 547978 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 39954 460226
rect 40010 460170 40078 460226
rect 40134 460170 40202 460226
rect 40258 460170 40326 460226
rect 40382 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 101394 460226
rect 101450 460170 101518 460226
rect 101574 460170 101642 460226
rect 101698 460170 101766 460226
rect 101822 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 209878 460226
rect 209934 460170 210002 460226
rect 210058 460170 240598 460226
rect 240654 460170 240722 460226
rect 240778 460170 271318 460226
rect 271374 460170 271442 460226
rect 271498 460170 302038 460226
rect 302094 460170 302162 460226
rect 302218 460170 332758 460226
rect 332814 460170 332882 460226
rect 332938 460170 363478 460226
rect 363534 460170 363602 460226
rect 363658 460170 394198 460226
rect 394254 460170 394322 460226
rect 394378 460170 424918 460226
rect 424974 460170 425042 460226
rect 425098 460170 455638 460226
rect 455694 460170 455762 460226
rect 455818 460170 486358 460226
rect 486414 460170 486482 460226
rect 486538 460170 517078 460226
rect 517134 460170 517202 460226
rect 517258 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 547798 460226
rect 547854 460170 547922 460226
rect 547978 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 39954 460102
rect 40010 460046 40078 460102
rect 40134 460046 40202 460102
rect 40258 460046 40326 460102
rect 40382 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 101394 460102
rect 101450 460046 101518 460102
rect 101574 460046 101642 460102
rect 101698 460046 101766 460102
rect 101822 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 209878 460102
rect 209934 460046 210002 460102
rect 210058 460046 240598 460102
rect 240654 460046 240722 460102
rect 240778 460046 271318 460102
rect 271374 460046 271442 460102
rect 271498 460046 302038 460102
rect 302094 460046 302162 460102
rect 302218 460046 332758 460102
rect 332814 460046 332882 460102
rect 332938 460046 363478 460102
rect 363534 460046 363602 460102
rect 363658 460046 394198 460102
rect 394254 460046 394322 460102
rect 394378 460046 424918 460102
rect 424974 460046 425042 460102
rect 425098 460046 455638 460102
rect 455694 460046 455762 460102
rect 455818 460046 486358 460102
rect 486414 460046 486482 460102
rect 486538 460046 517078 460102
rect 517134 460046 517202 460102
rect 517258 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 547798 460102
rect 547854 460046 547922 460102
rect 547978 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 39954 459978
rect 40010 459922 40078 459978
rect 40134 459922 40202 459978
rect 40258 459922 40326 459978
rect 40382 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 101394 459978
rect 101450 459922 101518 459978
rect 101574 459922 101642 459978
rect 101698 459922 101766 459978
rect 101822 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 209878 459978
rect 209934 459922 210002 459978
rect 210058 459922 240598 459978
rect 240654 459922 240722 459978
rect 240778 459922 271318 459978
rect 271374 459922 271442 459978
rect 271498 459922 302038 459978
rect 302094 459922 302162 459978
rect 302218 459922 332758 459978
rect 332814 459922 332882 459978
rect 332938 459922 363478 459978
rect 363534 459922 363602 459978
rect 363658 459922 394198 459978
rect 394254 459922 394322 459978
rect 394378 459922 424918 459978
rect 424974 459922 425042 459978
rect 425098 459922 455638 459978
rect 455694 459922 455762 459978
rect 455818 459922 486358 459978
rect 486414 459922 486482 459978
rect 486538 459922 517078 459978
rect 517134 459922 517202 459978
rect 517258 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 547798 459978
rect 547854 459922 547922 459978
rect 547978 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 194518 454350
rect 194574 454294 194642 454350
rect 194698 454294 225238 454350
rect 225294 454294 225362 454350
rect 225418 454294 255958 454350
rect 256014 454294 256082 454350
rect 256138 454294 286678 454350
rect 286734 454294 286802 454350
rect 286858 454294 317398 454350
rect 317454 454294 317522 454350
rect 317578 454294 348118 454350
rect 348174 454294 348242 454350
rect 348298 454294 378838 454350
rect 378894 454294 378962 454350
rect 379018 454294 409558 454350
rect 409614 454294 409682 454350
rect 409738 454294 440278 454350
rect 440334 454294 440402 454350
rect 440458 454294 470998 454350
rect 471054 454294 471122 454350
rect 471178 454294 501718 454350
rect 501774 454294 501842 454350
rect 501898 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 532438 454350
rect 532494 454294 532562 454350
rect 532618 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 194518 454226
rect 194574 454170 194642 454226
rect 194698 454170 225238 454226
rect 225294 454170 225362 454226
rect 225418 454170 255958 454226
rect 256014 454170 256082 454226
rect 256138 454170 286678 454226
rect 286734 454170 286802 454226
rect 286858 454170 317398 454226
rect 317454 454170 317522 454226
rect 317578 454170 348118 454226
rect 348174 454170 348242 454226
rect 348298 454170 378838 454226
rect 378894 454170 378962 454226
rect 379018 454170 409558 454226
rect 409614 454170 409682 454226
rect 409738 454170 440278 454226
rect 440334 454170 440402 454226
rect 440458 454170 470998 454226
rect 471054 454170 471122 454226
rect 471178 454170 501718 454226
rect 501774 454170 501842 454226
rect 501898 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 532438 454226
rect 532494 454170 532562 454226
rect 532618 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 194518 454102
rect 194574 454046 194642 454102
rect 194698 454046 225238 454102
rect 225294 454046 225362 454102
rect 225418 454046 255958 454102
rect 256014 454046 256082 454102
rect 256138 454046 286678 454102
rect 286734 454046 286802 454102
rect 286858 454046 317398 454102
rect 317454 454046 317522 454102
rect 317578 454046 348118 454102
rect 348174 454046 348242 454102
rect 348298 454046 378838 454102
rect 378894 454046 378962 454102
rect 379018 454046 409558 454102
rect 409614 454046 409682 454102
rect 409738 454046 440278 454102
rect 440334 454046 440402 454102
rect 440458 454046 470998 454102
rect 471054 454046 471122 454102
rect 471178 454046 501718 454102
rect 501774 454046 501842 454102
rect 501898 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 532438 454102
rect 532494 454046 532562 454102
rect 532618 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 194518 453978
rect 194574 453922 194642 453978
rect 194698 453922 225238 453978
rect 225294 453922 225362 453978
rect 225418 453922 255958 453978
rect 256014 453922 256082 453978
rect 256138 453922 286678 453978
rect 286734 453922 286802 453978
rect 286858 453922 317398 453978
rect 317454 453922 317522 453978
rect 317578 453922 348118 453978
rect 348174 453922 348242 453978
rect 348298 453922 378838 453978
rect 378894 453922 378962 453978
rect 379018 453922 409558 453978
rect 409614 453922 409682 453978
rect 409738 453922 440278 453978
rect 440334 453922 440402 453978
rect 440458 453922 470998 453978
rect 471054 453922 471122 453978
rect 471178 453922 501718 453978
rect 501774 453922 501842 453978
rect 501898 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 532438 453978
rect 532494 453922 532562 453978
rect 532618 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 39954 442350
rect 40010 442294 40078 442350
rect 40134 442294 40202 442350
rect 40258 442294 40326 442350
rect 40382 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 101394 442350
rect 101450 442294 101518 442350
rect 101574 442294 101642 442350
rect 101698 442294 101766 442350
rect 101822 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 209878 442350
rect 209934 442294 210002 442350
rect 210058 442294 240598 442350
rect 240654 442294 240722 442350
rect 240778 442294 271318 442350
rect 271374 442294 271442 442350
rect 271498 442294 302038 442350
rect 302094 442294 302162 442350
rect 302218 442294 332758 442350
rect 332814 442294 332882 442350
rect 332938 442294 363478 442350
rect 363534 442294 363602 442350
rect 363658 442294 394198 442350
rect 394254 442294 394322 442350
rect 394378 442294 424918 442350
rect 424974 442294 425042 442350
rect 425098 442294 455638 442350
rect 455694 442294 455762 442350
rect 455818 442294 486358 442350
rect 486414 442294 486482 442350
rect 486538 442294 517078 442350
rect 517134 442294 517202 442350
rect 517258 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 547798 442350
rect 547854 442294 547922 442350
rect 547978 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 39954 442226
rect 40010 442170 40078 442226
rect 40134 442170 40202 442226
rect 40258 442170 40326 442226
rect 40382 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 101394 442226
rect 101450 442170 101518 442226
rect 101574 442170 101642 442226
rect 101698 442170 101766 442226
rect 101822 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 209878 442226
rect 209934 442170 210002 442226
rect 210058 442170 240598 442226
rect 240654 442170 240722 442226
rect 240778 442170 271318 442226
rect 271374 442170 271442 442226
rect 271498 442170 302038 442226
rect 302094 442170 302162 442226
rect 302218 442170 332758 442226
rect 332814 442170 332882 442226
rect 332938 442170 363478 442226
rect 363534 442170 363602 442226
rect 363658 442170 394198 442226
rect 394254 442170 394322 442226
rect 394378 442170 424918 442226
rect 424974 442170 425042 442226
rect 425098 442170 455638 442226
rect 455694 442170 455762 442226
rect 455818 442170 486358 442226
rect 486414 442170 486482 442226
rect 486538 442170 517078 442226
rect 517134 442170 517202 442226
rect 517258 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 547798 442226
rect 547854 442170 547922 442226
rect 547978 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 39954 442102
rect 40010 442046 40078 442102
rect 40134 442046 40202 442102
rect 40258 442046 40326 442102
rect 40382 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 101394 442102
rect 101450 442046 101518 442102
rect 101574 442046 101642 442102
rect 101698 442046 101766 442102
rect 101822 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 209878 442102
rect 209934 442046 210002 442102
rect 210058 442046 240598 442102
rect 240654 442046 240722 442102
rect 240778 442046 271318 442102
rect 271374 442046 271442 442102
rect 271498 442046 302038 442102
rect 302094 442046 302162 442102
rect 302218 442046 332758 442102
rect 332814 442046 332882 442102
rect 332938 442046 363478 442102
rect 363534 442046 363602 442102
rect 363658 442046 394198 442102
rect 394254 442046 394322 442102
rect 394378 442046 424918 442102
rect 424974 442046 425042 442102
rect 425098 442046 455638 442102
rect 455694 442046 455762 442102
rect 455818 442046 486358 442102
rect 486414 442046 486482 442102
rect 486538 442046 517078 442102
rect 517134 442046 517202 442102
rect 517258 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 547798 442102
rect 547854 442046 547922 442102
rect 547978 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 39954 441978
rect 40010 441922 40078 441978
rect 40134 441922 40202 441978
rect 40258 441922 40326 441978
rect 40382 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 101394 441978
rect 101450 441922 101518 441978
rect 101574 441922 101642 441978
rect 101698 441922 101766 441978
rect 101822 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 209878 441978
rect 209934 441922 210002 441978
rect 210058 441922 240598 441978
rect 240654 441922 240722 441978
rect 240778 441922 271318 441978
rect 271374 441922 271442 441978
rect 271498 441922 302038 441978
rect 302094 441922 302162 441978
rect 302218 441922 332758 441978
rect 332814 441922 332882 441978
rect 332938 441922 363478 441978
rect 363534 441922 363602 441978
rect 363658 441922 394198 441978
rect 394254 441922 394322 441978
rect 394378 441922 424918 441978
rect 424974 441922 425042 441978
rect 425098 441922 455638 441978
rect 455694 441922 455762 441978
rect 455818 441922 486358 441978
rect 486414 441922 486482 441978
rect 486538 441922 517078 441978
rect 517134 441922 517202 441978
rect 517258 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 547798 441978
rect 547854 441922 547922 441978
rect 547978 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 194518 436350
rect 194574 436294 194642 436350
rect 194698 436294 225238 436350
rect 225294 436294 225362 436350
rect 225418 436294 255958 436350
rect 256014 436294 256082 436350
rect 256138 436294 286678 436350
rect 286734 436294 286802 436350
rect 286858 436294 317398 436350
rect 317454 436294 317522 436350
rect 317578 436294 348118 436350
rect 348174 436294 348242 436350
rect 348298 436294 378838 436350
rect 378894 436294 378962 436350
rect 379018 436294 409558 436350
rect 409614 436294 409682 436350
rect 409738 436294 440278 436350
rect 440334 436294 440402 436350
rect 440458 436294 470998 436350
rect 471054 436294 471122 436350
rect 471178 436294 501718 436350
rect 501774 436294 501842 436350
rect 501898 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 532438 436350
rect 532494 436294 532562 436350
rect 532618 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 194518 436226
rect 194574 436170 194642 436226
rect 194698 436170 225238 436226
rect 225294 436170 225362 436226
rect 225418 436170 255958 436226
rect 256014 436170 256082 436226
rect 256138 436170 286678 436226
rect 286734 436170 286802 436226
rect 286858 436170 317398 436226
rect 317454 436170 317522 436226
rect 317578 436170 348118 436226
rect 348174 436170 348242 436226
rect 348298 436170 378838 436226
rect 378894 436170 378962 436226
rect 379018 436170 409558 436226
rect 409614 436170 409682 436226
rect 409738 436170 440278 436226
rect 440334 436170 440402 436226
rect 440458 436170 470998 436226
rect 471054 436170 471122 436226
rect 471178 436170 501718 436226
rect 501774 436170 501842 436226
rect 501898 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 532438 436226
rect 532494 436170 532562 436226
rect 532618 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 194518 436102
rect 194574 436046 194642 436102
rect 194698 436046 225238 436102
rect 225294 436046 225362 436102
rect 225418 436046 255958 436102
rect 256014 436046 256082 436102
rect 256138 436046 286678 436102
rect 286734 436046 286802 436102
rect 286858 436046 317398 436102
rect 317454 436046 317522 436102
rect 317578 436046 348118 436102
rect 348174 436046 348242 436102
rect 348298 436046 378838 436102
rect 378894 436046 378962 436102
rect 379018 436046 409558 436102
rect 409614 436046 409682 436102
rect 409738 436046 440278 436102
rect 440334 436046 440402 436102
rect 440458 436046 470998 436102
rect 471054 436046 471122 436102
rect 471178 436046 501718 436102
rect 501774 436046 501842 436102
rect 501898 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 532438 436102
rect 532494 436046 532562 436102
rect 532618 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 194518 435978
rect 194574 435922 194642 435978
rect 194698 435922 225238 435978
rect 225294 435922 225362 435978
rect 225418 435922 255958 435978
rect 256014 435922 256082 435978
rect 256138 435922 286678 435978
rect 286734 435922 286802 435978
rect 286858 435922 317398 435978
rect 317454 435922 317522 435978
rect 317578 435922 348118 435978
rect 348174 435922 348242 435978
rect 348298 435922 378838 435978
rect 378894 435922 378962 435978
rect 379018 435922 409558 435978
rect 409614 435922 409682 435978
rect 409738 435922 440278 435978
rect 440334 435922 440402 435978
rect 440458 435922 470998 435978
rect 471054 435922 471122 435978
rect 471178 435922 501718 435978
rect 501774 435922 501842 435978
rect 501898 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 532438 435978
rect 532494 435922 532562 435978
rect 532618 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 39954 424350
rect 40010 424294 40078 424350
rect 40134 424294 40202 424350
rect 40258 424294 40326 424350
rect 40382 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 101394 424350
rect 101450 424294 101518 424350
rect 101574 424294 101642 424350
rect 101698 424294 101766 424350
rect 101822 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 209878 424350
rect 209934 424294 210002 424350
rect 210058 424294 240598 424350
rect 240654 424294 240722 424350
rect 240778 424294 271318 424350
rect 271374 424294 271442 424350
rect 271498 424294 302038 424350
rect 302094 424294 302162 424350
rect 302218 424294 332758 424350
rect 332814 424294 332882 424350
rect 332938 424294 363478 424350
rect 363534 424294 363602 424350
rect 363658 424294 394198 424350
rect 394254 424294 394322 424350
rect 394378 424294 424918 424350
rect 424974 424294 425042 424350
rect 425098 424294 455638 424350
rect 455694 424294 455762 424350
rect 455818 424294 486358 424350
rect 486414 424294 486482 424350
rect 486538 424294 517078 424350
rect 517134 424294 517202 424350
rect 517258 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 547798 424350
rect 547854 424294 547922 424350
rect 547978 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 39954 424226
rect 40010 424170 40078 424226
rect 40134 424170 40202 424226
rect 40258 424170 40326 424226
rect 40382 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 101394 424226
rect 101450 424170 101518 424226
rect 101574 424170 101642 424226
rect 101698 424170 101766 424226
rect 101822 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 209878 424226
rect 209934 424170 210002 424226
rect 210058 424170 240598 424226
rect 240654 424170 240722 424226
rect 240778 424170 271318 424226
rect 271374 424170 271442 424226
rect 271498 424170 302038 424226
rect 302094 424170 302162 424226
rect 302218 424170 332758 424226
rect 332814 424170 332882 424226
rect 332938 424170 363478 424226
rect 363534 424170 363602 424226
rect 363658 424170 394198 424226
rect 394254 424170 394322 424226
rect 394378 424170 424918 424226
rect 424974 424170 425042 424226
rect 425098 424170 455638 424226
rect 455694 424170 455762 424226
rect 455818 424170 486358 424226
rect 486414 424170 486482 424226
rect 486538 424170 517078 424226
rect 517134 424170 517202 424226
rect 517258 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 547798 424226
rect 547854 424170 547922 424226
rect 547978 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 39954 424102
rect 40010 424046 40078 424102
rect 40134 424046 40202 424102
rect 40258 424046 40326 424102
rect 40382 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 101394 424102
rect 101450 424046 101518 424102
rect 101574 424046 101642 424102
rect 101698 424046 101766 424102
rect 101822 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 209878 424102
rect 209934 424046 210002 424102
rect 210058 424046 240598 424102
rect 240654 424046 240722 424102
rect 240778 424046 271318 424102
rect 271374 424046 271442 424102
rect 271498 424046 302038 424102
rect 302094 424046 302162 424102
rect 302218 424046 332758 424102
rect 332814 424046 332882 424102
rect 332938 424046 363478 424102
rect 363534 424046 363602 424102
rect 363658 424046 394198 424102
rect 394254 424046 394322 424102
rect 394378 424046 424918 424102
rect 424974 424046 425042 424102
rect 425098 424046 455638 424102
rect 455694 424046 455762 424102
rect 455818 424046 486358 424102
rect 486414 424046 486482 424102
rect 486538 424046 517078 424102
rect 517134 424046 517202 424102
rect 517258 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 547798 424102
rect 547854 424046 547922 424102
rect 547978 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 39954 423978
rect 40010 423922 40078 423978
rect 40134 423922 40202 423978
rect 40258 423922 40326 423978
rect 40382 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 101394 423978
rect 101450 423922 101518 423978
rect 101574 423922 101642 423978
rect 101698 423922 101766 423978
rect 101822 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 209878 423978
rect 209934 423922 210002 423978
rect 210058 423922 240598 423978
rect 240654 423922 240722 423978
rect 240778 423922 271318 423978
rect 271374 423922 271442 423978
rect 271498 423922 302038 423978
rect 302094 423922 302162 423978
rect 302218 423922 332758 423978
rect 332814 423922 332882 423978
rect 332938 423922 363478 423978
rect 363534 423922 363602 423978
rect 363658 423922 394198 423978
rect 394254 423922 394322 423978
rect 394378 423922 424918 423978
rect 424974 423922 425042 423978
rect 425098 423922 455638 423978
rect 455694 423922 455762 423978
rect 455818 423922 486358 423978
rect 486414 423922 486482 423978
rect 486538 423922 517078 423978
rect 517134 423922 517202 423978
rect 517258 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 547798 423978
rect 547854 423922 547922 423978
rect 547978 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect 190636 421858 192404 421874
rect 190636 421802 190652 421858
rect 190708 421802 192332 421858
rect 192388 421802 192404 421858
rect 190636 421786 192404 421802
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 194518 418350
rect 194574 418294 194642 418350
rect 194698 418294 225238 418350
rect 225294 418294 225362 418350
rect 225418 418294 255958 418350
rect 256014 418294 256082 418350
rect 256138 418294 286678 418350
rect 286734 418294 286802 418350
rect 286858 418294 317398 418350
rect 317454 418294 317522 418350
rect 317578 418294 348118 418350
rect 348174 418294 348242 418350
rect 348298 418294 378838 418350
rect 378894 418294 378962 418350
rect 379018 418294 409558 418350
rect 409614 418294 409682 418350
rect 409738 418294 440278 418350
rect 440334 418294 440402 418350
rect 440458 418294 470998 418350
rect 471054 418294 471122 418350
rect 471178 418294 501718 418350
rect 501774 418294 501842 418350
rect 501898 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 532438 418350
rect 532494 418294 532562 418350
rect 532618 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 194518 418226
rect 194574 418170 194642 418226
rect 194698 418170 225238 418226
rect 225294 418170 225362 418226
rect 225418 418170 255958 418226
rect 256014 418170 256082 418226
rect 256138 418170 286678 418226
rect 286734 418170 286802 418226
rect 286858 418170 317398 418226
rect 317454 418170 317522 418226
rect 317578 418170 348118 418226
rect 348174 418170 348242 418226
rect 348298 418170 378838 418226
rect 378894 418170 378962 418226
rect 379018 418170 409558 418226
rect 409614 418170 409682 418226
rect 409738 418170 440278 418226
rect 440334 418170 440402 418226
rect 440458 418170 470998 418226
rect 471054 418170 471122 418226
rect 471178 418170 501718 418226
rect 501774 418170 501842 418226
rect 501898 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 532438 418226
rect 532494 418170 532562 418226
rect 532618 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 194518 418102
rect 194574 418046 194642 418102
rect 194698 418046 225238 418102
rect 225294 418046 225362 418102
rect 225418 418046 255958 418102
rect 256014 418046 256082 418102
rect 256138 418046 286678 418102
rect 286734 418046 286802 418102
rect 286858 418046 317398 418102
rect 317454 418046 317522 418102
rect 317578 418046 348118 418102
rect 348174 418046 348242 418102
rect 348298 418046 378838 418102
rect 378894 418046 378962 418102
rect 379018 418046 409558 418102
rect 409614 418046 409682 418102
rect 409738 418046 440278 418102
rect 440334 418046 440402 418102
rect 440458 418046 470998 418102
rect 471054 418046 471122 418102
rect 471178 418046 501718 418102
rect 501774 418046 501842 418102
rect 501898 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 532438 418102
rect 532494 418046 532562 418102
rect 532618 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 194518 417978
rect 194574 417922 194642 417978
rect 194698 417922 225238 417978
rect 225294 417922 225362 417978
rect 225418 417922 255958 417978
rect 256014 417922 256082 417978
rect 256138 417922 286678 417978
rect 286734 417922 286802 417978
rect 286858 417922 317398 417978
rect 317454 417922 317522 417978
rect 317578 417922 348118 417978
rect 348174 417922 348242 417978
rect 348298 417922 378838 417978
rect 378894 417922 378962 417978
rect 379018 417922 409558 417978
rect 409614 417922 409682 417978
rect 409738 417922 440278 417978
rect 440334 417922 440402 417978
rect 440458 417922 470998 417978
rect 471054 417922 471122 417978
rect 471178 417922 501718 417978
rect 501774 417922 501842 417978
rect 501898 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 532438 417978
rect 532494 417922 532562 417978
rect 532618 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect 357180 411058 568724 411074
rect 357180 411002 357196 411058
rect 357252 411002 568652 411058
rect 568708 411002 568724 411058
rect 357180 410986 568724 411002
rect 334220 410878 556180 410894
rect 334220 410822 334236 410878
rect 334292 410822 556108 410878
rect 556164 410822 556180 410878
rect 334220 410806 556180 410822
rect 324140 410698 556516 410714
rect 324140 410642 324156 410698
rect 324212 410642 556444 410698
rect 556500 410642 556516 410698
rect 324140 410626 556516 410642
rect 358748 409978 519220 409994
rect 358748 409922 358764 409978
rect 358820 409922 519148 409978
rect 519204 409922 519220 409978
rect 358748 409906 519220 409922
rect 357292 409618 514964 409634
rect 357292 409562 357308 409618
rect 357364 409562 514892 409618
rect 514948 409562 514964 409618
rect 357292 409546 514964 409562
rect 358076 409438 584740 409454
rect 358076 409382 358092 409438
rect 358148 409382 584668 409438
rect 584724 409382 584740 409438
rect 358076 409366 584740 409382
rect 329180 409258 556292 409274
rect 329180 409202 329196 409258
rect 329252 409202 556220 409258
rect 556276 409202 556292 409258
rect 329180 409186 556292 409202
rect 357628 409078 585524 409094
rect 357628 409022 357644 409078
rect 357700 409022 585452 409078
rect 585508 409022 585524 409078
rect 357628 409006 585524 409022
rect 356172 408178 567044 408194
rect 356172 408122 356188 408178
rect 356244 408122 566972 408178
rect 567028 408122 567044 408178
rect 356172 408106 567044 408122
rect 243500 407638 357716 407654
rect 243500 407582 243516 407638
rect 243572 407582 357644 407638
rect 357700 407582 357716 407638
rect 243500 407566 357716 407582
rect 277100 407458 551252 407474
rect 277100 407402 277116 407458
rect 277172 407402 551180 407458
rect 551236 407402 551252 407458
rect 277100 407386 551252 407402
rect 360428 407098 533892 407114
rect 360428 407042 360444 407098
rect 360500 407042 533820 407098
rect 533876 407042 533892 407098
rect 360428 407026 533892 407042
rect 248876 406918 357828 406934
rect 248876 406862 248892 406918
rect 248948 406862 357756 406918
rect 357812 406862 357828 406918
rect 248876 406846 357828 406862
rect 358972 406918 539268 406934
rect 358972 406862 358988 406918
rect 359044 406862 539196 406918
rect 539252 406862 539268 406918
rect 358972 406846 539268 406862
rect 227596 406738 557860 406754
rect 227596 406682 227612 406738
rect 227668 406682 557788 406738
rect 557844 406682 557860 406738
rect 227596 406666 557860 406682
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 39954 406350
rect 40010 406294 40078 406350
rect 40134 406294 40202 406350
rect 40258 406294 40326 406350
rect 40382 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 101394 406350
rect 101450 406294 101518 406350
rect 101574 406294 101642 406350
rect 101698 406294 101766 406350
rect 101822 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 285714 406350
rect 285770 406294 285838 406350
rect 285894 406294 285962 406350
rect 286018 406294 286086 406350
rect 286142 406294 316434 406350
rect 316490 406294 316558 406350
rect 316614 406294 316682 406350
rect 316738 406294 316806 406350
rect 316862 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 39954 406226
rect 40010 406170 40078 406226
rect 40134 406170 40202 406226
rect 40258 406170 40326 406226
rect 40382 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 101394 406226
rect 101450 406170 101518 406226
rect 101574 406170 101642 406226
rect 101698 406170 101766 406226
rect 101822 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 285714 406226
rect 285770 406170 285838 406226
rect 285894 406170 285962 406226
rect 286018 406170 286086 406226
rect 286142 406170 316434 406226
rect 316490 406170 316558 406226
rect 316614 406170 316682 406226
rect 316738 406170 316806 406226
rect 316862 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 39954 406102
rect 40010 406046 40078 406102
rect 40134 406046 40202 406102
rect 40258 406046 40326 406102
rect 40382 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 101394 406102
rect 101450 406046 101518 406102
rect 101574 406046 101642 406102
rect 101698 406046 101766 406102
rect 101822 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 285714 406102
rect 285770 406046 285838 406102
rect 285894 406046 285962 406102
rect 286018 406046 286086 406102
rect 286142 406046 316434 406102
rect 316490 406046 316558 406102
rect 316614 406046 316682 406102
rect 316738 406046 316806 406102
rect 316862 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 39954 405978
rect 40010 405922 40078 405978
rect 40134 405922 40202 405978
rect 40258 405922 40326 405978
rect 40382 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 101394 405978
rect 101450 405922 101518 405978
rect 101574 405922 101642 405978
rect 101698 405922 101766 405978
rect 101822 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 285714 405978
rect 285770 405922 285838 405978
rect 285894 405922 285962 405978
rect 286018 405922 286086 405978
rect 286142 405922 316434 405978
rect 316490 405922 316558 405978
rect 316614 405922 316682 405978
rect 316738 405922 316806 405978
rect 316862 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect 330860 405658 552820 405674
rect 330860 405602 330876 405658
rect 330932 405602 552748 405658
rect 552804 405602 552820 405658
rect 330860 405586 552820 405602
rect 209900 404578 560324 404594
rect 209900 404522 209916 404578
rect 209972 404522 560252 404578
rect 560308 404522 560324 404578
rect 209900 404506 560324 404522
rect 208220 404398 565364 404414
rect 208220 404342 208236 404398
rect 208292 404342 565292 404398
rect 565348 404342 565364 404398
rect 208220 404326 565364 404342
rect 206540 404218 570404 404234
rect 206540 404162 206556 404218
rect 206612 404162 570332 404218
rect 570388 404162 570404 404218
rect 206540 404146 570404 404162
rect 186156 404038 590564 404054
rect 186156 403982 186172 404038
rect 186228 403982 590492 404038
rect 590548 403982 590564 404038
rect 186156 403966 590564 403982
rect 185932 402418 590676 402434
rect 185932 402362 185948 402418
rect 186004 402362 590604 402418
rect 590660 402362 590676 402418
rect 185932 402346 590676 402362
rect 196460 402058 572084 402074
rect 196460 402002 196476 402058
rect 196532 402002 572012 402058
rect 572068 402002 572084 402058
rect 196460 401986 572084 402002
rect 198140 401878 573764 401894
rect 198140 401822 198156 401878
rect 198212 401822 573692 401878
rect 573748 401822 573764 401878
rect 198140 401806 573764 401822
rect 199820 401698 575444 401714
rect 199820 401642 199836 401698
rect 199892 401642 575372 401698
rect 575428 401642 575444 401698
rect 199820 401626 575444 401642
rect 319100 400618 549460 400634
rect 319100 400562 319116 400618
rect 319172 400562 549388 400618
rect 549444 400562 549460 400618
rect 319100 400546 549460 400562
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 97674 400350
rect 97730 400294 97798 400350
rect 97854 400294 97922 400350
rect 97978 400294 98046 400350
rect 98102 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 281994 400350
rect 282050 400294 282118 400350
rect 282174 400294 282242 400350
rect 282298 400294 282366 400350
rect 282422 400294 312714 400350
rect 312770 400294 312838 400350
rect 312894 400294 312962 400350
rect 313018 400294 313086 400350
rect 313142 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 97674 400226
rect 97730 400170 97798 400226
rect 97854 400170 97922 400226
rect 97978 400170 98046 400226
rect 98102 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 281994 400226
rect 282050 400170 282118 400226
rect 282174 400170 282242 400226
rect 282298 400170 282366 400226
rect 282422 400170 312714 400226
rect 312770 400170 312838 400226
rect 312894 400170 312962 400226
rect 313018 400170 313086 400226
rect 313142 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 97674 400102
rect 97730 400046 97798 400102
rect 97854 400046 97922 400102
rect 97978 400046 98046 400102
rect 98102 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 281994 400102
rect 282050 400046 282118 400102
rect 282174 400046 282242 400102
rect 282298 400046 282366 400102
rect 282422 400046 312714 400102
rect 312770 400046 312838 400102
rect 312894 400046 312962 400102
rect 313018 400046 313086 400102
rect 313142 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 97674 399978
rect 97730 399922 97798 399978
rect 97854 399922 97922 399978
rect 97978 399922 98046 399978
rect 98102 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 281994 399978
rect 282050 399922 282118 399978
rect 282174 399922 282242 399978
rect 282298 399922 282366 399978
rect 282422 399922 312714 399978
rect 312770 399922 312838 399978
rect 312894 399922 312962 399978
rect 313018 399922 313086 399978
rect 313142 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect 320780 399358 556404 399374
rect 320780 399302 320796 399358
rect 320852 399302 556332 399358
rect 556388 399302 556404 399358
rect 320780 399286 556404 399302
rect 307340 399178 551140 399194
rect 307340 399122 307356 399178
rect 307412 399122 551068 399178
rect 551124 399122 551140 399178
rect 307340 399106 551140 399122
rect 305660 398998 549572 399014
rect 305660 398942 305676 398998
rect 305732 398942 549500 398998
rect 549556 398942 549572 398998
rect 305660 398926 549572 398942
rect 344076 398278 559540 398294
rect 344076 398222 344092 398278
rect 344148 398222 559468 398278
rect 559524 398222 559540 398278
rect 344076 398206 559540 398222
rect 349004 397198 526500 397214
rect 349004 397142 349020 397198
rect 349076 397142 526428 397198
rect 526484 397142 526500 397198
rect 349004 397126 526500 397142
rect 353484 397018 532548 397034
rect 353484 396962 353500 397018
rect 353556 396962 532476 397018
rect 532532 396962 532548 397018
rect 353484 396946 532548 396962
rect 355836 396838 556740 396854
rect 355836 396782 355852 396838
rect 355908 396782 556668 396838
rect 556724 396782 556740 396838
rect 355836 396766 556740 396782
rect 345532 396658 550692 396674
rect 345532 396602 345548 396658
rect 345604 396602 550620 396658
rect 550676 396602 550692 396658
rect 345532 396586 550692 396602
rect 362108 395578 375524 395594
rect 362108 395522 362124 395578
rect 362180 395522 375452 395578
rect 375508 395522 375524 395578
rect 362108 395506 375524 395522
rect 344188 395398 559652 395414
rect 344188 395342 344204 395398
rect 344260 395342 559580 395398
rect 559636 395342 559652 395398
rect 344188 395326 559652 395342
rect 231628 395218 581380 395234
rect 231628 395162 231644 395218
rect 231700 395162 581308 395218
rect 581364 395162 581380 395218
rect 231628 395146 581380 395162
rect 231740 395038 583060 395054
rect 231740 394982 231756 395038
rect 231812 394982 582988 395038
rect 583044 394982 583060 395038
rect 231740 394966 583060 394982
rect 354380 394858 538596 394874
rect 354380 394802 354396 394858
rect 354452 394802 538524 394858
rect 538580 394802 538596 394858
rect 354380 394786 538596 394802
rect 230060 393778 579700 393794
rect 230060 393722 230076 393778
rect 230132 393722 579628 393778
rect 579684 393722 579700 393778
rect 230060 393706 579700 393722
rect 199708 393598 570404 393614
rect 199708 393542 199724 393598
rect 199780 393542 570332 393598
rect 570388 393542 570404 393598
rect 199708 393526 570404 393542
rect 201500 393418 577124 393434
rect 201500 393362 201516 393418
rect 201572 393362 577052 393418
rect 577108 393362 577124 393418
rect 201500 393346 577124 393362
rect 198028 393238 585524 393254
rect 198028 393182 198044 393238
rect 198100 393182 585452 393238
rect 585508 393182 585524 393238
rect 198028 393166 585524 393182
rect 341948 392338 441828 392354
rect 341948 392282 341964 392338
rect 342020 392282 441756 392338
rect 441812 392282 441828 392338
rect 341948 392266 441828 392282
rect 204860 392158 590564 392174
rect 204860 392102 204876 392158
rect 204932 392102 590492 392158
rect 590548 392102 590564 392158
rect 204860 392086 590564 392102
rect 201388 391978 361972 391994
rect 201388 391922 201404 391978
rect 201460 391922 361900 391978
rect 361956 391922 361972 391978
rect 201388 391906 361972 391922
rect 197468 391798 362196 391814
rect 197468 391742 197484 391798
rect 197540 391742 362124 391798
rect 362180 391742 362196 391798
rect 197468 391726 362196 391742
rect 215052 391438 361748 391454
rect 215052 391382 215068 391438
rect 215124 391382 216636 391438
rect 216692 391382 361676 391438
rect 361732 391382 361748 391438
rect 215052 391366 361748 391382
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 39954 388350
rect 40010 388294 40078 388350
rect 40134 388294 40202 388350
rect 40258 388294 40326 388350
rect 40382 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 101394 388350
rect 101450 388294 101518 388350
rect 101574 388294 101642 388350
rect 101698 388294 101766 388350
rect 101822 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 285714 388350
rect 285770 388294 285838 388350
rect 285894 388294 285962 388350
rect 286018 388294 286086 388350
rect 286142 388294 316434 388350
rect 316490 388294 316558 388350
rect 316614 388294 316682 388350
rect 316738 388294 316806 388350
rect 316862 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 379878 388350
rect 379934 388294 380002 388350
rect 380058 388294 410598 388350
rect 410654 388294 410722 388350
rect 410778 388294 441318 388350
rect 441374 388294 441442 388350
rect 441498 388294 472038 388350
rect 472094 388294 472162 388350
rect 472218 388294 502758 388350
rect 502814 388294 502882 388350
rect 502938 388294 533478 388350
rect 533534 388294 533602 388350
rect 533658 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 39954 388226
rect 40010 388170 40078 388226
rect 40134 388170 40202 388226
rect 40258 388170 40326 388226
rect 40382 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 101394 388226
rect 101450 388170 101518 388226
rect 101574 388170 101642 388226
rect 101698 388170 101766 388226
rect 101822 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 285714 388226
rect 285770 388170 285838 388226
rect 285894 388170 285962 388226
rect 286018 388170 286086 388226
rect 286142 388170 316434 388226
rect 316490 388170 316558 388226
rect 316614 388170 316682 388226
rect 316738 388170 316806 388226
rect 316862 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 379878 388226
rect 379934 388170 380002 388226
rect 380058 388170 410598 388226
rect 410654 388170 410722 388226
rect 410778 388170 441318 388226
rect 441374 388170 441442 388226
rect 441498 388170 472038 388226
rect 472094 388170 472162 388226
rect 472218 388170 502758 388226
rect 502814 388170 502882 388226
rect 502938 388170 533478 388226
rect 533534 388170 533602 388226
rect 533658 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 39954 388102
rect 40010 388046 40078 388102
rect 40134 388046 40202 388102
rect 40258 388046 40326 388102
rect 40382 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 101394 388102
rect 101450 388046 101518 388102
rect 101574 388046 101642 388102
rect 101698 388046 101766 388102
rect 101822 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 285714 388102
rect 285770 388046 285838 388102
rect 285894 388046 285962 388102
rect 286018 388046 286086 388102
rect 286142 388046 316434 388102
rect 316490 388046 316558 388102
rect 316614 388046 316682 388102
rect 316738 388046 316806 388102
rect 316862 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 379878 388102
rect 379934 388046 380002 388102
rect 380058 388046 410598 388102
rect 410654 388046 410722 388102
rect 410778 388046 441318 388102
rect 441374 388046 441442 388102
rect 441498 388046 472038 388102
rect 472094 388046 472162 388102
rect 472218 388046 502758 388102
rect 502814 388046 502882 388102
rect 502938 388046 533478 388102
rect 533534 388046 533602 388102
rect 533658 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 39954 387978
rect 40010 387922 40078 387978
rect 40134 387922 40202 387978
rect 40258 387922 40326 387978
rect 40382 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 101394 387978
rect 101450 387922 101518 387978
rect 101574 387922 101642 387978
rect 101698 387922 101766 387978
rect 101822 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 285714 387978
rect 285770 387922 285838 387978
rect 285894 387922 285962 387978
rect 286018 387922 286086 387978
rect 286142 387922 316434 387978
rect 316490 387922 316558 387978
rect 316614 387922 316682 387978
rect 316738 387922 316806 387978
rect 316862 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 379878 387978
rect 379934 387922 380002 387978
rect 380058 387922 410598 387978
rect 410654 387922 410722 387978
rect 410778 387922 441318 387978
rect 441374 387922 441442 387978
rect 441498 387922 472038 387978
rect 472094 387922 472162 387978
rect 472218 387922 502758 387978
rect 502814 387922 502882 387978
rect 502938 387922 533478 387978
rect 533534 387922 533602 387978
rect 533658 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect 357852 383158 362196 383174
rect 357852 383102 357868 383158
rect 357924 383102 362124 383158
rect 362180 383102 362196 383158
rect 357852 383086 362196 383102
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 281994 382350
rect 282050 382294 282118 382350
rect 282174 382294 282242 382350
rect 282298 382294 282366 382350
rect 282422 382294 312714 382350
rect 312770 382294 312838 382350
rect 312894 382294 312962 382350
rect 313018 382294 313086 382350
rect 313142 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 364518 382350
rect 364574 382294 364642 382350
rect 364698 382294 395238 382350
rect 395294 382294 395362 382350
rect 395418 382294 425958 382350
rect 426014 382294 426082 382350
rect 426138 382294 456678 382350
rect 456734 382294 456802 382350
rect 456858 382294 487398 382350
rect 487454 382294 487522 382350
rect 487578 382294 518118 382350
rect 518174 382294 518242 382350
rect 518298 382294 548838 382350
rect 548894 382294 548962 382350
rect 549018 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 281994 382226
rect 282050 382170 282118 382226
rect 282174 382170 282242 382226
rect 282298 382170 282366 382226
rect 282422 382170 312714 382226
rect 312770 382170 312838 382226
rect 312894 382170 312962 382226
rect 313018 382170 313086 382226
rect 313142 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 364518 382226
rect 364574 382170 364642 382226
rect 364698 382170 395238 382226
rect 395294 382170 395362 382226
rect 395418 382170 425958 382226
rect 426014 382170 426082 382226
rect 426138 382170 456678 382226
rect 456734 382170 456802 382226
rect 456858 382170 487398 382226
rect 487454 382170 487522 382226
rect 487578 382170 518118 382226
rect 518174 382170 518242 382226
rect 518298 382170 548838 382226
rect 548894 382170 548962 382226
rect 549018 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 281994 382102
rect 282050 382046 282118 382102
rect 282174 382046 282242 382102
rect 282298 382046 282366 382102
rect 282422 382046 312714 382102
rect 312770 382046 312838 382102
rect 312894 382046 312962 382102
rect 313018 382046 313086 382102
rect 313142 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 364518 382102
rect 364574 382046 364642 382102
rect 364698 382046 395238 382102
rect 395294 382046 395362 382102
rect 395418 382046 425958 382102
rect 426014 382046 426082 382102
rect 426138 382046 456678 382102
rect 456734 382046 456802 382102
rect 456858 382046 487398 382102
rect 487454 382046 487522 382102
rect 487578 382046 518118 382102
rect 518174 382046 518242 382102
rect 518298 382046 548838 382102
rect 548894 382046 548962 382102
rect 549018 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 281994 381978
rect 282050 381922 282118 381978
rect 282174 381922 282242 381978
rect 282298 381922 282366 381978
rect 282422 381922 312714 381978
rect 312770 381922 312838 381978
rect 312894 381922 312962 381978
rect 313018 381922 313086 381978
rect 313142 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 364518 381978
rect 364574 381922 364642 381978
rect 364698 381922 395238 381978
rect 395294 381922 395362 381978
rect 395418 381922 425958 381978
rect 426014 381922 426082 381978
rect 426138 381922 456678 381978
rect 456734 381922 456802 381978
rect 456858 381922 487398 381978
rect 487454 381922 487522 381978
rect 487578 381922 518118 381978
rect 518174 381922 518242 381978
rect 518298 381922 548838 381978
rect 548894 381922 548962 381978
rect 549018 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect 236108 379738 350324 379754
rect 236108 379682 236124 379738
rect 236180 379682 350252 379738
rect 350308 379682 350324 379738
rect 236108 379666 350324 379682
rect 184476 378838 342932 378854
rect 184476 378782 184492 378838
rect 184548 378782 342860 378838
rect 342916 378782 342932 378838
rect 184476 378766 342932 378782
rect 4156 376318 325964 376334
rect 4156 376262 4172 376318
rect 4228 376262 323372 376318
rect 323428 376262 325964 376318
rect 4156 376246 325964 376262
rect 325876 375434 325964 376246
rect 325876 375418 348644 375434
rect 325876 375362 348572 375418
rect 348628 375362 348644 375418
rect 325876 375346 348644 375362
rect 199372 373798 237092 373814
rect 199372 373742 199388 373798
rect 199444 373742 237020 373798
rect 237076 373742 237092 373798
rect 199372 373726 237092 373742
rect 281356 373798 340356 373814
rect 281356 373742 281372 373798
rect 281428 373742 340284 373798
rect 340340 373742 340356 373798
rect 281356 373726 340356 373742
rect 276316 373078 342148 373094
rect 276316 373022 276332 373078
rect 276388 373022 342076 373078
rect 342132 373022 342148 373078
rect 276316 373006 342148 373022
rect 286396 372178 350660 372194
rect 286396 372122 286412 372178
rect 286468 372122 350588 372178
rect 350644 372122 350660 372178
rect 286396 372106 350660 372122
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 39954 370350
rect 40010 370294 40078 370350
rect 40134 370294 40202 370350
rect 40258 370294 40326 370350
rect 40382 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 101394 370350
rect 101450 370294 101518 370350
rect 101574 370294 101642 370350
rect 101698 370294 101766 370350
rect 101822 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 209878 370350
rect 209934 370294 210002 370350
rect 210058 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 240598 370350
rect 240654 370294 240722 370350
rect 240778 370294 254994 370350
rect 255050 370294 255118 370350
rect 255174 370294 255242 370350
rect 255298 370294 255366 370350
rect 255422 370294 271318 370350
rect 271374 370294 271442 370350
rect 271498 370294 285714 370350
rect 285770 370294 285838 370350
rect 285894 370294 285962 370350
rect 286018 370294 286086 370350
rect 286142 370294 302038 370350
rect 302094 370294 302162 370350
rect 302218 370294 316434 370350
rect 316490 370294 316558 370350
rect 316614 370294 316682 370350
rect 316738 370294 316806 370350
rect 316862 370294 332758 370350
rect 332814 370294 332882 370350
rect 332938 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 379878 370350
rect 379934 370294 380002 370350
rect 380058 370294 410598 370350
rect 410654 370294 410722 370350
rect 410778 370294 441318 370350
rect 441374 370294 441442 370350
rect 441498 370294 472038 370350
rect 472094 370294 472162 370350
rect 472218 370294 502758 370350
rect 502814 370294 502882 370350
rect 502938 370294 533478 370350
rect 533534 370294 533602 370350
rect 533658 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 39954 370226
rect 40010 370170 40078 370226
rect 40134 370170 40202 370226
rect 40258 370170 40326 370226
rect 40382 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 101394 370226
rect 101450 370170 101518 370226
rect 101574 370170 101642 370226
rect 101698 370170 101766 370226
rect 101822 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 209878 370226
rect 209934 370170 210002 370226
rect 210058 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 240598 370226
rect 240654 370170 240722 370226
rect 240778 370170 254994 370226
rect 255050 370170 255118 370226
rect 255174 370170 255242 370226
rect 255298 370170 255366 370226
rect 255422 370170 271318 370226
rect 271374 370170 271442 370226
rect 271498 370170 285714 370226
rect 285770 370170 285838 370226
rect 285894 370170 285962 370226
rect 286018 370170 286086 370226
rect 286142 370170 302038 370226
rect 302094 370170 302162 370226
rect 302218 370170 316434 370226
rect 316490 370170 316558 370226
rect 316614 370170 316682 370226
rect 316738 370170 316806 370226
rect 316862 370170 332758 370226
rect 332814 370170 332882 370226
rect 332938 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 379878 370226
rect 379934 370170 380002 370226
rect 380058 370170 410598 370226
rect 410654 370170 410722 370226
rect 410778 370170 441318 370226
rect 441374 370170 441442 370226
rect 441498 370170 472038 370226
rect 472094 370170 472162 370226
rect 472218 370170 502758 370226
rect 502814 370170 502882 370226
rect 502938 370170 533478 370226
rect 533534 370170 533602 370226
rect 533658 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 39954 370102
rect 40010 370046 40078 370102
rect 40134 370046 40202 370102
rect 40258 370046 40326 370102
rect 40382 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 101394 370102
rect 101450 370046 101518 370102
rect 101574 370046 101642 370102
rect 101698 370046 101766 370102
rect 101822 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 209878 370102
rect 209934 370046 210002 370102
rect 210058 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 240598 370102
rect 240654 370046 240722 370102
rect 240778 370046 254994 370102
rect 255050 370046 255118 370102
rect 255174 370046 255242 370102
rect 255298 370046 255366 370102
rect 255422 370046 271318 370102
rect 271374 370046 271442 370102
rect 271498 370046 285714 370102
rect 285770 370046 285838 370102
rect 285894 370046 285962 370102
rect 286018 370046 286086 370102
rect 286142 370046 302038 370102
rect 302094 370046 302162 370102
rect 302218 370046 316434 370102
rect 316490 370046 316558 370102
rect 316614 370046 316682 370102
rect 316738 370046 316806 370102
rect 316862 370046 332758 370102
rect 332814 370046 332882 370102
rect 332938 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 379878 370102
rect 379934 370046 380002 370102
rect 380058 370046 410598 370102
rect 410654 370046 410722 370102
rect 410778 370046 441318 370102
rect 441374 370046 441442 370102
rect 441498 370046 472038 370102
rect 472094 370046 472162 370102
rect 472218 370046 502758 370102
rect 502814 370046 502882 370102
rect 502938 370046 533478 370102
rect 533534 370046 533602 370102
rect 533658 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 39954 369978
rect 40010 369922 40078 369978
rect 40134 369922 40202 369978
rect 40258 369922 40326 369978
rect 40382 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 101394 369978
rect 101450 369922 101518 369978
rect 101574 369922 101642 369978
rect 101698 369922 101766 369978
rect 101822 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 209878 369978
rect 209934 369922 210002 369978
rect 210058 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 240598 369978
rect 240654 369922 240722 369978
rect 240778 369922 254994 369978
rect 255050 369922 255118 369978
rect 255174 369922 255242 369978
rect 255298 369922 255366 369978
rect 255422 369922 271318 369978
rect 271374 369922 271442 369978
rect 271498 369922 285714 369978
rect 285770 369922 285838 369978
rect 285894 369922 285962 369978
rect 286018 369922 286086 369978
rect 286142 369922 302038 369978
rect 302094 369922 302162 369978
rect 302218 369922 316434 369978
rect 316490 369922 316558 369978
rect 316614 369922 316682 369978
rect 316738 369922 316806 369978
rect 316862 369922 332758 369978
rect 332814 369922 332882 369978
rect 332938 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 379878 369978
rect 379934 369922 380002 369978
rect 380058 369922 410598 369978
rect 410654 369922 410722 369978
rect 410778 369922 441318 369978
rect 441374 369922 441442 369978
rect 441498 369922 472038 369978
rect 472094 369922 472162 369978
rect 472218 369922 502758 369978
rect 502814 369922 502882 369978
rect 502938 369922 533478 369978
rect 533534 369922 533602 369978
rect 533658 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect 329068 369118 357156 369134
rect 329068 369062 329084 369118
rect 329140 369062 357084 369118
rect 357140 369062 357156 369118
rect 329068 369046 357156 369062
rect 266236 368938 337724 368954
rect 266236 368882 266252 368938
rect 266308 368882 337724 368938
rect 266236 368866 337724 368882
rect 337636 368774 337724 368866
rect 199260 368758 235300 368774
rect 199260 368702 199276 368758
rect 199332 368702 235228 368758
rect 235284 368702 235300 368758
rect 199260 368686 235300 368702
rect 238460 368758 336100 368774
rect 238460 368702 238476 368758
rect 238532 368702 336028 368758
rect 336084 368702 336100 368758
rect 238460 368686 336100 368702
rect 337636 368758 354356 368774
rect 337636 368702 338268 368758
rect 338324 368702 354284 368758
rect 354340 368702 354356 368758
rect 337636 368686 354356 368702
rect 93980 367138 276404 367154
rect 93980 367082 93996 367138
rect 94052 367082 276332 367138
rect 276388 367082 276404 367138
rect 93980 367066 276404 367082
rect 272060 366598 355476 366614
rect 272060 366542 272076 366598
rect 272132 366542 355404 366598
rect 355460 366542 355476 366598
rect 272060 366526 355476 366542
rect 63740 366418 344500 366434
rect 63740 366362 63756 366418
rect 63812 366362 344428 366418
rect 344484 366362 344500 366418
rect 63740 366346 344500 366362
rect 78860 365878 272148 365894
rect 78860 365822 78876 365878
rect 78932 365822 270508 365878
rect 270564 365822 272076 365878
rect 272132 365822 272148 365878
rect 78860 365806 272148 365822
rect -1916 364416 597980 364446
rect -1916 364360 159114 364416
rect 159170 364360 159238 364416
rect 159294 364360 159362 364416
rect 159418 364360 159486 364416
rect 159542 364360 597980 364416
rect -1916 364350 597980 364360
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 194518 364350
rect 194574 364294 194642 364350
rect 194698 364294 225238 364350
rect 225294 364294 225362 364350
rect 225418 364294 255958 364350
rect 256014 364294 256082 364350
rect 256138 364294 286678 364350
rect 286734 364294 286802 364350
rect 286858 364294 317398 364350
rect 317454 364294 317522 364350
rect 317578 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 364518 364350
rect 364574 364294 364642 364350
rect 364698 364294 395238 364350
rect 395294 364294 395362 364350
rect 395418 364294 425958 364350
rect 426014 364294 426082 364350
rect 426138 364294 456678 364350
rect 456734 364294 456802 364350
rect 456858 364294 487398 364350
rect 487454 364294 487522 364350
rect 487578 364294 518118 364350
rect 518174 364294 518242 364350
rect 518298 364294 548838 364350
rect 548894 364294 548962 364350
rect 549018 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364292 597980 364294
rect -1916 364236 159114 364292
rect 159170 364236 159238 364292
rect 159294 364236 159362 364292
rect 159418 364236 159486 364292
rect 159542 364236 597980 364292
rect -1916 364226 597980 364236
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 194518 364226
rect 194574 364170 194642 364226
rect 194698 364170 225238 364226
rect 225294 364170 225362 364226
rect 225418 364170 255958 364226
rect 256014 364170 256082 364226
rect 256138 364170 286678 364226
rect 286734 364170 286802 364226
rect 286858 364170 317398 364226
rect 317454 364170 317522 364226
rect 317578 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 364518 364226
rect 364574 364170 364642 364226
rect 364698 364170 395238 364226
rect 395294 364170 395362 364226
rect 395418 364170 425958 364226
rect 426014 364170 426082 364226
rect 426138 364170 456678 364226
rect 456734 364170 456802 364226
rect 456858 364170 487398 364226
rect 487454 364170 487522 364226
rect 487578 364170 518118 364226
rect 518174 364170 518242 364226
rect 518298 364170 548838 364226
rect 548894 364170 548962 364226
rect 549018 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 194518 364102
rect 194574 364046 194642 364102
rect 194698 364046 225238 364102
rect 225294 364046 225362 364102
rect 225418 364046 255958 364102
rect 256014 364046 256082 364102
rect 256138 364046 286678 364102
rect 286734 364046 286802 364102
rect 286858 364046 317398 364102
rect 317454 364046 317522 364102
rect 317578 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 364518 364102
rect 364574 364046 364642 364102
rect 364698 364046 395238 364102
rect 395294 364046 395362 364102
rect 395418 364046 425958 364102
rect 426014 364046 426082 364102
rect 426138 364046 456678 364102
rect 456734 364046 456802 364102
rect 456858 364046 487398 364102
rect 487454 364046 487522 364102
rect 487578 364046 518118 364102
rect 518174 364046 518242 364102
rect 518298 364046 548838 364102
rect 548894 364046 548962 364102
rect 549018 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 194518 363978
rect 194574 363922 194642 363978
rect 194698 363922 225238 363978
rect 225294 363922 225362 363978
rect 225418 363922 255958 363978
rect 256014 363922 256082 363978
rect 256138 363922 286678 363978
rect 286734 363922 286802 363978
rect 286858 363922 317398 363978
rect 317454 363922 317522 363978
rect 317578 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 364518 363978
rect 364574 363922 364642 363978
rect 364698 363922 395238 363978
rect 395294 363922 395362 363978
rect 395418 363922 425958 363978
rect 426014 363922 426082 363978
rect 426138 363922 456678 363978
rect 456734 363922 456802 363978
rect 456858 363922 487398 363978
rect 487454 363922 487522 363978
rect 487578 363922 518118 363978
rect 518174 363922 518242 363978
rect 518298 363922 548838 363978
rect 548894 363922 548962 363978
rect 549018 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect 335900 356158 356596 356174
rect 335900 356102 335916 356158
rect 335972 356102 356524 356158
rect 356580 356102 356596 356158
rect 335900 356086 356596 356102
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 39954 352350
rect 40010 352294 40078 352350
rect 40134 352294 40202 352350
rect 40258 352294 40326 352350
rect 40382 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 101394 352350
rect 101450 352294 101518 352350
rect 101574 352294 101642 352350
rect 101698 352294 101766 352350
rect 101822 352294 132114 352350
rect 132170 352294 132238 352350
rect 132294 352294 132362 352350
rect 132418 352294 132486 352350
rect 132542 352294 149878 352350
rect 149934 352294 150002 352350
rect 150058 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 209878 352350
rect 209934 352294 210002 352350
rect 210058 352294 240598 352350
rect 240654 352294 240722 352350
rect 240778 352294 271318 352350
rect 271374 352294 271442 352350
rect 271498 352294 302038 352350
rect 302094 352294 302162 352350
rect 302218 352294 332758 352350
rect 332814 352294 332882 352350
rect 332938 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 379878 352350
rect 379934 352294 380002 352350
rect 380058 352294 410598 352350
rect 410654 352294 410722 352350
rect 410778 352294 441318 352350
rect 441374 352294 441442 352350
rect 441498 352294 472038 352350
rect 472094 352294 472162 352350
rect 472218 352294 502758 352350
rect 502814 352294 502882 352350
rect 502938 352294 533478 352350
rect 533534 352294 533602 352350
rect 533658 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 39954 352226
rect 40010 352170 40078 352226
rect 40134 352170 40202 352226
rect 40258 352170 40326 352226
rect 40382 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 101394 352226
rect 101450 352170 101518 352226
rect 101574 352170 101642 352226
rect 101698 352170 101766 352226
rect 101822 352170 132114 352226
rect 132170 352170 132238 352226
rect 132294 352170 132362 352226
rect 132418 352170 132486 352226
rect 132542 352170 149878 352226
rect 149934 352170 150002 352226
rect 150058 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 209878 352226
rect 209934 352170 210002 352226
rect 210058 352170 240598 352226
rect 240654 352170 240722 352226
rect 240778 352170 271318 352226
rect 271374 352170 271442 352226
rect 271498 352170 302038 352226
rect 302094 352170 302162 352226
rect 302218 352170 332758 352226
rect 332814 352170 332882 352226
rect 332938 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 379878 352226
rect 379934 352170 380002 352226
rect 380058 352170 410598 352226
rect 410654 352170 410722 352226
rect 410778 352170 441318 352226
rect 441374 352170 441442 352226
rect 441498 352170 472038 352226
rect 472094 352170 472162 352226
rect 472218 352170 502758 352226
rect 502814 352170 502882 352226
rect 502938 352170 533478 352226
rect 533534 352170 533602 352226
rect 533658 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 39954 352102
rect 40010 352046 40078 352102
rect 40134 352046 40202 352102
rect 40258 352046 40326 352102
rect 40382 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 101394 352102
rect 101450 352046 101518 352102
rect 101574 352046 101642 352102
rect 101698 352046 101766 352102
rect 101822 352046 132114 352102
rect 132170 352046 132238 352102
rect 132294 352046 132362 352102
rect 132418 352046 132486 352102
rect 132542 352046 149878 352102
rect 149934 352046 150002 352102
rect 150058 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 209878 352102
rect 209934 352046 210002 352102
rect 210058 352046 240598 352102
rect 240654 352046 240722 352102
rect 240778 352046 271318 352102
rect 271374 352046 271442 352102
rect 271498 352046 302038 352102
rect 302094 352046 302162 352102
rect 302218 352046 332758 352102
rect 332814 352046 332882 352102
rect 332938 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 379878 352102
rect 379934 352046 380002 352102
rect 380058 352046 410598 352102
rect 410654 352046 410722 352102
rect 410778 352046 441318 352102
rect 441374 352046 441442 352102
rect 441498 352046 472038 352102
rect 472094 352046 472162 352102
rect 472218 352046 502758 352102
rect 502814 352046 502882 352102
rect 502938 352046 533478 352102
rect 533534 352046 533602 352102
rect 533658 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 39954 351978
rect 40010 351922 40078 351978
rect 40134 351922 40202 351978
rect 40258 351922 40326 351978
rect 40382 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 101394 351978
rect 101450 351922 101518 351978
rect 101574 351922 101642 351978
rect 101698 351922 101766 351978
rect 101822 351922 132114 351978
rect 132170 351922 132238 351978
rect 132294 351922 132362 351978
rect 132418 351922 132486 351978
rect 132542 351922 149878 351978
rect 149934 351922 150002 351978
rect 150058 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 209878 351978
rect 209934 351922 210002 351978
rect 210058 351922 240598 351978
rect 240654 351922 240722 351978
rect 240778 351922 271318 351978
rect 271374 351922 271442 351978
rect 271498 351922 302038 351978
rect 302094 351922 302162 351978
rect 302218 351922 332758 351978
rect 332814 351922 332882 351978
rect 332938 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 379878 351978
rect 379934 351922 380002 351978
rect 380058 351922 410598 351978
rect 410654 351922 410722 351978
rect 410778 351922 441318 351978
rect 441374 351922 441442 351978
rect 441498 351922 472038 351978
rect 472094 351922 472162 351978
rect 472218 351922 502758 351978
rect 502814 351922 502882 351978
rect 502938 351922 533478 351978
rect 533534 351922 533602 351978
rect 533658 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 134518 346350
rect 134574 346294 134642 346350
rect 134698 346294 165238 346350
rect 165294 346294 165362 346350
rect 165418 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 194518 346350
rect 194574 346294 194642 346350
rect 194698 346294 225238 346350
rect 225294 346294 225362 346350
rect 225418 346294 255958 346350
rect 256014 346294 256082 346350
rect 256138 346294 286678 346350
rect 286734 346294 286802 346350
rect 286858 346294 317398 346350
rect 317454 346294 317522 346350
rect 317578 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 364518 346350
rect 364574 346294 364642 346350
rect 364698 346294 395238 346350
rect 395294 346294 395362 346350
rect 395418 346294 425958 346350
rect 426014 346294 426082 346350
rect 426138 346294 456678 346350
rect 456734 346294 456802 346350
rect 456858 346294 487398 346350
rect 487454 346294 487522 346350
rect 487578 346294 518118 346350
rect 518174 346294 518242 346350
rect 518298 346294 548838 346350
rect 548894 346294 548962 346350
rect 549018 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 134518 346226
rect 134574 346170 134642 346226
rect 134698 346170 165238 346226
rect 165294 346170 165362 346226
rect 165418 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 194518 346226
rect 194574 346170 194642 346226
rect 194698 346170 225238 346226
rect 225294 346170 225362 346226
rect 225418 346170 255958 346226
rect 256014 346170 256082 346226
rect 256138 346170 286678 346226
rect 286734 346170 286802 346226
rect 286858 346170 317398 346226
rect 317454 346170 317522 346226
rect 317578 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 364518 346226
rect 364574 346170 364642 346226
rect 364698 346170 395238 346226
rect 395294 346170 395362 346226
rect 395418 346170 425958 346226
rect 426014 346170 426082 346226
rect 426138 346170 456678 346226
rect 456734 346170 456802 346226
rect 456858 346170 487398 346226
rect 487454 346170 487522 346226
rect 487578 346170 518118 346226
rect 518174 346170 518242 346226
rect 518298 346170 548838 346226
rect 548894 346170 548962 346226
rect 549018 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 134518 346102
rect 134574 346046 134642 346102
rect 134698 346046 165238 346102
rect 165294 346046 165362 346102
rect 165418 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 194518 346102
rect 194574 346046 194642 346102
rect 194698 346046 225238 346102
rect 225294 346046 225362 346102
rect 225418 346046 255958 346102
rect 256014 346046 256082 346102
rect 256138 346046 286678 346102
rect 286734 346046 286802 346102
rect 286858 346046 317398 346102
rect 317454 346046 317522 346102
rect 317578 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 364518 346102
rect 364574 346046 364642 346102
rect 364698 346046 395238 346102
rect 395294 346046 395362 346102
rect 395418 346046 425958 346102
rect 426014 346046 426082 346102
rect 426138 346046 456678 346102
rect 456734 346046 456802 346102
rect 456858 346046 487398 346102
rect 487454 346046 487522 346102
rect 487578 346046 518118 346102
rect 518174 346046 518242 346102
rect 518298 346046 548838 346102
rect 548894 346046 548962 346102
rect 549018 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 134518 345978
rect 134574 345922 134642 345978
rect 134698 345922 165238 345978
rect 165294 345922 165362 345978
rect 165418 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 194518 345978
rect 194574 345922 194642 345978
rect 194698 345922 225238 345978
rect 225294 345922 225362 345978
rect 225418 345922 255958 345978
rect 256014 345922 256082 345978
rect 256138 345922 286678 345978
rect 286734 345922 286802 345978
rect 286858 345922 317398 345978
rect 317454 345922 317522 345978
rect 317578 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 364518 345978
rect 364574 345922 364642 345978
rect 364698 345922 395238 345978
rect 395294 345922 395362 345978
rect 395418 345922 425958 345978
rect 426014 345922 426082 345978
rect 426138 345922 456678 345978
rect 456734 345922 456802 345978
rect 456858 345922 487398 345978
rect 487454 345922 487522 345978
rect 487578 345922 518118 345978
rect 518174 345922 518242 345978
rect 518298 345922 548838 345978
rect 548894 345922 548962 345978
rect 549018 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect 178092 340138 197668 340154
rect 178092 340082 178108 340138
rect 178164 340082 197596 340138
rect 197652 340082 197668 340138
rect 178092 340066 197668 340082
rect 338140 336358 339460 336374
rect 338140 336302 338156 336358
rect 338212 336302 339388 336358
rect 339444 336302 339460 336358
rect 338140 336286 339460 336302
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 39954 334350
rect 40010 334294 40078 334350
rect 40134 334294 40202 334350
rect 40258 334294 40326 334350
rect 40382 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 101394 334350
rect 101450 334294 101518 334350
rect 101574 334294 101642 334350
rect 101698 334294 101766 334350
rect 101822 334294 132114 334350
rect 132170 334294 132238 334350
rect 132294 334294 132362 334350
rect 132418 334294 132486 334350
rect 132542 334294 149878 334350
rect 149934 334294 150002 334350
rect 150058 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 209878 334350
rect 209934 334294 210002 334350
rect 210058 334294 240598 334350
rect 240654 334294 240722 334350
rect 240778 334294 271318 334350
rect 271374 334294 271442 334350
rect 271498 334294 302038 334350
rect 302094 334294 302162 334350
rect 302218 334294 332758 334350
rect 332814 334294 332882 334350
rect 332938 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 379878 334350
rect 379934 334294 380002 334350
rect 380058 334294 410598 334350
rect 410654 334294 410722 334350
rect 410778 334294 441318 334350
rect 441374 334294 441442 334350
rect 441498 334294 472038 334350
rect 472094 334294 472162 334350
rect 472218 334294 502758 334350
rect 502814 334294 502882 334350
rect 502938 334294 533478 334350
rect 533534 334294 533602 334350
rect 533658 334294 562194 334350
rect 562250 334294 562318 334350
rect 562374 334294 562442 334350
rect 562498 334294 562566 334350
rect 562622 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 39954 334226
rect 40010 334170 40078 334226
rect 40134 334170 40202 334226
rect 40258 334170 40326 334226
rect 40382 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 101394 334226
rect 101450 334170 101518 334226
rect 101574 334170 101642 334226
rect 101698 334170 101766 334226
rect 101822 334170 132114 334226
rect 132170 334170 132238 334226
rect 132294 334170 132362 334226
rect 132418 334170 132486 334226
rect 132542 334170 149878 334226
rect 149934 334170 150002 334226
rect 150058 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 209878 334226
rect 209934 334170 210002 334226
rect 210058 334170 240598 334226
rect 240654 334170 240722 334226
rect 240778 334170 271318 334226
rect 271374 334170 271442 334226
rect 271498 334170 302038 334226
rect 302094 334170 302162 334226
rect 302218 334170 332758 334226
rect 332814 334170 332882 334226
rect 332938 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 379878 334226
rect 379934 334170 380002 334226
rect 380058 334170 410598 334226
rect 410654 334170 410722 334226
rect 410778 334170 441318 334226
rect 441374 334170 441442 334226
rect 441498 334170 472038 334226
rect 472094 334170 472162 334226
rect 472218 334170 502758 334226
rect 502814 334170 502882 334226
rect 502938 334170 533478 334226
rect 533534 334170 533602 334226
rect 533658 334170 562194 334226
rect 562250 334170 562318 334226
rect 562374 334170 562442 334226
rect 562498 334170 562566 334226
rect 562622 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 39954 334102
rect 40010 334046 40078 334102
rect 40134 334046 40202 334102
rect 40258 334046 40326 334102
rect 40382 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 101394 334102
rect 101450 334046 101518 334102
rect 101574 334046 101642 334102
rect 101698 334046 101766 334102
rect 101822 334046 132114 334102
rect 132170 334046 132238 334102
rect 132294 334046 132362 334102
rect 132418 334046 132486 334102
rect 132542 334046 149878 334102
rect 149934 334046 150002 334102
rect 150058 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 209878 334102
rect 209934 334046 210002 334102
rect 210058 334046 240598 334102
rect 240654 334046 240722 334102
rect 240778 334046 271318 334102
rect 271374 334046 271442 334102
rect 271498 334046 302038 334102
rect 302094 334046 302162 334102
rect 302218 334046 332758 334102
rect 332814 334046 332882 334102
rect 332938 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 379878 334102
rect 379934 334046 380002 334102
rect 380058 334046 410598 334102
rect 410654 334046 410722 334102
rect 410778 334046 441318 334102
rect 441374 334046 441442 334102
rect 441498 334046 472038 334102
rect 472094 334046 472162 334102
rect 472218 334046 502758 334102
rect 502814 334046 502882 334102
rect 502938 334046 533478 334102
rect 533534 334046 533602 334102
rect 533658 334046 562194 334102
rect 562250 334046 562318 334102
rect 562374 334046 562442 334102
rect 562498 334046 562566 334102
rect 562622 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 39954 333978
rect 40010 333922 40078 333978
rect 40134 333922 40202 333978
rect 40258 333922 40326 333978
rect 40382 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 101394 333978
rect 101450 333922 101518 333978
rect 101574 333922 101642 333978
rect 101698 333922 101766 333978
rect 101822 333922 132114 333978
rect 132170 333922 132238 333978
rect 132294 333922 132362 333978
rect 132418 333922 132486 333978
rect 132542 333922 149878 333978
rect 149934 333922 150002 333978
rect 150058 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 209878 333978
rect 209934 333922 210002 333978
rect 210058 333922 240598 333978
rect 240654 333922 240722 333978
rect 240778 333922 271318 333978
rect 271374 333922 271442 333978
rect 271498 333922 302038 333978
rect 302094 333922 302162 333978
rect 302218 333922 332758 333978
rect 332814 333922 332882 333978
rect 332938 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 379878 333978
rect 379934 333922 380002 333978
rect 380058 333922 410598 333978
rect 410654 333922 410722 333978
rect 410778 333922 441318 333978
rect 441374 333922 441442 333978
rect 441498 333922 472038 333978
rect 472094 333922 472162 333978
rect 472218 333922 502758 333978
rect 502814 333922 502882 333978
rect 502938 333922 533478 333978
rect 533534 333922 533602 333978
rect 533658 333922 562194 333978
rect 562250 333922 562318 333978
rect 562374 333922 562442 333978
rect 562498 333922 562566 333978
rect 562622 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 134518 328350
rect 134574 328294 134642 328350
rect 134698 328294 165238 328350
rect 165294 328294 165362 328350
rect 165418 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 194518 328350
rect 194574 328294 194642 328350
rect 194698 328294 225238 328350
rect 225294 328294 225362 328350
rect 225418 328294 255958 328350
rect 256014 328294 256082 328350
rect 256138 328294 286678 328350
rect 286734 328294 286802 328350
rect 286858 328294 317398 328350
rect 317454 328294 317522 328350
rect 317578 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 364518 328350
rect 364574 328294 364642 328350
rect 364698 328294 395238 328350
rect 395294 328294 395362 328350
rect 395418 328294 425958 328350
rect 426014 328294 426082 328350
rect 426138 328294 456678 328350
rect 456734 328294 456802 328350
rect 456858 328294 487398 328350
rect 487454 328294 487522 328350
rect 487578 328294 518118 328350
rect 518174 328294 518242 328350
rect 518298 328294 548838 328350
rect 548894 328294 548962 328350
rect 549018 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 134518 328226
rect 134574 328170 134642 328226
rect 134698 328170 165238 328226
rect 165294 328170 165362 328226
rect 165418 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 194518 328226
rect 194574 328170 194642 328226
rect 194698 328170 225238 328226
rect 225294 328170 225362 328226
rect 225418 328170 255958 328226
rect 256014 328170 256082 328226
rect 256138 328170 286678 328226
rect 286734 328170 286802 328226
rect 286858 328170 317398 328226
rect 317454 328170 317522 328226
rect 317578 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 364518 328226
rect 364574 328170 364642 328226
rect 364698 328170 395238 328226
rect 395294 328170 395362 328226
rect 395418 328170 425958 328226
rect 426014 328170 426082 328226
rect 426138 328170 456678 328226
rect 456734 328170 456802 328226
rect 456858 328170 487398 328226
rect 487454 328170 487522 328226
rect 487578 328170 518118 328226
rect 518174 328170 518242 328226
rect 518298 328170 548838 328226
rect 548894 328170 548962 328226
rect 549018 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 134518 328102
rect 134574 328046 134642 328102
rect 134698 328046 165238 328102
rect 165294 328046 165362 328102
rect 165418 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 194518 328102
rect 194574 328046 194642 328102
rect 194698 328046 225238 328102
rect 225294 328046 225362 328102
rect 225418 328046 255958 328102
rect 256014 328046 256082 328102
rect 256138 328046 286678 328102
rect 286734 328046 286802 328102
rect 286858 328046 317398 328102
rect 317454 328046 317522 328102
rect 317578 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 364518 328102
rect 364574 328046 364642 328102
rect 364698 328046 395238 328102
rect 395294 328046 395362 328102
rect 395418 328046 425958 328102
rect 426014 328046 426082 328102
rect 426138 328046 456678 328102
rect 456734 328046 456802 328102
rect 456858 328046 487398 328102
rect 487454 328046 487522 328102
rect 487578 328046 518118 328102
rect 518174 328046 518242 328102
rect 518298 328046 548838 328102
rect 548894 328046 548962 328102
rect 549018 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 134518 327978
rect 134574 327922 134642 327978
rect 134698 327922 165238 327978
rect 165294 327922 165362 327978
rect 165418 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 194518 327978
rect 194574 327922 194642 327978
rect 194698 327922 225238 327978
rect 225294 327922 225362 327978
rect 225418 327922 255958 327978
rect 256014 327922 256082 327978
rect 256138 327922 286678 327978
rect 286734 327922 286802 327978
rect 286858 327922 317398 327978
rect 317454 327922 317522 327978
rect 317578 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 364518 327978
rect 364574 327922 364642 327978
rect 364698 327922 395238 327978
rect 395294 327922 395362 327978
rect 395418 327922 425958 327978
rect 426014 327922 426082 327978
rect 426138 327922 456678 327978
rect 456734 327922 456802 327978
rect 456858 327922 487398 327978
rect 487454 327922 487522 327978
rect 487578 327922 518118 327978
rect 518174 327922 518242 327978
rect 518298 327922 548838 327978
rect 548894 327922 548962 327978
rect 549018 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect 342284 325918 356260 325934
rect 342284 325862 342300 325918
rect 342356 325862 356188 325918
rect 356244 325862 356260 325918
rect 342284 325846 356260 325862
rect 190636 323398 192404 323414
rect 190636 323342 190652 323398
rect 190708 323342 192332 323398
rect 192388 323342 192404 323398
rect 190636 323326 192404 323342
rect 172156 322678 187476 322694
rect 172156 322622 172172 322678
rect 172228 322622 187404 322678
rect 187460 322622 187476 322678
rect 172156 322606 187476 322622
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 39954 316350
rect 40010 316294 40078 316350
rect 40134 316294 40202 316350
rect 40258 316294 40326 316350
rect 40382 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 101394 316350
rect 101450 316294 101518 316350
rect 101574 316294 101642 316350
rect 101698 316294 101766 316350
rect 101822 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 209878 316350
rect 209934 316294 210002 316350
rect 210058 316294 240598 316350
rect 240654 316294 240722 316350
rect 240778 316294 271318 316350
rect 271374 316294 271442 316350
rect 271498 316294 302038 316350
rect 302094 316294 302162 316350
rect 302218 316294 332758 316350
rect 332814 316294 332882 316350
rect 332938 316294 347154 316350
rect 347210 316294 347278 316350
rect 347334 316294 347402 316350
rect 347458 316294 347526 316350
rect 347582 316294 379878 316350
rect 379934 316294 380002 316350
rect 380058 316294 410598 316350
rect 410654 316294 410722 316350
rect 410778 316294 441318 316350
rect 441374 316294 441442 316350
rect 441498 316294 472038 316350
rect 472094 316294 472162 316350
rect 472218 316294 502758 316350
rect 502814 316294 502882 316350
rect 502938 316294 533478 316350
rect 533534 316294 533602 316350
rect 533658 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 39954 316226
rect 40010 316170 40078 316226
rect 40134 316170 40202 316226
rect 40258 316170 40326 316226
rect 40382 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 101394 316226
rect 101450 316170 101518 316226
rect 101574 316170 101642 316226
rect 101698 316170 101766 316226
rect 101822 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 209878 316226
rect 209934 316170 210002 316226
rect 210058 316170 240598 316226
rect 240654 316170 240722 316226
rect 240778 316170 271318 316226
rect 271374 316170 271442 316226
rect 271498 316170 302038 316226
rect 302094 316170 302162 316226
rect 302218 316170 332758 316226
rect 332814 316170 332882 316226
rect 332938 316170 347154 316226
rect 347210 316170 347278 316226
rect 347334 316170 347402 316226
rect 347458 316170 347526 316226
rect 347582 316170 379878 316226
rect 379934 316170 380002 316226
rect 380058 316170 410598 316226
rect 410654 316170 410722 316226
rect 410778 316170 441318 316226
rect 441374 316170 441442 316226
rect 441498 316170 472038 316226
rect 472094 316170 472162 316226
rect 472218 316170 502758 316226
rect 502814 316170 502882 316226
rect 502938 316170 533478 316226
rect 533534 316170 533602 316226
rect 533658 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 39954 316102
rect 40010 316046 40078 316102
rect 40134 316046 40202 316102
rect 40258 316046 40326 316102
rect 40382 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 101394 316102
rect 101450 316046 101518 316102
rect 101574 316046 101642 316102
rect 101698 316046 101766 316102
rect 101822 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 209878 316102
rect 209934 316046 210002 316102
rect 210058 316046 240598 316102
rect 240654 316046 240722 316102
rect 240778 316046 271318 316102
rect 271374 316046 271442 316102
rect 271498 316046 302038 316102
rect 302094 316046 302162 316102
rect 302218 316046 332758 316102
rect 332814 316046 332882 316102
rect 332938 316046 347154 316102
rect 347210 316046 347278 316102
rect 347334 316046 347402 316102
rect 347458 316046 347526 316102
rect 347582 316046 379878 316102
rect 379934 316046 380002 316102
rect 380058 316046 410598 316102
rect 410654 316046 410722 316102
rect 410778 316046 441318 316102
rect 441374 316046 441442 316102
rect 441498 316046 472038 316102
rect 472094 316046 472162 316102
rect 472218 316046 502758 316102
rect 502814 316046 502882 316102
rect 502938 316046 533478 316102
rect 533534 316046 533602 316102
rect 533658 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 39954 315978
rect 40010 315922 40078 315978
rect 40134 315922 40202 315978
rect 40258 315922 40326 315978
rect 40382 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 101394 315978
rect 101450 315922 101518 315978
rect 101574 315922 101642 315978
rect 101698 315922 101766 315978
rect 101822 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 209878 315978
rect 209934 315922 210002 315978
rect 210058 315922 240598 315978
rect 240654 315922 240722 315978
rect 240778 315922 271318 315978
rect 271374 315922 271442 315978
rect 271498 315922 302038 315978
rect 302094 315922 302162 315978
rect 302218 315922 332758 315978
rect 332814 315922 332882 315978
rect 332938 315922 347154 315978
rect 347210 315922 347278 315978
rect 347334 315922 347402 315978
rect 347458 315922 347526 315978
rect 347582 315922 379878 315978
rect 379934 315922 380002 315978
rect 380058 315922 410598 315978
rect 410654 315922 410722 315978
rect 410778 315922 441318 315978
rect 441374 315922 441442 315978
rect 441498 315922 472038 315978
rect 472094 315922 472162 315978
rect 472218 315922 502758 315978
rect 502814 315922 502882 315978
rect 502938 315922 533478 315978
rect 533534 315922 533602 315978
rect 533658 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect 338812 313318 339460 313334
rect 338812 313262 338828 313318
rect 338884 313262 339388 313318
rect 339444 313262 339460 313318
rect 338812 313246 339460 313262
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 194518 310350
rect 194574 310294 194642 310350
rect 194698 310294 225238 310350
rect 225294 310294 225362 310350
rect 225418 310294 255958 310350
rect 256014 310294 256082 310350
rect 256138 310294 286678 310350
rect 286734 310294 286802 310350
rect 286858 310294 317398 310350
rect 317454 310294 317522 310350
rect 317578 310294 343434 310350
rect 343490 310294 343558 310350
rect 343614 310294 343682 310350
rect 343738 310294 343806 310350
rect 343862 310294 364518 310350
rect 364574 310294 364642 310350
rect 364698 310294 395238 310350
rect 395294 310294 395362 310350
rect 395418 310294 425958 310350
rect 426014 310294 426082 310350
rect 426138 310294 456678 310350
rect 456734 310294 456802 310350
rect 456858 310294 487398 310350
rect 487454 310294 487522 310350
rect 487578 310294 518118 310350
rect 518174 310294 518242 310350
rect 518298 310294 548838 310350
rect 548894 310294 548962 310350
rect 549018 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 194518 310226
rect 194574 310170 194642 310226
rect 194698 310170 225238 310226
rect 225294 310170 225362 310226
rect 225418 310170 255958 310226
rect 256014 310170 256082 310226
rect 256138 310170 286678 310226
rect 286734 310170 286802 310226
rect 286858 310170 317398 310226
rect 317454 310170 317522 310226
rect 317578 310170 343434 310226
rect 343490 310170 343558 310226
rect 343614 310170 343682 310226
rect 343738 310170 343806 310226
rect 343862 310170 364518 310226
rect 364574 310170 364642 310226
rect 364698 310170 395238 310226
rect 395294 310170 395362 310226
rect 395418 310170 425958 310226
rect 426014 310170 426082 310226
rect 426138 310170 456678 310226
rect 456734 310170 456802 310226
rect 456858 310170 487398 310226
rect 487454 310170 487522 310226
rect 487578 310170 518118 310226
rect 518174 310170 518242 310226
rect 518298 310170 548838 310226
rect 548894 310170 548962 310226
rect 549018 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 194518 310102
rect 194574 310046 194642 310102
rect 194698 310046 225238 310102
rect 225294 310046 225362 310102
rect 225418 310046 255958 310102
rect 256014 310046 256082 310102
rect 256138 310046 286678 310102
rect 286734 310046 286802 310102
rect 286858 310046 317398 310102
rect 317454 310046 317522 310102
rect 317578 310046 343434 310102
rect 343490 310046 343558 310102
rect 343614 310046 343682 310102
rect 343738 310046 343806 310102
rect 343862 310046 364518 310102
rect 364574 310046 364642 310102
rect 364698 310046 395238 310102
rect 395294 310046 395362 310102
rect 395418 310046 425958 310102
rect 426014 310046 426082 310102
rect 426138 310046 456678 310102
rect 456734 310046 456802 310102
rect 456858 310046 487398 310102
rect 487454 310046 487522 310102
rect 487578 310046 518118 310102
rect 518174 310046 518242 310102
rect 518298 310046 548838 310102
rect 548894 310046 548962 310102
rect 549018 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 194518 309978
rect 194574 309922 194642 309978
rect 194698 309922 225238 309978
rect 225294 309922 225362 309978
rect 225418 309922 255958 309978
rect 256014 309922 256082 309978
rect 256138 309922 286678 309978
rect 286734 309922 286802 309978
rect 286858 309922 317398 309978
rect 317454 309922 317522 309978
rect 317578 309922 343434 309978
rect 343490 309922 343558 309978
rect 343614 309922 343682 309978
rect 343738 309922 343806 309978
rect 343862 309922 364518 309978
rect 364574 309922 364642 309978
rect 364698 309922 395238 309978
rect 395294 309922 395362 309978
rect 395418 309922 425958 309978
rect 426014 309922 426082 309978
rect 426138 309922 456678 309978
rect 456734 309922 456802 309978
rect 456858 309922 487398 309978
rect 487454 309922 487522 309978
rect 487578 309922 518118 309978
rect 518174 309922 518242 309978
rect 518298 309922 548838 309978
rect 548894 309922 548962 309978
rect 549018 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect 336908 308998 357380 309014
rect 336908 308942 336924 308998
rect 336980 308942 357308 308998
rect 357364 308942 357380 308998
rect 336908 308926 357380 308942
rect 359868 308638 359956 308654
rect 359868 308582 359884 308638
rect 359940 308582 359956 308638
rect 359868 308294 359956 308582
rect 360092 308638 360188 308654
rect 360092 308582 360108 308638
rect 360164 308582 360188 308638
rect 360092 308566 360188 308582
rect 360092 308458 360180 308566
rect 360092 308402 360108 308458
rect 360164 308402 360180 308458
rect 360092 308386 360180 308402
rect 359868 308278 360404 308294
rect 359868 308222 360332 308278
rect 360388 308222 360404 308278
rect 359868 308206 360404 308222
rect 337636 305038 339348 305054
rect 337636 304982 339276 305038
rect 339332 304982 339348 305038
rect 337636 304966 339348 304982
rect 337636 304874 337724 304966
rect 336684 304858 337724 304874
rect 336684 304802 336700 304858
rect 336756 304802 337724 304858
rect 336684 304786 337724 304802
rect -1916 298422 597980 298446
rect -1916 298366 70674 298422
rect 70730 298366 70798 298422
rect 70854 298366 70922 298422
rect 70978 298366 71046 298422
rect 71102 298366 597980 298422
rect -1916 298350 597980 298366
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 39954 298350
rect 40010 298294 40078 298350
rect 40134 298294 40202 298350
rect 40258 298294 40326 298350
rect 40382 298298 101394 298350
rect 40382 298294 70674 298298
rect -1916 298242 70674 298294
rect 70730 298242 70798 298298
rect 70854 298242 70922 298298
rect 70978 298242 71046 298298
rect 71102 298294 101394 298298
rect 101450 298294 101518 298350
rect 101574 298294 101642 298350
rect 101698 298294 101766 298350
rect 101822 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 209878 298350
rect 209934 298294 210002 298350
rect 210058 298294 240598 298350
rect 240654 298294 240722 298350
rect 240778 298294 271318 298350
rect 271374 298294 271442 298350
rect 271498 298294 302038 298350
rect 302094 298294 302162 298350
rect 302218 298294 332758 298350
rect 332814 298294 332882 298350
rect 332938 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 379878 298350
rect 379934 298294 380002 298350
rect 380058 298294 410598 298350
rect 410654 298294 410722 298350
rect 410778 298294 441318 298350
rect 441374 298294 441442 298350
rect 441498 298294 472038 298350
rect 472094 298294 472162 298350
rect 472218 298294 502758 298350
rect 502814 298294 502882 298350
rect 502938 298294 533478 298350
rect 533534 298294 533602 298350
rect 533658 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 71102 298242 597980 298294
rect -1916 298226 597980 298242
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 39954 298226
rect 40010 298170 40078 298226
rect 40134 298170 40202 298226
rect 40258 298170 40326 298226
rect 40382 298174 101394 298226
rect 40382 298170 70674 298174
rect -1916 298118 70674 298170
rect 70730 298118 70798 298174
rect 70854 298118 70922 298174
rect 70978 298118 71046 298174
rect 71102 298170 101394 298174
rect 101450 298170 101518 298226
rect 101574 298170 101642 298226
rect 101698 298170 101766 298226
rect 101822 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 209878 298226
rect 209934 298170 210002 298226
rect 210058 298170 240598 298226
rect 240654 298170 240722 298226
rect 240778 298170 271318 298226
rect 271374 298170 271442 298226
rect 271498 298170 302038 298226
rect 302094 298170 302162 298226
rect 302218 298170 332758 298226
rect 332814 298170 332882 298226
rect 332938 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 379878 298226
rect 379934 298170 380002 298226
rect 380058 298170 410598 298226
rect 410654 298170 410722 298226
rect 410778 298170 441318 298226
rect 441374 298170 441442 298226
rect 441498 298170 472038 298226
rect 472094 298170 472162 298226
rect 472218 298170 502758 298226
rect 502814 298170 502882 298226
rect 502938 298170 533478 298226
rect 533534 298170 533602 298226
rect 533658 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 71102 298118 597980 298170
rect -1916 298102 597980 298118
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 39954 298102
rect 40010 298046 40078 298102
rect 40134 298046 40202 298102
rect 40258 298046 40326 298102
rect 40382 298046 101394 298102
rect 101450 298046 101518 298102
rect 101574 298046 101642 298102
rect 101698 298046 101766 298102
rect 101822 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 209878 298102
rect 209934 298046 210002 298102
rect 210058 298046 240598 298102
rect 240654 298046 240722 298102
rect 240778 298046 271318 298102
rect 271374 298046 271442 298102
rect 271498 298046 302038 298102
rect 302094 298046 302162 298102
rect 302218 298046 332758 298102
rect 332814 298046 332882 298102
rect 332938 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 379878 298102
rect 379934 298046 380002 298102
rect 380058 298046 410598 298102
rect 410654 298046 410722 298102
rect 410778 298046 441318 298102
rect 441374 298046 441442 298102
rect 441498 298046 472038 298102
rect 472094 298046 472162 298102
rect 472218 298046 502758 298102
rect 502814 298046 502882 298102
rect 502938 298046 533478 298102
rect 533534 298046 533602 298102
rect 533658 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 39954 297978
rect 40010 297922 40078 297978
rect 40134 297922 40202 297978
rect 40258 297922 40326 297978
rect 40382 297922 101394 297978
rect 101450 297922 101518 297978
rect 101574 297922 101642 297978
rect 101698 297922 101766 297978
rect 101822 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 209878 297978
rect 209934 297922 210002 297978
rect 210058 297922 240598 297978
rect 240654 297922 240722 297978
rect 240778 297922 271318 297978
rect 271374 297922 271442 297978
rect 271498 297922 302038 297978
rect 302094 297922 302162 297978
rect 302218 297922 332758 297978
rect 332814 297922 332882 297978
rect 332938 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 379878 297978
rect 379934 297922 380002 297978
rect 380058 297922 410598 297978
rect 410654 297922 410722 297978
rect 410778 297922 441318 297978
rect 441374 297922 441442 297978
rect 441498 297922 472038 297978
rect 472094 297922 472162 297978
rect 472218 297922 502758 297978
rect 502814 297922 502882 297978
rect 502938 297922 533478 297978
rect 533534 297922 533602 297978
rect 533658 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect 356508 296758 360292 296774
rect 356508 296702 356524 296758
rect 356580 296702 360220 296758
rect 360276 296702 360292 296758
rect 356508 296686 360292 296702
rect 342732 292618 362084 292634
rect 342732 292562 342748 292618
rect 342804 292562 362012 292618
rect 362068 292562 362084 292618
rect 342732 292546 362084 292562
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 44518 292350
rect 44574 292294 44642 292350
rect 44698 292294 75238 292350
rect 75294 292294 75362 292350
rect 75418 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 194518 292350
rect 194574 292294 194642 292350
rect 194698 292294 225238 292350
rect 225294 292294 225362 292350
rect 225418 292294 255958 292350
rect 256014 292294 256082 292350
rect 256138 292294 286678 292350
rect 286734 292294 286802 292350
rect 286858 292294 317398 292350
rect 317454 292294 317522 292350
rect 317578 292294 343434 292350
rect 343490 292294 343558 292350
rect 343614 292294 343682 292350
rect 343738 292294 343806 292350
rect 343862 292294 364518 292350
rect 364574 292294 364642 292350
rect 364698 292294 395238 292350
rect 395294 292294 395362 292350
rect 395418 292294 425958 292350
rect 426014 292294 426082 292350
rect 426138 292294 456678 292350
rect 456734 292294 456802 292350
rect 456858 292294 487398 292350
rect 487454 292294 487522 292350
rect 487578 292294 518118 292350
rect 518174 292294 518242 292350
rect 518298 292294 548838 292350
rect 548894 292294 548962 292350
rect 549018 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 44518 292226
rect 44574 292170 44642 292226
rect 44698 292170 75238 292226
rect 75294 292170 75362 292226
rect 75418 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 194518 292226
rect 194574 292170 194642 292226
rect 194698 292170 225238 292226
rect 225294 292170 225362 292226
rect 225418 292170 255958 292226
rect 256014 292170 256082 292226
rect 256138 292170 286678 292226
rect 286734 292170 286802 292226
rect 286858 292170 317398 292226
rect 317454 292170 317522 292226
rect 317578 292170 343434 292226
rect 343490 292170 343558 292226
rect 343614 292170 343682 292226
rect 343738 292170 343806 292226
rect 343862 292170 364518 292226
rect 364574 292170 364642 292226
rect 364698 292170 395238 292226
rect 395294 292170 395362 292226
rect 395418 292170 425958 292226
rect 426014 292170 426082 292226
rect 426138 292170 456678 292226
rect 456734 292170 456802 292226
rect 456858 292170 487398 292226
rect 487454 292170 487522 292226
rect 487578 292170 518118 292226
rect 518174 292170 518242 292226
rect 518298 292170 548838 292226
rect 548894 292170 548962 292226
rect 549018 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 44518 292102
rect 44574 292046 44642 292102
rect 44698 292046 75238 292102
rect 75294 292046 75362 292102
rect 75418 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 194518 292102
rect 194574 292046 194642 292102
rect 194698 292046 225238 292102
rect 225294 292046 225362 292102
rect 225418 292046 255958 292102
rect 256014 292046 256082 292102
rect 256138 292046 286678 292102
rect 286734 292046 286802 292102
rect 286858 292046 317398 292102
rect 317454 292046 317522 292102
rect 317578 292046 343434 292102
rect 343490 292046 343558 292102
rect 343614 292046 343682 292102
rect 343738 292046 343806 292102
rect 343862 292046 364518 292102
rect 364574 292046 364642 292102
rect 364698 292046 395238 292102
rect 395294 292046 395362 292102
rect 395418 292046 425958 292102
rect 426014 292046 426082 292102
rect 426138 292046 456678 292102
rect 456734 292046 456802 292102
rect 456858 292046 487398 292102
rect 487454 292046 487522 292102
rect 487578 292046 518118 292102
rect 518174 292046 518242 292102
rect 518298 292046 548838 292102
rect 548894 292046 548962 292102
rect 549018 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 44518 291978
rect 44574 291922 44642 291978
rect 44698 291922 75238 291978
rect 75294 291922 75362 291978
rect 75418 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 194518 291978
rect 194574 291922 194642 291978
rect 194698 291922 225238 291978
rect 225294 291922 225362 291978
rect 225418 291922 255958 291978
rect 256014 291922 256082 291978
rect 256138 291922 286678 291978
rect 286734 291922 286802 291978
rect 286858 291922 317398 291978
rect 317454 291922 317522 291978
rect 317578 291922 343434 291978
rect 343490 291922 343558 291978
rect 343614 291922 343682 291978
rect 343738 291922 343806 291978
rect 343862 291922 364518 291978
rect 364574 291922 364642 291978
rect 364698 291922 395238 291978
rect 395294 291922 395362 291978
rect 395418 291922 425958 291978
rect 426014 291922 426082 291978
rect 426138 291922 456678 291978
rect 456734 291922 456802 291978
rect 456858 291922 487398 291978
rect 487454 291922 487522 291978
rect 487578 291922 518118 291978
rect 518174 291922 518242 291978
rect 518298 291922 548838 291978
rect 548894 291922 548962 291978
rect 549018 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect 187276 289018 197668 289034
rect 187276 288962 187292 289018
rect 187348 288962 197596 289018
rect 197652 288962 197668 289018
rect 187276 288946 197668 288962
rect 342732 287398 360068 287414
rect 342732 287342 342748 287398
rect 342804 287342 359996 287398
rect 360052 287342 360068 287398
rect 342732 287326 360068 287342
rect 187164 287218 197556 287234
rect 187164 287162 187180 287218
rect 187236 287162 197484 287218
rect 197540 287162 197556 287218
rect 187164 287146 197556 287162
rect 188060 285778 197780 285794
rect 188060 285722 188076 285778
rect 188132 285722 197708 285778
rect 197764 285722 197780 285778
rect 188060 285706 197780 285722
rect 336908 284698 339460 284714
rect 336908 284642 336924 284698
rect 336980 284642 339388 284698
rect 339444 284642 339460 284698
rect 336908 284626 339460 284642
rect 170476 281458 197556 281474
rect 170476 281402 170492 281458
rect 170548 281402 187852 281458
rect 187908 281402 197484 281458
rect 197540 281402 197556 281458
rect 170476 281386 197556 281402
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 39954 280350
rect 40010 280294 40078 280350
rect 40134 280294 40202 280350
rect 40258 280294 40326 280350
rect 40382 280294 59878 280350
rect 59934 280294 60002 280350
rect 60058 280294 90598 280350
rect 90654 280294 90722 280350
rect 90778 280294 101394 280350
rect 101450 280294 101518 280350
rect 101574 280294 101642 280350
rect 101698 280294 101766 280350
rect 101822 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 147078 280350
rect 147134 280294 147202 280350
rect 147258 280294 152902 280350
rect 152958 280294 153026 280350
rect 153082 280294 158726 280350
rect 158782 280294 158850 280350
rect 158906 280294 164550 280350
rect 164606 280294 164674 280350
rect 164730 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 209878 280350
rect 209934 280294 210002 280350
rect 210058 280294 240598 280350
rect 240654 280294 240722 280350
rect 240778 280294 271318 280350
rect 271374 280294 271442 280350
rect 271498 280294 302038 280350
rect 302094 280294 302162 280350
rect 302218 280294 332758 280350
rect 332814 280294 332882 280350
rect 332938 280294 347154 280350
rect 347210 280294 347278 280350
rect 347334 280294 347402 280350
rect 347458 280294 347526 280350
rect 347582 280294 379878 280350
rect 379934 280294 380002 280350
rect 380058 280294 410598 280350
rect 410654 280294 410722 280350
rect 410778 280294 441318 280350
rect 441374 280294 441442 280350
rect 441498 280294 472038 280350
rect 472094 280294 472162 280350
rect 472218 280294 502758 280350
rect 502814 280294 502882 280350
rect 502938 280294 533478 280350
rect 533534 280294 533602 280350
rect 533658 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 39954 280226
rect 40010 280170 40078 280226
rect 40134 280170 40202 280226
rect 40258 280170 40326 280226
rect 40382 280170 59878 280226
rect 59934 280170 60002 280226
rect 60058 280170 90598 280226
rect 90654 280170 90722 280226
rect 90778 280170 101394 280226
rect 101450 280170 101518 280226
rect 101574 280170 101642 280226
rect 101698 280170 101766 280226
rect 101822 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 147078 280226
rect 147134 280170 147202 280226
rect 147258 280170 152902 280226
rect 152958 280170 153026 280226
rect 153082 280170 158726 280226
rect 158782 280170 158850 280226
rect 158906 280170 164550 280226
rect 164606 280170 164674 280226
rect 164730 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 209878 280226
rect 209934 280170 210002 280226
rect 210058 280170 240598 280226
rect 240654 280170 240722 280226
rect 240778 280170 271318 280226
rect 271374 280170 271442 280226
rect 271498 280170 302038 280226
rect 302094 280170 302162 280226
rect 302218 280170 332758 280226
rect 332814 280170 332882 280226
rect 332938 280170 347154 280226
rect 347210 280170 347278 280226
rect 347334 280170 347402 280226
rect 347458 280170 347526 280226
rect 347582 280170 379878 280226
rect 379934 280170 380002 280226
rect 380058 280170 410598 280226
rect 410654 280170 410722 280226
rect 410778 280170 441318 280226
rect 441374 280170 441442 280226
rect 441498 280170 472038 280226
rect 472094 280170 472162 280226
rect 472218 280170 502758 280226
rect 502814 280170 502882 280226
rect 502938 280170 533478 280226
rect 533534 280170 533602 280226
rect 533658 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 39954 280102
rect 40010 280046 40078 280102
rect 40134 280046 40202 280102
rect 40258 280046 40326 280102
rect 40382 280046 59878 280102
rect 59934 280046 60002 280102
rect 60058 280046 90598 280102
rect 90654 280046 90722 280102
rect 90778 280046 101394 280102
rect 101450 280046 101518 280102
rect 101574 280046 101642 280102
rect 101698 280046 101766 280102
rect 101822 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 147078 280102
rect 147134 280046 147202 280102
rect 147258 280046 152902 280102
rect 152958 280046 153026 280102
rect 153082 280046 158726 280102
rect 158782 280046 158850 280102
rect 158906 280046 164550 280102
rect 164606 280046 164674 280102
rect 164730 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 209878 280102
rect 209934 280046 210002 280102
rect 210058 280046 240598 280102
rect 240654 280046 240722 280102
rect 240778 280046 271318 280102
rect 271374 280046 271442 280102
rect 271498 280046 302038 280102
rect 302094 280046 302162 280102
rect 302218 280046 332758 280102
rect 332814 280046 332882 280102
rect 332938 280046 347154 280102
rect 347210 280046 347278 280102
rect 347334 280046 347402 280102
rect 347458 280046 347526 280102
rect 347582 280046 379878 280102
rect 379934 280046 380002 280102
rect 380058 280046 410598 280102
rect 410654 280046 410722 280102
rect 410778 280046 441318 280102
rect 441374 280046 441442 280102
rect 441498 280046 472038 280102
rect 472094 280046 472162 280102
rect 472218 280046 502758 280102
rect 502814 280046 502882 280102
rect 502938 280046 533478 280102
rect 533534 280046 533602 280102
rect 533658 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 39954 279978
rect 40010 279922 40078 279978
rect 40134 279922 40202 279978
rect 40258 279922 40326 279978
rect 40382 279922 59878 279978
rect 59934 279922 60002 279978
rect 60058 279922 90598 279978
rect 90654 279922 90722 279978
rect 90778 279922 101394 279978
rect 101450 279922 101518 279978
rect 101574 279922 101642 279978
rect 101698 279922 101766 279978
rect 101822 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 147078 279978
rect 147134 279922 147202 279978
rect 147258 279922 152902 279978
rect 152958 279922 153026 279978
rect 153082 279922 158726 279978
rect 158782 279922 158850 279978
rect 158906 279922 164550 279978
rect 164606 279922 164674 279978
rect 164730 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 209878 279978
rect 209934 279922 210002 279978
rect 210058 279922 240598 279978
rect 240654 279922 240722 279978
rect 240778 279922 271318 279978
rect 271374 279922 271442 279978
rect 271498 279922 302038 279978
rect 302094 279922 302162 279978
rect 302218 279922 332758 279978
rect 332814 279922 332882 279978
rect 332938 279922 347154 279978
rect 347210 279922 347278 279978
rect 347334 279922 347402 279978
rect 347458 279922 347526 279978
rect 347582 279922 379878 279978
rect 379934 279922 380002 279978
rect 380058 279922 410598 279978
rect 410654 279922 410722 279978
rect 410778 279922 441318 279978
rect 441374 279922 441442 279978
rect 441498 279922 472038 279978
rect 472094 279922 472162 279978
rect 472218 279922 502758 279978
rect 502814 279922 502882 279978
rect 502938 279922 533478 279978
rect 533534 279922 533602 279978
rect 533658 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect 337244 279658 339460 279674
rect 337244 279602 337260 279658
rect 337316 279602 339388 279658
rect 339444 279602 339460 279658
rect 337244 279586 339460 279602
rect 337020 277318 339348 277334
rect 337020 277262 337036 277318
rect 337092 277262 339276 277318
rect 339332 277262 339348 277318
rect 337020 277246 339348 277262
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 44518 274350
rect 44574 274294 44642 274350
rect 44698 274294 75238 274350
rect 75294 274294 75362 274350
rect 75418 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 144166 274350
rect 144222 274294 144290 274350
rect 144346 274294 149990 274350
rect 150046 274294 150114 274350
rect 150170 274294 155814 274350
rect 155870 274294 155938 274350
rect 155994 274294 161638 274350
rect 161694 274294 161762 274350
rect 161818 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 194518 274350
rect 194574 274294 194642 274350
rect 194698 274294 225238 274350
rect 225294 274294 225362 274350
rect 225418 274294 255958 274350
rect 256014 274294 256082 274350
rect 256138 274294 286678 274350
rect 286734 274294 286802 274350
rect 286858 274294 317398 274350
rect 317454 274294 317522 274350
rect 317578 274294 343434 274350
rect 343490 274294 343558 274350
rect 343614 274294 343682 274350
rect 343738 274294 343806 274350
rect 343862 274294 364518 274350
rect 364574 274294 364642 274350
rect 364698 274294 395238 274350
rect 395294 274294 395362 274350
rect 395418 274294 425958 274350
rect 426014 274294 426082 274350
rect 426138 274294 456678 274350
rect 456734 274294 456802 274350
rect 456858 274294 487398 274350
rect 487454 274294 487522 274350
rect 487578 274294 518118 274350
rect 518174 274294 518242 274350
rect 518298 274294 548838 274350
rect 548894 274294 548962 274350
rect 549018 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 44518 274226
rect 44574 274170 44642 274226
rect 44698 274170 75238 274226
rect 75294 274170 75362 274226
rect 75418 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 144166 274226
rect 144222 274170 144290 274226
rect 144346 274170 149990 274226
rect 150046 274170 150114 274226
rect 150170 274170 155814 274226
rect 155870 274170 155938 274226
rect 155994 274170 161638 274226
rect 161694 274170 161762 274226
rect 161818 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 194518 274226
rect 194574 274170 194642 274226
rect 194698 274170 225238 274226
rect 225294 274170 225362 274226
rect 225418 274170 255958 274226
rect 256014 274170 256082 274226
rect 256138 274170 286678 274226
rect 286734 274170 286802 274226
rect 286858 274170 317398 274226
rect 317454 274170 317522 274226
rect 317578 274170 343434 274226
rect 343490 274170 343558 274226
rect 343614 274170 343682 274226
rect 343738 274170 343806 274226
rect 343862 274170 364518 274226
rect 364574 274170 364642 274226
rect 364698 274170 395238 274226
rect 395294 274170 395362 274226
rect 395418 274170 425958 274226
rect 426014 274170 426082 274226
rect 426138 274170 456678 274226
rect 456734 274170 456802 274226
rect 456858 274170 487398 274226
rect 487454 274170 487522 274226
rect 487578 274170 518118 274226
rect 518174 274170 518242 274226
rect 518298 274170 548838 274226
rect 548894 274170 548962 274226
rect 549018 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 44518 274102
rect 44574 274046 44642 274102
rect 44698 274046 75238 274102
rect 75294 274046 75362 274102
rect 75418 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 144166 274102
rect 144222 274046 144290 274102
rect 144346 274046 149990 274102
rect 150046 274046 150114 274102
rect 150170 274046 155814 274102
rect 155870 274046 155938 274102
rect 155994 274046 161638 274102
rect 161694 274046 161762 274102
rect 161818 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 194518 274102
rect 194574 274046 194642 274102
rect 194698 274046 225238 274102
rect 225294 274046 225362 274102
rect 225418 274046 255958 274102
rect 256014 274046 256082 274102
rect 256138 274046 286678 274102
rect 286734 274046 286802 274102
rect 286858 274046 317398 274102
rect 317454 274046 317522 274102
rect 317578 274046 343434 274102
rect 343490 274046 343558 274102
rect 343614 274046 343682 274102
rect 343738 274046 343806 274102
rect 343862 274046 364518 274102
rect 364574 274046 364642 274102
rect 364698 274046 395238 274102
rect 395294 274046 395362 274102
rect 395418 274046 425958 274102
rect 426014 274046 426082 274102
rect 426138 274046 456678 274102
rect 456734 274046 456802 274102
rect 456858 274046 487398 274102
rect 487454 274046 487522 274102
rect 487578 274046 518118 274102
rect 518174 274046 518242 274102
rect 518298 274046 548838 274102
rect 548894 274046 548962 274102
rect 549018 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 44518 273978
rect 44574 273922 44642 273978
rect 44698 273922 75238 273978
rect 75294 273922 75362 273978
rect 75418 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 144166 273978
rect 144222 273922 144290 273978
rect 144346 273922 149990 273978
rect 150046 273922 150114 273978
rect 150170 273922 155814 273978
rect 155870 273922 155938 273978
rect 155994 273922 161638 273978
rect 161694 273922 161762 273978
rect 161818 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 194518 273978
rect 194574 273922 194642 273978
rect 194698 273922 225238 273978
rect 225294 273922 225362 273978
rect 225418 273922 255958 273978
rect 256014 273922 256082 273978
rect 256138 273922 286678 273978
rect 286734 273922 286802 273978
rect 286858 273922 317398 273978
rect 317454 273922 317522 273978
rect 317578 273922 343434 273978
rect 343490 273922 343558 273978
rect 343614 273922 343682 273978
rect 343738 273922 343806 273978
rect 343862 273922 364518 273978
rect 364574 273922 364642 273978
rect 364698 273922 395238 273978
rect 395294 273922 395362 273978
rect 395418 273922 425958 273978
rect 426014 273922 426082 273978
rect 426138 273922 456678 273978
rect 456734 273922 456802 273978
rect 456858 273922 487398 273978
rect 487454 273922 487522 273978
rect 487578 273922 518118 273978
rect 518174 273922 518242 273978
rect 518298 273922 548838 273978
rect 548894 273922 548962 273978
rect 549018 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect 186380 268858 198116 268874
rect 186380 268802 186396 268858
rect 186452 268802 198044 268858
rect 198100 268802 198116 268858
rect 186380 268786 198116 268802
rect 337636 267418 339348 267434
rect 337636 267362 339276 267418
rect 339332 267362 339348 267418
rect 337636 267346 339348 267362
rect 337636 267254 337724 267346
rect 337132 267238 337724 267254
rect 337132 267182 337148 267238
rect 337204 267182 337724 267238
rect 337132 267166 337724 267182
rect 338700 264358 339460 264374
rect 338700 264302 338716 264358
rect 338772 264302 339388 264358
rect 339444 264302 339460 264358
rect 338700 264286 339460 264302
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 39954 262350
rect 40010 262294 40078 262350
rect 40134 262294 40202 262350
rect 40258 262294 40326 262350
rect 40382 262294 59878 262350
rect 59934 262294 60002 262350
rect 60058 262294 90598 262350
rect 90654 262294 90722 262350
rect 90778 262294 101394 262350
rect 101450 262294 101518 262350
rect 101574 262294 101642 262350
rect 101698 262294 101766 262350
rect 101822 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 209878 262350
rect 209934 262294 210002 262350
rect 210058 262294 240598 262350
rect 240654 262294 240722 262350
rect 240778 262294 271318 262350
rect 271374 262294 271442 262350
rect 271498 262294 302038 262350
rect 302094 262294 302162 262350
rect 302218 262294 332758 262350
rect 332814 262294 332882 262350
rect 332938 262294 347154 262350
rect 347210 262294 347278 262350
rect 347334 262294 347402 262350
rect 347458 262294 347526 262350
rect 347582 262294 379878 262350
rect 379934 262294 380002 262350
rect 380058 262294 410598 262350
rect 410654 262294 410722 262350
rect 410778 262294 441318 262350
rect 441374 262294 441442 262350
rect 441498 262294 472038 262350
rect 472094 262294 472162 262350
rect 472218 262294 502758 262350
rect 502814 262294 502882 262350
rect 502938 262294 533478 262350
rect 533534 262294 533602 262350
rect 533658 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 39954 262226
rect 40010 262170 40078 262226
rect 40134 262170 40202 262226
rect 40258 262170 40326 262226
rect 40382 262170 59878 262226
rect 59934 262170 60002 262226
rect 60058 262170 90598 262226
rect 90654 262170 90722 262226
rect 90778 262170 101394 262226
rect 101450 262170 101518 262226
rect 101574 262170 101642 262226
rect 101698 262170 101766 262226
rect 101822 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 209878 262226
rect 209934 262170 210002 262226
rect 210058 262170 240598 262226
rect 240654 262170 240722 262226
rect 240778 262170 271318 262226
rect 271374 262170 271442 262226
rect 271498 262170 302038 262226
rect 302094 262170 302162 262226
rect 302218 262170 332758 262226
rect 332814 262170 332882 262226
rect 332938 262170 347154 262226
rect 347210 262170 347278 262226
rect 347334 262170 347402 262226
rect 347458 262170 347526 262226
rect 347582 262170 379878 262226
rect 379934 262170 380002 262226
rect 380058 262170 410598 262226
rect 410654 262170 410722 262226
rect 410778 262170 441318 262226
rect 441374 262170 441442 262226
rect 441498 262170 472038 262226
rect 472094 262170 472162 262226
rect 472218 262170 502758 262226
rect 502814 262170 502882 262226
rect 502938 262170 533478 262226
rect 533534 262170 533602 262226
rect 533658 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 39954 262102
rect 40010 262046 40078 262102
rect 40134 262046 40202 262102
rect 40258 262046 40326 262102
rect 40382 262046 59878 262102
rect 59934 262046 60002 262102
rect 60058 262046 90598 262102
rect 90654 262046 90722 262102
rect 90778 262046 101394 262102
rect 101450 262046 101518 262102
rect 101574 262046 101642 262102
rect 101698 262046 101766 262102
rect 101822 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 209878 262102
rect 209934 262046 210002 262102
rect 210058 262046 240598 262102
rect 240654 262046 240722 262102
rect 240778 262046 271318 262102
rect 271374 262046 271442 262102
rect 271498 262046 302038 262102
rect 302094 262046 302162 262102
rect 302218 262046 332758 262102
rect 332814 262046 332882 262102
rect 332938 262046 347154 262102
rect 347210 262046 347278 262102
rect 347334 262046 347402 262102
rect 347458 262046 347526 262102
rect 347582 262046 379878 262102
rect 379934 262046 380002 262102
rect 380058 262046 410598 262102
rect 410654 262046 410722 262102
rect 410778 262046 441318 262102
rect 441374 262046 441442 262102
rect 441498 262046 472038 262102
rect 472094 262046 472162 262102
rect 472218 262046 502758 262102
rect 502814 262046 502882 262102
rect 502938 262046 533478 262102
rect 533534 262046 533602 262102
rect 533658 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 39954 261978
rect 40010 261922 40078 261978
rect 40134 261922 40202 261978
rect 40258 261922 40326 261978
rect 40382 261922 59878 261978
rect 59934 261922 60002 261978
rect 60058 261922 90598 261978
rect 90654 261922 90722 261978
rect 90778 261922 101394 261978
rect 101450 261922 101518 261978
rect 101574 261922 101642 261978
rect 101698 261922 101766 261978
rect 101822 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 209878 261978
rect 209934 261922 210002 261978
rect 210058 261922 240598 261978
rect 240654 261922 240722 261978
rect 240778 261922 271318 261978
rect 271374 261922 271442 261978
rect 271498 261922 302038 261978
rect 302094 261922 302162 261978
rect 302218 261922 332758 261978
rect 332814 261922 332882 261978
rect 332938 261922 347154 261978
rect 347210 261922 347278 261978
rect 347334 261922 347402 261978
rect 347458 261922 347526 261978
rect 347582 261922 379878 261978
rect 379934 261922 380002 261978
rect 380058 261922 410598 261978
rect 410654 261922 410722 261978
rect 410778 261922 441318 261978
rect 441374 261922 441442 261978
rect 441498 261922 472038 261978
rect 472094 261922 472162 261978
rect 472218 261922 502758 261978
rect 502814 261922 502882 261978
rect 502938 261922 533478 261978
rect 533534 261922 533602 261978
rect 533658 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect 338588 258778 339572 258794
rect 338588 258722 338604 258778
rect 338660 258722 339500 258778
rect 339556 258722 339572 258778
rect 338588 258706 339572 258722
rect 337356 257878 339572 257894
rect 337356 257822 337372 257878
rect 337428 257822 339500 257878
rect 339556 257822 339572 257878
rect 337356 257806 339572 257822
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 44518 256350
rect 44574 256294 44642 256350
rect 44698 256294 75238 256350
rect 75294 256294 75362 256350
rect 75418 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 194518 256350
rect 194574 256294 194642 256350
rect 194698 256294 225238 256350
rect 225294 256294 225362 256350
rect 225418 256294 255958 256350
rect 256014 256294 256082 256350
rect 256138 256294 286678 256350
rect 286734 256294 286802 256350
rect 286858 256294 317398 256350
rect 317454 256294 317522 256350
rect 317578 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 364518 256350
rect 364574 256294 364642 256350
rect 364698 256294 395238 256350
rect 395294 256294 395362 256350
rect 395418 256294 425958 256350
rect 426014 256294 426082 256350
rect 426138 256294 456678 256350
rect 456734 256294 456802 256350
rect 456858 256294 487398 256350
rect 487454 256294 487522 256350
rect 487578 256294 518118 256350
rect 518174 256294 518242 256350
rect 518298 256294 548838 256350
rect 548894 256294 548962 256350
rect 549018 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 44518 256226
rect 44574 256170 44642 256226
rect 44698 256170 75238 256226
rect 75294 256170 75362 256226
rect 75418 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 194518 256226
rect 194574 256170 194642 256226
rect 194698 256170 225238 256226
rect 225294 256170 225362 256226
rect 225418 256170 255958 256226
rect 256014 256170 256082 256226
rect 256138 256170 286678 256226
rect 286734 256170 286802 256226
rect 286858 256170 317398 256226
rect 317454 256170 317522 256226
rect 317578 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 364518 256226
rect 364574 256170 364642 256226
rect 364698 256170 395238 256226
rect 395294 256170 395362 256226
rect 395418 256170 425958 256226
rect 426014 256170 426082 256226
rect 426138 256170 456678 256226
rect 456734 256170 456802 256226
rect 456858 256170 487398 256226
rect 487454 256170 487522 256226
rect 487578 256170 518118 256226
rect 518174 256170 518242 256226
rect 518298 256170 548838 256226
rect 548894 256170 548962 256226
rect 549018 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 44518 256102
rect 44574 256046 44642 256102
rect 44698 256046 75238 256102
rect 75294 256046 75362 256102
rect 75418 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 194518 256102
rect 194574 256046 194642 256102
rect 194698 256046 225238 256102
rect 225294 256046 225362 256102
rect 225418 256046 255958 256102
rect 256014 256046 256082 256102
rect 256138 256046 286678 256102
rect 286734 256046 286802 256102
rect 286858 256046 317398 256102
rect 317454 256046 317522 256102
rect 317578 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 364518 256102
rect 364574 256046 364642 256102
rect 364698 256046 395238 256102
rect 395294 256046 395362 256102
rect 395418 256046 425958 256102
rect 426014 256046 426082 256102
rect 426138 256046 456678 256102
rect 456734 256046 456802 256102
rect 456858 256046 487398 256102
rect 487454 256046 487522 256102
rect 487578 256046 518118 256102
rect 518174 256046 518242 256102
rect 518298 256046 548838 256102
rect 548894 256046 548962 256102
rect 549018 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 44518 255978
rect 44574 255922 44642 255978
rect 44698 255922 75238 255978
rect 75294 255922 75362 255978
rect 75418 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 194518 255978
rect 194574 255922 194642 255978
rect 194698 255922 225238 255978
rect 225294 255922 225362 255978
rect 225418 255922 255958 255978
rect 256014 255922 256082 255978
rect 256138 255922 286678 255978
rect 286734 255922 286802 255978
rect 286858 255922 317398 255978
rect 317454 255922 317522 255978
rect 317578 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 364518 255978
rect 364574 255922 364642 255978
rect 364698 255922 395238 255978
rect 395294 255922 395362 255978
rect 395418 255922 425958 255978
rect 426014 255922 426082 255978
rect 426138 255922 456678 255978
rect 456734 255922 456802 255978
rect 456858 255922 487398 255978
rect 487454 255922 487522 255978
rect 487578 255922 518118 255978
rect 518174 255922 518242 255978
rect 518298 255922 548838 255978
rect 548894 255922 548962 255978
rect 549018 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect 338812 255718 339348 255734
rect 338812 255662 338828 255718
rect 338884 255662 339276 255718
rect 339332 255662 339348 255718
rect 338812 255646 339348 255662
rect 359308 255718 360516 255734
rect 359308 255662 359324 255718
rect 359380 255662 360444 255718
rect 360500 255662 360516 255718
rect 359308 255646 360516 255662
rect 337468 254818 339348 254834
rect 337468 254762 337484 254818
rect 337540 254762 339276 254818
rect 339332 254762 339348 254818
rect 337468 254746 339348 254762
rect 338364 254638 339348 254654
rect 338364 254582 338380 254638
rect 338436 254582 339276 254638
rect 339332 254582 339348 254638
rect 338364 254566 339348 254582
rect 335788 253558 337332 253574
rect 335788 253502 335804 253558
rect 335860 253502 337260 253558
rect 337316 253502 337332 253558
rect 335788 253486 337332 253502
rect 336796 253018 345172 253034
rect 336796 252962 336812 253018
rect 336868 252962 345100 253018
rect 345156 252962 345172 253018
rect 336796 252946 345172 252962
rect 190636 249778 197892 249794
rect 190636 249722 190652 249778
rect 190708 249722 197820 249778
rect 197876 249722 197892 249778
rect 190636 249706 197892 249722
rect 338924 248878 339348 248894
rect 338924 248822 338940 248878
rect 338996 248822 339276 248878
rect 339332 248822 339348 248878
rect 338924 248806 339348 248822
rect 190636 248698 194308 248714
rect 190636 248642 190652 248698
rect 190708 248642 194236 248698
rect 194292 248642 194308 248698
rect 190636 248626 194308 248642
rect 338252 248698 339124 248714
rect 338252 248642 338268 248698
rect 338324 248642 339052 248698
rect 339108 248642 339124 248698
rect 338252 248626 339124 248642
rect 190636 247258 198004 247274
rect 190636 247202 190652 247258
rect 190708 247202 197932 247258
rect 197988 247202 198004 247258
rect 190636 247186 198004 247202
rect 4156 247078 46244 247094
rect 4156 247022 4172 247078
rect 4228 247022 46172 247078
rect 46228 247022 46244 247078
rect 4156 247006 46244 247022
rect 337580 246358 339460 246374
rect 337580 246302 337596 246358
rect 337652 246302 339388 246358
rect 339444 246302 339460 246358
rect 337580 246286 339460 246302
rect 337244 244738 341252 244754
rect 337244 244682 337260 244738
rect 337316 244682 341180 244738
rect 341236 244682 341252 244738
rect 337244 244666 341252 244682
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 39954 244350
rect 40010 244294 40078 244350
rect 40134 244294 40202 244350
rect 40258 244294 40326 244350
rect 40382 244294 59878 244350
rect 59934 244294 60002 244350
rect 60058 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 90598 244350
rect 90654 244294 90722 244350
rect 90778 244294 101394 244350
rect 101450 244294 101518 244350
rect 101574 244294 101642 244350
rect 101698 244294 101766 244350
rect 101822 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 209878 244350
rect 209934 244294 210002 244350
rect 210058 244294 240598 244350
rect 240654 244294 240722 244350
rect 240778 244294 271318 244350
rect 271374 244294 271442 244350
rect 271498 244294 302038 244350
rect 302094 244294 302162 244350
rect 302218 244294 332758 244350
rect 332814 244294 332882 244350
rect 332938 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 379878 244350
rect 379934 244294 380002 244350
rect 380058 244294 410598 244350
rect 410654 244294 410722 244350
rect 410778 244294 441318 244350
rect 441374 244294 441442 244350
rect 441498 244294 472038 244350
rect 472094 244294 472162 244350
rect 472218 244294 502758 244350
rect 502814 244294 502882 244350
rect 502938 244294 533478 244350
rect 533534 244294 533602 244350
rect 533658 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 39954 244226
rect 40010 244170 40078 244226
rect 40134 244170 40202 244226
rect 40258 244170 40326 244226
rect 40382 244170 59878 244226
rect 59934 244170 60002 244226
rect 60058 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 90598 244226
rect 90654 244170 90722 244226
rect 90778 244170 101394 244226
rect 101450 244170 101518 244226
rect 101574 244170 101642 244226
rect 101698 244170 101766 244226
rect 101822 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 209878 244226
rect 209934 244170 210002 244226
rect 210058 244170 240598 244226
rect 240654 244170 240722 244226
rect 240778 244170 271318 244226
rect 271374 244170 271442 244226
rect 271498 244170 302038 244226
rect 302094 244170 302162 244226
rect 302218 244170 332758 244226
rect 332814 244170 332882 244226
rect 332938 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 379878 244226
rect 379934 244170 380002 244226
rect 380058 244170 410598 244226
rect 410654 244170 410722 244226
rect 410778 244170 441318 244226
rect 441374 244170 441442 244226
rect 441498 244170 472038 244226
rect 472094 244170 472162 244226
rect 472218 244170 502758 244226
rect 502814 244170 502882 244226
rect 502938 244170 533478 244226
rect 533534 244170 533602 244226
rect 533658 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 39954 244102
rect 40010 244046 40078 244102
rect 40134 244046 40202 244102
rect 40258 244046 40326 244102
rect 40382 244046 59878 244102
rect 59934 244046 60002 244102
rect 60058 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 90598 244102
rect 90654 244046 90722 244102
rect 90778 244046 101394 244102
rect 101450 244046 101518 244102
rect 101574 244046 101642 244102
rect 101698 244046 101766 244102
rect 101822 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 209878 244102
rect 209934 244046 210002 244102
rect 210058 244046 240598 244102
rect 240654 244046 240722 244102
rect 240778 244046 271318 244102
rect 271374 244046 271442 244102
rect 271498 244046 302038 244102
rect 302094 244046 302162 244102
rect 302218 244046 332758 244102
rect 332814 244046 332882 244102
rect 332938 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 379878 244102
rect 379934 244046 380002 244102
rect 380058 244046 410598 244102
rect 410654 244046 410722 244102
rect 410778 244046 441318 244102
rect 441374 244046 441442 244102
rect 441498 244046 472038 244102
rect 472094 244046 472162 244102
rect 472218 244046 502758 244102
rect 502814 244046 502882 244102
rect 502938 244046 533478 244102
rect 533534 244046 533602 244102
rect 533658 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 39954 243978
rect 40010 243922 40078 243978
rect 40134 243922 40202 243978
rect 40258 243922 40326 243978
rect 40382 243922 59878 243978
rect 59934 243922 60002 243978
rect 60058 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 90598 243978
rect 90654 243922 90722 243978
rect 90778 243922 101394 243978
rect 101450 243922 101518 243978
rect 101574 243922 101642 243978
rect 101698 243922 101766 243978
rect 101822 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 209878 243978
rect 209934 243922 210002 243978
rect 210058 243922 240598 243978
rect 240654 243922 240722 243978
rect 240778 243922 271318 243978
rect 271374 243922 271442 243978
rect 271498 243922 302038 243978
rect 302094 243922 302162 243978
rect 302218 243922 332758 243978
rect 332814 243922 332882 243978
rect 332938 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 379878 243978
rect 379934 243922 380002 243978
rect 380058 243922 410598 243978
rect 410654 243922 410722 243978
rect 410778 243922 441318 243978
rect 441374 243922 441442 243978
rect 441498 243922 472038 243978
rect 472094 243922 472162 243978
rect 472218 243922 502758 243978
rect 502814 243922 502882 243978
rect 502938 243922 533478 243978
rect 533534 243922 533602 243978
rect 533658 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect 190860 243118 346292 243134
rect 190860 243062 190876 243118
rect 190932 243062 346220 243118
rect 346276 243062 346292 243118
rect 190860 243046 346292 243062
rect 323244 242758 355924 242774
rect 323244 242702 323260 242758
rect 323316 242702 355852 242758
rect 355908 242702 355924 242758
rect 323244 242686 355924 242702
rect 190636 242038 278084 242054
rect 190636 241982 190652 242038
rect 190708 241982 278012 242038
rect 278068 241982 278084 242038
rect 190636 241966 278084 241982
rect 334220 242038 348532 242054
rect 334220 241982 334236 242038
rect 334292 241982 348460 242038
rect 348516 241982 348532 242038
rect 334220 241966 348532 241982
rect 336796 241858 339572 241874
rect 336796 241802 336812 241858
rect 336868 241802 339500 241858
rect 339556 241802 339572 241858
rect 336796 241786 339572 241802
rect 336572 241678 340468 241694
rect 336572 241622 336588 241678
rect 336644 241622 340396 241678
rect 340452 241622 340468 241678
rect 336572 241606 340468 241622
rect 35180 241138 343156 241154
rect 35180 241082 35196 241138
rect 35252 241082 343084 241138
rect 343140 241082 343156 241138
rect 35180 241066 343156 241082
rect 284940 240778 335988 240794
rect 284940 240722 284956 240778
rect 285012 240722 335916 240778
rect 335972 240722 335988 240778
rect 284940 240706 335988 240722
rect 281356 240598 334196 240614
rect 281356 240542 281372 240598
rect 281428 240542 334124 240598
rect 334180 240542 334196 240598
rect 281356 240526 334196 240542
rect 284716 240418 337780 240434
rect 284716 240362 284732 240418
rect 284788 240362 337708 240418
rect 337764 240362 337780 240418
rect 284716 240346 337780 240362
rect 320556 240238 353572 240254
rect 320556 240182 320572 240238
rect 320628 240182 353500 240238
rect 353556 240182 353572 240238
rect 320556 240166 353572 240182
rect 319884 240058 349092 240074
rect 319884 240002 319900 240058
rect 319956 240002 349020 240058
rect 349076 240002 349092 240058
rect 319884 239986 349092 240002
rect 279676 239338 338452 239354
rect 279676 239282 279692 239338
rect 279748 239282 338380 239338
rect 338436 239282 338452 239338
rect 279676 239266 338452 239282
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 364518 238350
rect 364574 238294 364642 238350
rect 364698 238294 395238 238350
rect 395294 238294 395362 238350
rect 395418 238294 425958 238350
rect 426014 238294 426082 238350
rect 426138 238294 456678 238350
rect 456734 238294 456802 238350
rect 456858 238294 487398 238350
rect 487454 238294 487522 238350
rect 487578 238294 518118 238350
rect 518174 238294 518242 238350
rect 518298 238294 548838 238350
rect 548894 238294 548962 238350
rect 549018 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 364518 238226
rect 364574 238170 364642 238226
rect 364698 238170 395238 238226
rect 395294 238170 395362 238226
rect 395418 238170 425958 238226
rect 426014 238170 426082 238226
rect 426138 238170 456678 238226
rect 456734 238170 456802 238226
rect 456858 238170 487398 238226
rect 487454 238170 487522 238226
rect 487578 238170 518118 238226
rect 518174 238170 518242 238226
rect 518298 238170 548838 238226
rect 548894 238170 548962 238226
rect 549018 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 364518 238102
rect 364574 238046 364642 238102
rect 364698 238046 395238 238102
rect 395294 238046 395362 238102
rect 395418 238046 425958 238102
rect 426014 238046 426082 238102
rect 426138 238046 456678 238102
rect 456734 238046 456802 238102
rect 456858 238046 487398 238102
rect 487454 238046 487522 238102
rect 487578 238046 518118 238102
rect 518174 238046 518242 238102
rect 518298 238046 548838 238102
rect 548894 238046 548962 238102
rect 549018 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 364518 237978
rect 364574 237922 364642 237978
rect 364698 237922 395238 237978
rect 395294 237922 395362 237978
rect 395418 237922 425958 237978
rect 426014 237922 426082 237978
rect 426138 237922 456678 237978
rect 456734 237922 456802 237978
rect 456858 237922 487398 237978
rect 487454 237922 487522 237978
rect 487578 237922 518118 237978
rect 518174 237922 518242 237978
rect 518298 237922 548838 237978
rect 548894 237922 548962 237978
rect 549018 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect 76956 237718 110084 237734
rect 76956 237662 76972 237718
rect 77028 237662 110012 237718
rect 110068 237662 110084 237718
rect 76956 237646 110084 237662
rect 321228 237718 354468 237734
rect 321228 237662 321244 237718
rect 321300 237662 354396 237718
rect 354452 237662 354468 237718
rect 321228 237646 354468 237662
rect 72924 237538 100004 237554
rect 72924 237482 72940 237538
rect 72996 237482 99932 237538
rect 99988 237482 100004 237538
rect 72924 237466 100004 237482
rect 321900 237538 348980 237554
rect 321900 237482 321916 237538
rect 321972 237482 348908 237538
rect 348964 237482 348980 237538
rect 321900 237466 348980 237482
rect 242604 237178 275620 237194
rect 242604 237122 242620 237178
rect 242676 237122 275548 237178
rect 275604 237122 275620 237178
rect 242604 237106 275620 237122
rect 241932 236998 275732 237014
rect 241932 236942 241948 236998
rect 242004 236942 275660 236998
rect 275716 236942 275732 236998
rect 241932 236926 275732 236942
rect 285164 236098 342932 236114
rect 285164 236042 285180 236098
rect 285236 236042 342860 236098
rect 342916 236042 342932 236098
rect 285164 236026 342932 236042
rect 359644 235918 361860 235934
rect 359644 235862 359660 235918
rect 359716 235862 359996 235918
rect 360052 235862 361788 235918
rect 361844 235862 361860 235918
rect 359644 235846 361860 235862
rect 196516 235198 355924 235214
rect 196516 235142 354508 235198
rect 354564 235142 355852 235198
rect 355908 235142 355924 235198
rect 196516 235126 355924 235142
rect 196516 235034 196604 235126
rect 190636 235018 196604 235034
rect 190636 234962 190652 235018
rect 190708 234962 196604 235018
rect 190636 234946 196604 234962
rect 314956 234658 337556 234674
rect 314956 234602 314972 234658
rect 315028 234602 337484 234658
rect 337540 234602 337556 234658
rect 314956 234586 337556 234602
rect 41340 234478 233284 234494
rect 41340 234422 41356 234478
rect 41412 234422 233212 234478
rect 233268 234422 233284 234478
rect 41340 234406 233284 234422
rect 235884 234478 270580 234494
rect 235884 234422 235900 234478
rect 235956 234422 270508 234478
rect 270564 234422 270580 234478
rect 235884 234406 270580 234422
rect 283036 234478 343044 234494
rect 283036 234422 283052 234478
rect 283108 234422 342972 234478
rect 343028 234422 343044 234478
rect 283036 234406 343044 234422
rect 16700 234298 341812 234314
rect 16700 234242 16716 234298
rect 16772 234242 341740 234298
rect 341796 234242 341812 234298
rect 16700 234226 341812 234242
rect 219980 231418 269796 231434
rect 219980 231362 219996 231418
rect 220052 231362 269724 231418
rect 269780 231362 269796 231418
rect 219980 231346 269796 231362
rect 218300 231238 270916 231254
rect 218300 231182 218316 231238
rect 218372 231182 270844 231238
rect 270900 231182 270916 231238
rect 218300 231166 270916 231182
rect 25100 231058 228580 231074
rect 25100 231002 25116 231058
rect 25172 231002 228508 231058
rect 228564 231002 228580 231058
rect 25100 230986 228580 231002
rect 311596 231058 342708 231074
rect 311596 231002 311612 231058
rect 311668 231002 342636 231058
rect 342692 231002 342708 231058
rect 311596 230986 342708 231002
rect 311820 230698 320084 230714
rect 311820 230642 311836 230698
rect 311892 230642 320012 230698
rect 320068 230642 320084 230698
rect 311820 230626 320084 230642
rect 312044 230518 337724 230534
rect 312044 230462 312060 230518
rect 312116 230462 337724 230518
rect 312044 230446 337724 230462
rect 337636 230354 337724 230446
rect 35068 230338 329268 230354
rect 35068 230282 35084 230338
rect 35140 230282 329196 230338
rect 329252 230282 329268 230338
rect 35068 230266 329268 230282
rect 337636 230338 359172 230354
rect 337636 230282 357868 230338
rect 357924 230282 359100 230338
rect 359156 230282 359172 230338
rect 337636 230266 359172 230282
rect 236780 227818 269908 227834
rect 236780 227762 236796 227818
rect 236852 227762 269836 227818
rect 269892 227762 269908 227818
rect 236780 227746 269908 227762
rect 18380 227638 339796 227654
rect 18380 227582 18396 227638
rect 18452 227582 339724 227638
rect 339780 227582 339796 227638
rect 18380 227566 339796 227582
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 39954 226350
rect 40010 226294 40078 226350
rect 40134 226294 40202 226350
rect 40258 226294 40326 226350
rect 40382 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 101394 226350
rect 101450 226294 101518 226350
rect 101574 226294 101642 226350
rect 101698 226294 101766 226350
rect 101822 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 379878 226350
rect 379934 226294 380002 226350
rect 380058 226294 410598 226350
rect 410654 226294 410722 226350
rect 410778 226294 441318 226350
rect 441374 226294 441442 226350
rect 441498 226294 472038 226350
rect 472094 226294 472162 226350
rect 472218 226294 502758 226350
rect 502814 226294 502882 226350
rect 502938 226294 533478 226350
rect 533534 226294 533602 226350
rect 533658 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 39954 226226
rect 40010 226170 40078 226226
rect 40134 226170 40202 226226
rect 40258 226170 40326 226226
rect 40382 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 101394 226226
rect 101450 226170 101518 226226
rect 101574 226170 101642 226226
rect 101698 226170 101766 226226
rect 101822 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 379878 226226
rect 379934 226170 380002 226226
rect 380058 226170 410598 226226
rect 410654 226170 410722 226226
rect 410778 226170 441318 226226
rect 441374 226170 441442 226226
rect 441498 226170 472038 226226
rect 472094 226170 472162 226226
rect 472218 226170 502758 226226
rect 502814 226170 502882 226226
rect 502938 226170 533478 226226
rect 533534 226170 533602 226226
rect 533658 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 39954 226102
rect 40010 226046 40078 226102
rect 40134 226046 40202 226102
rect 40258 226046 40326 226102
rect 40382 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 101394 226102
rect 101450 226046 101518 226102
rect 101574 226046 101642 226102
rect 101698 226046 101766 226102
rect 101822 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 379878 226102
rect 379934 226046 380002 226102
rect 380058 226046 410598 226102
rect 410654 226046 410722 226102
rect 410778 226046 441318 226102
rect 441374 226046 441442 226102
rect 441498 226046 472038 226102
rect 472094 226046 472162 226102
rect 472218 226046 502758 226102
rect 502814 226046 502882 226102
rect 502938 226046 533478 226102
rect 533534 226046 533602 226102
rect 533658 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 39954 225978
rect 40010 225922 40078 225978
rect 40134 225922 40202 225978
rect 40258 225922 40326 225978
rect 40382 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 101394 225978
rect 101450 225922 101518 225978
rect 101574 225922 101642 225978
rect 101698 225922 101766 225978
rect 101822 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 379878 225978
rect 379934 225922 380002 225978
rect 380058 225922 410598 225978
rect 410654 225922 410722 225978
rect 410778 225922 441318 225978
rect 441374 225922 441442 225978
rect 441498 225922 472038 225978
rect 472094 225922 472162 225978
rect 472218 225922 502758 225978
rect 502814 225922 502882 225978
rect 502938 225922 533478 225978
rect 533534 225922 533602 225978
rect 533658 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect 20060 224218 341588 224234
rect 20060 224162 20076 224218
rect 20132 224162 341516 224218
rect 341572 224162 341588 224218
rect 20060 224146 341588 224162
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 364518 220350
rect 364574 220294 364642 220350
rect 364698 220294 395238 220350
rect 395294 220294 395362 220350
rect 395418 220294 425958 220350
rect 426014 220294 426082 220350
rect 426138 220294 456678 220350
rect 456734 220294 456802 220350
rect 456858 220294 487398 220350
rect 487454 220294 487522 220350
rect 487578 220294 518118 220350
rect 518174 220294 518242 220350
rect 518298 220294 548838 220350
rect 548894 220294 548962 220350
rect 549018 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 364518 220226
rect 364574 220170 364642 220226
rect 364698 220170 395238 220226
rect 395294 220170 395362 220226
rect 395418 220170 425958 220226
rect 426014 220170 426082 220226
rect 426138 220170 456678 220226
rect 456734 220170 456802 220226
rect 456858 220170 487398 220226
rect 487454 220170 487522 220226
rect 487578 220170 518118 220226
rect 518174 220170 518242 220226
rect 518298 220170 548838 220226
rect 548894 220170 548962 220226
rect 549018 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 364518 220102
rect 364574 220046 364642 220102
rect 364698 220046 395238 220102
rect 395294 220046 395362 220102
rect 395418 220046 425958 220102
rect 426014 220046 426082 220102
rect 426138 220046 456678 220102
rect 456734 220046 456802 220102
rect 456858 220046 487398 220102
rect 487454 220046 487522 220102
rect 487578 220046 518118 220102
rect 518174 220046 518242 220102
rect 518298 220046 548838 220102
rect 548894 220046 548962 220102
rect 549018 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 364518 219978
rect 364574 219922 364642 219978
rect 364698 219922 395238 219978
rect 395294 219922 395362 219978
rect 395418 219922 425958 219978
rect 426014 219922 426082 219978
rect 426138 219922 456678 219978
rect 456734 219922 456802 219978
rect 456858 219922 487398 219978
rect 487454 219922 487522 219978
rect 487578 219922 518118 219978
rect 518174 219922 518242 219978
rect 518298 219922 548838 219978
rect 548894 219922 548962 219978
rect 549018 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect 192316 214498 289844 214514
rect 192316 214442 192332 214498
rect 192388 214442 289772 214498
rect 289828 214442 289844 214498
rect 192316 214426 289844 214442
rect 197916 214318 354468 214334
rect 197916 214262 197932 214318
rect 197988 214262 354396 214318
rect 354452 214262 354468 214318
rect 197916 214246 354468 214262
rect 187836 214138 359284 214154
rect 187836 214082 187852 214138
rect 187908 214082 359212 214138
rect 359268 214082 359284 214138
rect 187836 214066 359284 214082
rect 196460 211438 288164 211454
rect 196460 211382 196476 211438
rect 196532 211382 288092 211438
rect 288148 211382 288164 211438
rect 196460 211366 288164 211382
rect 199260 211258 315156 211274
rect 199260 211202 199276 211258
rect 199332 211202 315084 211258
rect 315140 211202 315156 211258
rect 199260 211186 315156 211202
rect 185484 211078 343044 211094
rect 185484 211022 185500 211078
rect 185556 211022 342972 211078
rect 343028 211022 343044 211078
rect 185484 211006 343044 211022
rect 197804 210898 355252 210914
rect 197804 210842 197820 210898
rect 197876 210842 355180 210898
rect 355236 210842 355252 210898
rect 197804 210826 355252 210842
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 39954 208350
rect 40010 208294 40078 208350
rect 40134 208294 40202 208350
rect 40258 208294 40326 208350
rect 40382 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 379878 208350
rect 379934 208294 380002 208350
rect 380058 208294 410598 208350
rect 410654 208294 410722 208350
rect 410778 208294 441318 208350
rect 441374 208294 441442 208350
rect 441498 208294 472038 208350
rect 472094 208294 472162 208350
rect 472218 208294 502758 208350
rect 502814 208294 502882 208350
rect 502938 208294 533478 208350
rect 533534 208294 533602 208350
rect 533658 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 39954 208226
rect 40010 208170 40078 208226
rect 40134 208170 40202 208226
rect 40258 208170 40326 208226
rect 40382 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 379878 208226
rect 379934 208170 380002 208226
rect 380058 208170 410598 208226
rect 410654 208170 410722 208226
rect 410778 208170 441318 208226
rect 441374 208170 441442 208226
rect 441498 208170 472038 208226
rect 472094 208170 472162 208226
rect 472218 208170 502758 208226
rect 502814 208170 502882 208226
rect 502938 208170 533478 208226
rect 533534 208170 533602 208226
rect 533658 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 39954 208102
rect 40010 208046 40078 208102
rect 40134 208046 40202 208102
rect 40258 208046 40326 208102
rect 40382 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 379878 208102
rect 379934 208046 380002 208102
rect 380058 208046 410598 208102
rect 410654 208046 410722 208102
rect 410778 208046 441318 208102
rect 441374 208046 441442 208102
rect 441498 208046 472038 208102
rect 472094 208046 472162 208102
rect 472218 208046 502758 208102
rect 502814 208046 502882 208102
rect 502938 208046 533478 208102
rect 533534 208046 533602 208102
rect 533658 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 39954 207978
rect 40010 207922 40078 207978
rect 40134 207922 40202 207978
rect 40258 207922 40326 207978
rect 40382 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 379878 207978
rect 379934 207922 380002 207978
rect 380058 207922 410598 207978
rect 410654 207922 410722 207978
rect 410778 207922 441318 207978
rect 441374 207922 441442 207978
rect 441498 207922 472038 207978
rect 472094 207922 472162 207978
rect 472218 207922 502758 207978
rect 502814 207922 502882 207978
rect 502938 207922 533478 207978
rect 533534 207922 533602 207978
rect 533658 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect 4156 206578 49716 206594
rect 4156 206522 4172 206578
rect 4228 206522 49644 206578
rect 49700 206522 49716 206578
rect 4156 206506 49716 206522
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 44518 202350
rect 44574 202294 44642 202350
rect 44698 202294 75238 202350
rect 75294 202294 75362 202350
rect 75418 202294 105958 202350
rect 106014 202294 106082 202350
rect 106138 202294 136678 202350
rect 136734 202294 136802 202350
rect 136858 202294 167398 202350
rect 167454 202294 167522 202350
rect 167578 202294 198118 202350
rect 198174 202294 198242 202350
rect 198298 202294 228838 202350
rect 228894 202294 228962 202350
rect 229018 202294 259558 202350
rect 259614 202294 259682 202350
rect 259738 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 364518 202350
rect 364574 202294 364642 202350
rect 364698 202294 395238 202350
rect 395294 202294 395362 202350
rect 395418 202294 425958 202350
rect 426014 202294 426082 202350
rect 426138 202294 456678 202350
rect 456734 202294 456802 202350
rect 456858 202294 487398 202350
rect 487454 202294 487522 202350
rect 487578 202294 518118 202350
rect 518174 202294 518242 202350
rect 518298 202294 548838 202350
rect 548894 202294 548962 202350
rect 549018 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 44518 202226
rect 44574 202170 44642 202226
rect 44698 202170 75238 202226
rect 75294 202170 75362 202226
rect 75418 202170 105958 202226
rect 106014 202170 106082 202226
rect 106138 202170 136678 202226
rect 136734 202170 136802 202226
rect 136858 202170 167398 202226
rect 167454 202170 167522 202226
rect 167578 202170 198118 202226
rect 198174 202170 198242 202226
rect 198298 202170 228838 202226
rect 228894 202170 228962 202226
rect 229018 202170 259558 202226
rect 259614 202170 259682 202226
rect 259738 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 364518 202226
rect 364574 202170 364642 202226
rect 364698 202170 395238 202226
rect 395294 202170 395362 202226
rect 395418 202170 425958 202226
rect 426014 202170 426082 202226
rect 426138 202170 456678 202226
rect 456734 202170 456802 202226
rect 456858 202170 487398 202226
rect 487454 202170 487522 202226
rect 487578 202170 518118 202226
rect 518174 202170 518242 202226
rect 518298 202170 548838 202226
rect 548894 202170 548962 202226
rect 549018 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 44518 202102
rect 44574 202046 44642 202102
rect 44698 202046 75238 202102
rect 75294 202046 75362 202102
rect 75418 202046 105958 202102
rect 106014 202046 106082 202102
rect 106138 202046 136678 202102
rect 136734 202046 136802 202102
rect 136858 202046 167398 202102
rect 167454 202046 167522 202102
rect 167578 202046 198118 202102
rect 198174 202046 198242 202102
rect 198298 202046 228838 202102
rect 228894 202046 228962 202102
rect 229018 202046 259558 202102
rect 259614 202046 259682 202102
rect 259738 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 364518 202102
rect 364574 202046 364642 202102
rect 364698 202046 395238 202102
rect 395294 202046 395362 202102
rect 395418 202046 425958 202102
rect 426014 202046 426082 202102
rect 426138 202046 456678 202102
rect 456734 202046 456802 202102
rect 456858 202046 487398 202102
rect 487454 202046 487522 202102
rect 487578 202046 518118 202102
rect 518174 202046 518242 202102
rect 518298 202046 548838 202102
rect 548894 202046 548962 202102
rect 549018 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 44518 201978
rect 44574 201922 44642 201978
rect 44698 201922 75238 201978
rect 75294 201922 75362 201978
rect 75418 201922 105958 201978
rect 106014 201922 106082 201978
rect 106138 201922 136678 201978
rect 136734 201922 136802 201978
rect 136858 201922 167398 201978
rect 167454 201922 167522 201978
rect 167578 201922 198118 201978
rect 198174 201922 198242 201978
rect 198298 201922 228838 201978
rect 228894 201922 228962 201978
rect 229018 201922 259558 201978
rect 259614 201922 259682 201978
rect 259738 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 364518 201978
rect 364574 201922 364642 201978
rect 364698 201922 395238 201978
rect 395294 201922 395362 201978
rect 395418 201922 425958 201978
rect 426014 201922 426082 201978
rect 426138 201922 456678 201978
rect 456734 201922 456802 201978
rect 456858 201922 487398 201978
rect 487454 201922 487522 201978
rect 487578 201922 518118 201978
rect 518174 201922 518242 201978
rect 518298 201922 548838 201978
rect 548894 201922 548962 201978
rect 549018 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect 345980 196678 350884 196694
rect 345980 196622 345996 196678
rect 346052 196622 350812 196678
rect 350868 196622 350884 196678
rect 345980 196606 350884 196622
rect 345420 195778 362196 195794
rect 345420 195722 345436 195778
rect 345492 195722 362124 195778
rect 362180 195722 362196 195778
rect 345420 195706 362196 195722
rect 339932 193978 361972 193994
rect 339932 193922 339948 193978
rect 340004 193922 361900 193978
rect 361956 193922 361972 193978
rect 339932 193906 361972 193922
rect 339260 193258 346404 193274
rect 339260 193202 339276 193258
rect 339332 193202 346332 193258
rect 346388 193202 346404 193258
rect 339260 193186 346404 193202
rect 344300 192718 351444 192734
rect 344300 192662 344316 192718
rect 344372 192662 351372 192718
rect 351428 192662 351444 192718
rect 344300 192646 351444 192662
rect 341836 192538 352788 192554
rect 341836 192482 341852 192538
rect 341908 192482 352716 192538
rect 352772 192482 352788 192538
rect 341836 192466 352788 192482
rect 345308 192358 358612 192374
rect 345308 192302 345324 192358
rect 345380 192302 358540 192358
rect 358596 192302 358612 192358
rect 345308 192286 358612 192302
rect 344860 191818 347076 191834
rect 344860 191762 344876 191818
rect 344932 191762 347004 191818
rect 347060 191762 347076 191818
rect 344860 191746 347076 191762
rect 359756 191818 360628 191834
rect 359756 191762 359772 191818
rect 359828 191762 360556 191818
rect 360612 191762 360628 191818
rect 359756 191746 360628 191762
rect 344076 191638 346292 191654
rect 344076 191582 344092 191638
rect 344148 191582 346220 191638
rect 346276 191582 346292 191638
rect 344076 191566 346292 191582
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 39954 190350
rect 40010 190294 40078 190350
rect 40134 190294 40202 190350
rect 40258 190294 40326 190350
rect 40382 190294 59878 190350
rect 59934 190294 60002 190350
rect 60058 190294 90598 190350
rect 90654 190294 90722 190350
rect 90778 190294 121318 190350
rect 121374 190294 121442 190350
rect 121498 190294 152038 190350
rect 152094 190294 152162 190350
rect 152218 190294 182758 190350
rect 182814 190294 182882 190350
rect 182938 190294 213478 190350
rect 213534 190294 213602 190350
rect 213658 190294 244198 190350
rect 244254 190294 244322 190350
rect 244378 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 319822 190350
rect 319878 190294 319946 190350
rect 320002 190294 328390 190350
rect 328446 190294 328514 190350
rect 328570 190294 336958 190350
rect 337014 190294 337082 190350
rect 337138 190294 345526 190350
rect 345582 190294 345650 190350
rect 345706 190294 379878 190350
rect 379934 190294 380002 190350
rect 380058 190294 410598 190350
rect 410654 190294 410722 190350
rect 410778 190294 441318 190350
rect 441374 190294 441442 190350
rect 441498 190294 472038 190350
rect 472094 190294 472162 190350
rect 472218 190294 502758 190350
rect 502814 190294 502882 190350
rect 502938 190294 533478 190350
rect 533534 190294 533602 190350
rect 533658 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 39954 190226
rect 40010 190170 40078 190226
rect 40134 190170 40202 190226
rect 40258 190170 40326 190226
rect 40382 190170 59878 190226
rect 59934 190170 60002 190226
rect 60058 190170 90598 190226
rect 90654 190170 90722 190226
rect 90778 190170 121318 190226
rect 121374 190170 121442 190226
rect 121498 190170 152038 190226
rect 152094 190170 152162 190226
rect 152218 190170 182758 190226
rect 182814 190170 182882 190226
rect 182938 190170 213478 190226
rect 213534 190170 213602 190226
rect 213658 190170 244198 190226
rect 244254 190170 244322 190226
rect 244378 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 319822 190226
rect 319878 190170 319946 190226
rect 320002 190170 328390 190226
rect 328446 190170 328514 190226
rect 328570 190170 336958 190226
rect 337014 190170 337082 190226
rect 337138 190170 345526 190226
rect 345582 190170 345650 190226
rect 345706 190170 379878 190226
rect 379934 190170 380002 190226
rect 380058 190170 410598 190226
rect 410654 190170 410722 190226
rect 410778 190170 441318 190226
rect 441374 190170 441442 190226
rect 441498 190170 472038 190226
rect 472094 190170 472162 190226
rect 472218 190170 502758 190226
rect 502814 190170 502882 190226
rect 502938 190170 533478 190226
rect 533534 190170 533602 190226
rect 533658 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 39954 190102
rect 40010 190046 40078 190102
rect 40134 190046 40202 190102
rect 40258 190046 40326 190102
rect 40382 190046 59878 190102
rect 59934 190046 60002 190102
rect 60058 190046 90598 190102
rect 90654 190046 90722 190102
rect 90778 190046 121318 190102
rect 121374 190046 121442 190102
rect 121498 190046 152038 190102
rect 152094 190046 152162 190102
rect 152218 190046 182758 190102
rect 182814 190046 182882 190102
rect 182938 190046 213478 190102
rect 213534 190046 213602 190102
rect 213658 190046 244198 190102
rect 244254 190046 244322 190102
rect 244378 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 319822 190102
rect 319878 190046 319946 190102
rect 320002 190046 328390 190102
rect 328446 190046 328514 190102
rect 328570 190046 336958 190102
rect 337014 190046 337082 190102
rect 337138 190046 345526 190102
rect 345582 190046 345650 190102
rect 345706 190046 379878 190102
rect 379934 190046 380002 190102
rect 380058 190046 410598 190102
rect 410654 190046 410722 190102
rect 410778 190046 441318 190102
rect 441374 190046 441442 190102
rect 441498 190046 472038 190102
rect 472094 190046 472162 190102
rect 472218 190046 502758 190102
rect 502814 190046 502882 190102
rect 502938 190046 533478 190102
rect 533534 190046 533602 190102
rect 533658 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 39954 189978
rect 40010 189922 40078 189978
rect 40134 189922 40202 189978
rect 40258 189922 40326 189978
rect 40382 189922 59878 189978
rect 59934 189922 60002 189978
rect 60058 189922 90598 189978
rect 90654 189922 90722 189978
rect 90778 189922 121318 189978
rect 121374 189922 121442 189978
rect 121498 189922 152038 189978
rect 152094 189922 152162 189978
rect 152218 189922 182758 189978
rect 182814 189922 182882 189978
rect 182938 189922 213478 189978
rect 213534 189922 213602 189978
rect 213658 189922 244198 189978
rect 244254 189922 244322 189978
rect 244378 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 319822 189978
rect 319878 189922 319946 189978
rect 320002 189922 328390 189978
rect 328446 189922 328514 189978
rect 328570 189922 336958 189978
rect 337014 189922 337082 189978
rect 337138 189922 345526 189978
rect 345582 189922 345650 189978
rect 345706 189922 379878 189978
rect 379934 189922 380002 189978
rect 380058 189922 410598 189978
rect 410654 189922 410722 189978
rect 410778 189922 441318 189978
rect 441374 189922 441442 189978
rect 441498 189922 472038 189978
rect 472094 189922 472162 189978
rect 472218 189922 502758 189978
rect 502814 189922 502882 189978
rect 502938 189922 533478 189978
rect 533534 189922 533602 189978
rect 533658 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect 359756 186058 359844 186074
rect 359756 186002 359772 186058
rect 359828 186002 359844 186058
rect 359756 185894 359844 186002
rect 359756 185878 360068 185894
rect 359756 185822 359996 185878
rect 360052 185822 360068 185878
rect 359756 185806 360068 185822
rect 359756 185698 360292 185714
rect 359756 185642 359772 185698
rect 359828 185642 360220 185698
rect 360276 185642 360292 185698
rect 359756 185626 360292 185642
rect 361212 184618 361972 184634
rect 361212 184562 361228 184618
rect 361284 184562 361900 184618
rect 361956 184562 361972 184618
rect 361212 184546 361972 184562
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 44518 184350
rect 44574 184294 44642 184350
rect 44698 184294 75238 184350
rect 75294 184294 75362 184350
rect 75418 184294 105958 184350
rect 106014 184294 106082 184350
rect 106138 184294 136678 184350
rect 136734 184294 136802 184350
rect 136858 184294 167398 184350
rect 167454 184294 167522 184350
rect 167578 184294 198118 184350
rect 198174 184294 198242 184350
rect 198298 184294 228838 184350
rect 228894 184294 228962 184350
rect 229018 184294 259558 184350
rect 259614 184294 259682 184350
rect 259738 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 315538 184350
rect 315594 184294 315662 184350
rect 315718 184294 324106 184350
rect 324162 184294 324230 184350
rect 324286 184294 332674 184350
rect 332730 184294 332798 184350
rect 332854 184294 341242 184350
rect 341298 184294 341366 184350
rect 341422 184294 364518 184350
rect 364574 184294 364642 184350
rect 364698 184294 395238 184350
rect 395294 184294 395362 184350
rect 395418 184294 425958 184350
rect 426014 184294 426082 184350
rect 426138 184294 456678 184350
rect 456734 184294 456802 184350
rect 456858 184294 487398 184350
rect 487454 184294 487522 184350
rect 487578 184294 518118 184350
rect 518174 184294 518242 184350
rect 518298 184294 548838 184350
rect 548894 184294 548962 184350
rect 549018 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 44518 184226
rect 44574 184170 44642 184226
rect 44698 184170 75238 184226
rect 75294 184170 75362 184226
rect 75418 184170 105958 184226
rect 106014 184170 106082 184226
rect 106138 184170 136678 184226
rect 136734 184170 136802 184226
rect 136858 184170 167398 184226
rect 167454 184170 167522 184226
rect 167578 184170 198118 184226
rect 198174 184170 198242 184226
rect 198298 184170 228838 184226
rect 228894 184170 228962 184226
rect 229018 184170 259558 184226
rect 259614 184170 259682 184226
rect 259738 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 315538 184226
rect 315594 184170 315662 184226
rect 315718 184170 324106 184226
rect 324162 184170 324230 184226
rect 324286 184170 332674 184226
rect 332730 184170 332798 184226
rect 332854 184170 341242 184226
rect 341298 184170 341366 184226
rect 341422 184170 364518 184226
rect 364574 184170 364642 184226
rect 364698 184170 395238 184226
rect 395294 184170 395362 184226
rect 395418 184170 425958 184226
rect 426014 184170 426082 184226
rect 426138 184170 456678 184226
rect 456734 184170 456802 184226
rect 456858 184170 487398 184226
rect 487454 184170 487522 184226
rect 487578 184170 518118 184226
rect 518174 184170 518242 184226
rect 518298 184170 548838 184226
rect 548894 184170 548962 184226
rect 549018 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 44518 184102
rect 44574 184046 44642 184102
rect 44698 184046 75238 184102
rect 75294 184046 75362 184102
rect 75418 184046 105958 184102
rect 106014 184046 106082 184102
rect 106138 184046 136678 184102
rect 136734 184046 136802 184102
rect 136858 184046 167398 184102
rect 167454 184046 167522 184102
rect 167578 184046 198118 184102
rect 198174 184046 198242 184102
rect 198298 184046 228838 184102
rect 228894 184046 228962 184102
rect 229018 184046 259558 184102
rect 259614 184046 259682 184102
rect 259738 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 315538 184102
rect 315594 184046 315662 184102
rect 315718 184046 324106 184102
rect 324162 184046 324230 184102
rect 324286 184046 332674 184102
rect 332730 184046 332798 184102
rect 332854 184046 341242 184102
rect 341298 184046 341366 184102
rect 341422 184046 364518 184102
rect 364574 184046 364642 184102
rect 364698 184046 395238 184102
rect 395294 184046 395362 184102
rect 395418 184046 425958 184102
rect 426014 184046 426082 184102
rect 426138 184046 456678 184102
rect 456734 184046 456802 184102
rect 456858 184046 487398 184102
rect 487454 184046 487522 184102
rect 487578 184046 518118 184102
rect 518174 184046 518242 184102
rect 518298 184046 548838 184102
rect 548894 184046 548962 184102
rect 549018 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 44518 183978
rect 44574 183922 44642 183978
rect 44698 183922 75238 183978
rect 75294 183922 75362 183978
rect 75418 183922 105958 183978
rect 106014 183922 106082 183978
rect 106138 183922 136678 183978
rect 136734 183922 136802 183978
rect 136858 183922 167398 183978
rect 167454 183922 167522 183978
rect 167578 183922 198118 183978
rect 198174 183922 198242 183978
rect 198298 183922 228838 183978
rect 228894 183922 228962 183978
rect 229018 183922 259558 183978
rect 259614 183922 259682 183978
rect 259738 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 315538 183978
rect 315594 183922 315662 183978
rect 315718 183922 324106 183978
rect 324162 183922 324230 183978
rect 324286 183922 332674 183978
rect 332730 183922 332798 183978
rect 332854 183922 341242 183978
rect 341298 183922 341366 183978
rect 341422 183922 364518 183978
rect 364574 183922 364642 183978
rect 364698 183922 395238 183978
rect 395294 183922 395362 183978
rect 395418 183922 425958 183978
rect 426014 183922 426082 183978
rect 426138 183922 456678 183978
rect 456734 183922 456802 183978
rect 456858 183922 487398 183978
rect 487454 183922 487522 183978
rect 487578 183922 518118 183978
rect 518174 183922 518242 183978
rect 518298 183922 548838 183978
rect 548894 183922 548962 183978
rect 549018 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect 356956 181018 361636 181034
rect 356956 180962 356972 181018
rect 357028 180962 361564 181018
rect 361620 180962 361636 181018
rect 356956 180946 361636 180962
rect 359196 176338 361524 176354
rect 359196 176282 359212 176338
rect 359268 176282 361452 176338
rect 361508 176282 361524 176338
rect 359196 176266 361524 176282
rect 345868 175258 375300 175274
rect 345868 175202 345884 175258
rect 345940 175202 375228 175258
rect 375284 175202 375300 175258
rect 345868 175186 375300 175202
rect 345196 173998 417636 174014
rect 345196 173942 345212 173998
rect 345268 173942 417564 173998
rect 417620 173942 417636 173998
rect 345196 173926 417636 173942
rect 346988 173818 561220 173834
rect 346988 173762 347004 173818
rect 347060 173762 561148 173818
rect 561204 173762 561220 173818
rect 346988 173746 561220 173762
rect 358412 173098 490660 173114
rect 358412 173042 358428 173098
rect 358484 173042 490588 173098
rect 490644 173042 490660 173098
rect 358412 173026 490660 173042
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 59878 172350
rect 59934 172294 60002 172350
rect 60058 172294 90598 172350
rect 90654 172294 90722 172350
rect 90778 172294 121318 172350
rect 121374 172294 121442 172350
rect 121498 172294 152038 172350
rect 152094 172294 152162 172350
rect 152218 172294 182758 172350
rect 182814 172294 182882 172350
rect 182938 172294 213478 172350
rect 213534 172294 213602 172350
rect 213658 172294 244198 172350
rect 244254 172294 244322 172350
rect 244378 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 319822 172350
rect 319878 172294 319946 172350
rect 320002 172294 328390 172350
rect 328446 172294 328514 172350
rect 328570 172294 336958 172350
rect 337014 172294 337082 172350
rect 337138 172294 345526 172350
rect 345582 172294 345650 172350
rect 345706 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 408594 172350
rect 408650 172294 408718 172350
rect 408774 172294 408842 172350
rect 408898 172294 408966 172350
rect 409022 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 59878 172226
rect 59934 172170 60002 172226
rect 60058 172170 90598 172226
rect 90654 172170 90722 172226
rect 90778 172170 121318 172226
rect 121374 172170 121442 172226
rect 121498 172170 152038 172226
rect 152094 172170 152162 172226
rect 152218 172170 182758 172226
rect 182814 172170 182882 172226
rect 182938 172170 213478 172226
rect 213534 172170 213602 172226
rect 213658 172170 244198 172226
rect 244254 172170 244322 172226
rect 244378 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 319822 172226
rect 319878 172170 319946 172226
rect 320002 172170 328390 172226
rect 328446 172170 328514 172226
rect 328570 172170 336958 172226
rect 337014 172170 337082 172226
rect 337138 172170 345526 172226
rect 345582 172170 345650 172226
rect 345706 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 408594 172226
rect 408650 172170 408718 172226
rect 408774 172170 408842 172226
rect 408898 172170 408966 172226
rect 409022 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 59878 172102
rect 59934 172046 60002 172102
rect 60058 172046 90598 172102
rect 90654 172046 90722 172102
rect 90778 172046 121318 172102
rect 121374 172046 121442 172102
rect 121498 172046 152038 172102
rect 152094 172046 152162 172102
rect 152218 172046 182758 172102
rect 182814 172046 182882 172102
rect 182938 172046 213478 172102
rect 213534 172046 213602 172102
rect 213658 172046 244198 172102
rect 244254 172046 244322 172102
rect 244378 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 319822 172102
rect 319878 172046 319946 172102
rect 320002 172046 328390 172102
rect 328446 172046 328514 172102
rect 328570 172046 336958 172102
rect 337014 172046 337082 172102
rect 337138 172046 345526 172102
rect 345582 172046 345650 172102
rect 345706 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 408594 172102
rect 408650 172046 408718 172102
rect 408774 172046 408842 172102
rect 408898 172046 408966 172102
rect 409022 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 59878 171978
rect 59934 171922 60002 171978
rect 60058 171922 90598 171978
rect 90654 171922 90722 171978
rect 90778 171922 121318 171978
rect 121374 171922 121442 171978
rect 121498 171922 152038 171978
rect 152094 171922 152162 171978
rect 152218 171922 182758 171978
rect 182814 171922 182882 171978
rect 182938 171922 213478 171978
rect 213534 171922 213602 171978
rect 213658 171922 244198 171978
rect 244254 171922 244322 171978
rect 244378 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 319822 171978
rect 319878 171922 319946 171978
rect 320002 171922 328390 171978
rect 328446 171922 328514 171978
rect 328570 171922 336958 171978
rect 337014 171922 337082 171978
rect 337138 171922 345526 171978
rect 345582 171922 345650 171978
rect 345706 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 408594 171978
rect 408650 171922 408718 171978
rect 408774 171922 408842 171978
rect 408898 171922 408966 171978
rect 409022 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect 350796 170578 559652 170594
rect 350796 170522 350812 170578
rect 350868 170522 559580 170578
rect 559636 170522 559652 170578
rect 350796 170506 559652 170522
rect 358748 168778 488980 168794
rect 358748 168722 358764 168778
rect 358820 168722 488908 168778
rect 488964 168722 488980 168778
rect 358748 168706 488980 168722
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 44518 166350
rect 44574 166294 44642 166350
rect 44698 166294 75238 166350
rect 75294 166294 75362 166350
rect 75418 166294 105958 166350
rect 106014 166294 106082 166350
rect 106138 166294 136678 166350
rect 136734 166294 136802 166350
rect 136858 166294 167398 166350
rect 167454 166294 167522 166350
rect 167578 166294 198118 166350
rect 198174 166294 198242 166350
rect 198298 166294 228838 166350
rect 228894 166294 228962 166350
rect 229018 166294 259558 166350
rect 259614 166294 259682 166350
rect 259738 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 315538 166350
rect 315594 166294 315662 166350
rect 315718 166294 324106 166350
rect 324162 166294 324230 166350
rect 324286 166294 332674 166350
rect 332730 166294 332798 166350
rect 332854 166294 341242 166350
rect 341298 166294 341366 166350
rect 341422 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 404874 166350
rect 404930 166294 404998 166350
rect 405054 166294 405122 166350
rect 405178 166294 405246 166350
rect 405302 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 44518 166226
rect 44574 166170 44642 166226
rect 44698 166170 75238 166226
rect 75294 166170 75362 166226
rect 75418 166170 105958 166226
rect 106014 166170 106082 166226
rect 106138 166170 136678 166226
rect 136734 166170 136802 166226
rect 136858 166170 167398 166226
rect 167454 166170 167522 166226
rect 167578 166170 198118 166226
rect 198174 166170 198242 166226
rect 198298 166170 228838 166226
rect 228894 166170 228962 166226
rect 229018 166170 259558 166226
rect 259614 166170 259682 166226
rect 259738 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 315538 166226
rect 315594 166170 315662 166226
rect 315718 166170 324106 166226
rect 324162 166170 324230 166226
rect 324286 166170 332674 166226
rect 332730 166170 332798 166226
rect 332854 166170 341242 166226
rect 341298 166170 341366 166226
rect 341422 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 404874 166226
rect 404930 166170 404998 166226
rect 405054 166170 405122 166226
rect 405178 166170 405246 166226
rect 405302 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 44518 166102
rect 44574 166046 44642 166102
rect 44698 166046 75238 166102
rect 75294 166046 75362 166102
rect 75418 166046 105958 166102
rect 106014 166046 106082 166102
rect 106138 166046 136678 166102
rect 136734 166046 136802 166102
rect 136858 166046 167398 166102
rect 167454 166046 167522 166102
rect 167578 166046 198118 166102
rect 198174 166046 198242 166102
rect 198298 166046 228838 166102
rect 228894 166046 228962 166102
rect 229018 166046 259558 166102
rect 259614 166046 259682 166102
rect 259738 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 315538 166102
rect 315594 166046 315662 166102
rect 315718 166046 324106 166102
rect 324162 166046 324230 166102
rect 324286 166046 332674 166102
rect 332730 166046 332798 166102
rect 332854 166046 341242 166102
rect 341298 166046 341366 166102
rect 341422 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 404874 166102
rect 404930 166046 404998 166102
rect 405054 166046 405122 166102
rect 405178 166046 405246 166102
rect 405302 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 44518 165978
rect 44574 165922 44642 165978
rect 44698 165922 75238 165978
rect 75294 165922 75362 165978
rect 75418 165922 105958 165978
rect 106014 165922 106082 165978
rect 106138 165922 136678 165978
rect 136734 165922 136802 165978
rect 136858 165922 167398 165978
rect 167454 165922 167522 165978
rect 167578 165922 198118 165978
rect 198174 165922 198242 165978
rect 198298 165922 228838 165978
rect 228894 165922 228962 165978
rect 229018 165922 259558 165978
rect 259614 165922 259682 165978
rect 259738 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 315538 165978
rect 315594 165922 315662 165978
rect 315718 165922 324106 165978
rect 324162 165922 324230 165978
rect 324286 165922 332674 165978
rect 332730 165922 332798 165978
rect 332854 165922 341242 165978
rect 341298 165922 341366 165978
rect 341422 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 404874 165978
rect 404930 165922 404998 165978
rect 405054 165922 405122 165978
rect 405178 165922 405246 165978
rect 405302 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect 4156 164638 49604 164654
rect 4156 164582 4172 164638
rect 4228 164582 49532 164638
rect 49588 164582 49604 164638
rect 4156 164566 49604 164582
rect 298940 160678 566260 160694
rect 298940 160622 298956 160678
rect 299012 160622 566188 160678
rect 566244 160622 566260 160678
rect 298940 160606 566260 160622
rect 293788 160498 564692 160514
rect 293788 160442 293804 160498
rect 293860 160442 564620 160498
rect 564676 160442 564692 160498
rect 293788 160426 564692 160442
rect 300620 158878 561332 158894
rect 300620 158822 300636 158878
rect 300692 158822 561260 158878
rect 561316 158822 561332 158878
rect 300620 158806 561332 158822
rect 293900 158698 564580 158714
rect 293900 158642 293916 158698
rect 293972 158642 564508 158698
rect 564564 158642 564580 158698
rect 293900 158626 564580 158642
rect 324364 157798 349540 157814
rect 324364 157742 324380 157798
rect 324436 157742 349468 157798
rect 349524 157742 349540 157798
rect 324364 157726 349540 157742
rect 330636 157618 346180 157634
rect 330636 157562 330652 157618
rect 330708 157562 346108 157618
rect 346164 157562 346180 157618
rect 330636 157546 346180 157562
rect 332204 157438 347860 157454
rect 332204 157382 332220 157438
rect 332276 157382 347788 157438
rect 347844 157382 347860 157438
rect 332204 157366 347860 157382
rect 360092 157078 493236 157094
rect 360092 157022 360108 157078
rect 360164 157022 493164 157078
rect 493220 157022 493236 157078
rect 360092 157006 493236 157022
rect 295580 155458 564804 155474
rect 295580 155402 295596 155458
rect 295652 155402 564732 155458
rect 564788 155402 564804 155458
rect 295580 155386 564804 155402
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 59878 154350
rect 59934 154294 60002 154350
rect 60058 154294 90598 154350
rect 90654 154294 90722 154350
rect 90778 154294 121318 154350
rect 121374 154294 121442 154350
rect 121498 154294 152038 154350
rect 152094 154294 152162 154350
rect 152218 154294 182758 154350
rect 182814 154294 182882 154350
rect 182938 154294 213478 154350
rect 213534 154294 213602 154350
rect 213658 154294 244198 154350
rect 244254 154294 244322 154350
rect 244378 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 59878 154226
rect 59934 154170 60002 154226
rect 60058 154170 90598 154226
rect 90654 154170 90722 154226
rect 90778 154170 121318 154226
rect 121374 154170 121442 154226
rect 121498 154170 152038 154226
rect 152094 154170 152162 154226
rect 152218 154170 182758 154226
rect 182814 154170 182882 154226
rect 182938 154170 213478 154226
rect 213534 154170 213602 154226
rect 213658 154170 244198 154226
rect 244254 154170 244322 154226
rect 244378 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 59878 154102
rect 59934 154046 60002 154102
rect 60058 154046 90598 154102
rect 90654 154046 90722 154102
rect 90778 154046 121318 154102
rect 121374 154046 121442 154102
rect 121498 154046 152038 154102
rect 152094 154046 152162 154102
rect 152218 154046 182758 154102
rect 182814 154046 182882 154102
rect 182938 154046 213478 154102
rect 213534 154046 213602 154102
rect 213658 154046 244198 154102
rect 244254 154046 244322 154102
rect 244378 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 59878 153978
rect 59934 153922 60002 153978
rect 60058 153922 90598 153978
rect 90654 153922 90722 153978
rect 90778 153922 121318 153978
rect 121374 153922 121442 153978
rect 121498 153922 152038 153978
rect 152094 153922 152162 153978
rect 152218 153922 182758 153978
rect 182814 153922 182882 153978
rect 182938 153922 213478 153978
rect 213534 153922 213602 153978
rect 213658 153922 244198 153978
rect 244254 153922 244322 153978
rect 244378 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect 272508 153658 502644 153674
rect 272508 153602 272524 153658
rect 272580 153602 502572 153658
rect 502628 153602 502644 153658
rect 272508 153586 502644 153602
rect 356172 153478 503204 153494
rect 356172 153422 356188 153478
rect 356244 153422 503132 153478
rect 503188 153422 503204 153478
rect 356172 153406 503204 153422
rect 352924 150598 482148 150614
rect 352924 150542 352940 150598
rect 352996 150542 482076 150598
rect 482132 150542 482148 150598
rect 352924 150526 482148 150542
rect 277996 150418 590564 150434
rect 277996 150362 278012 150418
rect 278068 150362 590492 150418
rect 590548 150362 590564 150418
rect 277996 150346 590564 150362
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 44518 148350
rect 44574 148294 44642 148350
rect 44698 148294 75238 148350
rect 75294 148294 75362 148350
rect 75418 148294 105958 148350
rect 106014 148294 106082 148350
rect 106138 148294 136678 148350
rect 136734 148294 136802 148350
rect 136858 148294 167398 148350
rect 167454 148294 167522 148350
rect 167578 148294 198118 148350
rect 198174 148294 198242 148350
rect 198298 148294 228838 148350
rect 228894 148294 228962 148350
rect 229018 148294 259558 148350
rect 259614 148294 259682 148350
rect 259738 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 44518 148226
rect 44574 148170 44642 148226
rect 44698 148170 75238 148226
rect 75294 148170 75362 148226
rect 75418 148170 105958 148226
rect 106014 148170 106082 148226
rect 106138 148170 136678 148226
rect 136734 148170 136802 148226
rect 136858 148170 167398 148226
rect 167454 148170 167522 148226
rect 167578 148170 198118 148226
rect 198174 148170 198242 148226
rect 198298 148170 228838 148226
rect 228894 148170 228962 148226
rect 229018 148170 259558 148226
rect 259614 148170 259682 148226
rect 259738 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 44518 148102
rect 44574 148046 44642 148102
rect 44698 148046 75238 148102
rect 75294 148046 75362 148102
rect 75418 148046 105958 148102
rect 106014 148046 106082 148102
rect 106138 148046 136678 148102
rect 136734 148046 136802 148102
rect 136858 148046 167398 148102
rect 167454 148046 167522 148102
rect 167578 148046 198118 148102
rect 198174 148046 198242 148102
rect 198298 148046 228838 148102
rect 228894 148046 228962 148102
rect 229018 148046 259558 148102
rect 259614 148046 259682 148102
rect 259738 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 44518 147978
rect 44574 147922 44642 147978
rect 44698 147922 75238 147978
rect 75294 147922 75362 147978
rect 75418 147922 105958 147978
rect 106014 147922 106082 147978
rect 106138 147922 136678 147978
rect 136734 147922 136802 147978
rect 136858 147922 167398 147978
rect 167454 147922 167522 147978
rect 167578 147922 198118 147978
rect 198174 147922 198242 147978
rect 198298 147922 228838 147978
rect 228894 147922 228962 147978
rect 229018 147922 259558 147978
rect 259614 147922 259682 147978
rect 259738 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect 357404 147718 463444 147734
rect 357404 147662 357420 147718
rect 357476 147662 463372 147718
rect 463428 147662 463444 147718
rect 357404 147646 463444 147662
rect 330076 146998 357492 147014
rect 330076 146942 330092 146998
rect 330148 146942 357420 146998
rect 357476 146942 357492 146998
rect 330076 146926 357492 146942
rect 307340 146098 462100 146114
rect 307340 146042 307356 146098
rect 307412 146042 462028 146098
rect 462084 146042 462100 146098
rect 307340 146026 462100 146042
rect 268588 136918 415060 136934
rect 268588 136862 268604 136918
rect 268660 136862 414988 136918
rect 415044 136862 415060 136918
rect 268588 136846 415060 136862
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 39954 136350
rect 40010 136294 40078 136350
rect 40134 136294 40202 136350
rect 40258 136294 40326 136350
rect 40382 136294 59878 136350
rect 59934 136294 60002 136350
rect 60058 136294 90598 136350
rect 90654 136294 90722 136350
rect 90778 136294 121318 136350
rect 121374 136294 121442 136350
rect 121498 136294 152038 136350
rect 152094 136294 152162 136350
rect 152218 136294 182758 136350
rect 182814 136294 182882 136350
rect 182938 136294 213478 136350
rect 213534 136294 213602 136350
rect 213658 136294 244198 136350
rect 244254 136294 244322 136350
rect 244378 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 479878 136350
rect 479934 136294 480002 136350
rect 480058 136294 510598 136350
rect 510654 136294 510722 136350
rect 510778 136294 541318 136350
rect 541374 136294 541442 136350
rect 541498 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 39954 136226
rect 40010 136170 40078 136226
rect 40134 136170 40202 136226
rect 40258 136170 40326 136226
rect 40382 136170 59878 136226
rect 59934 136170 60002 136226
rect 60058 136170 90598 136226
rect 90654 136170 90722 136226
rect 90778 136170 121318 136226
rect 121374 136170 121442 136226
rect 121498 136170 152038 136226
rect 152094 136170 152162 136226
rect 152218 136170 182758 136226
rect 182814 136170 182882 136226
rect 182938 136170 213478 136226
rect 213534 136170 213602 136226
rect 213658 136170 244198 136226
rect 244254 136170 244322 136226
rect 244378 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 479878 136226
rect 479934 136170 480002 136226
rect 480058 136170 510598 136226
rect 510654 136170 510722 136226
rect 510778 136170 541318 136226
rect 541374 136170 541442 136226
rect 541498 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 39954 136102
rect 40010 136046 40078 136102
rect 40134 136046 40202 136102
rect 40258 136046 40326 136102
rect 40382 136046 59878 136102
rect 59934 136046 60002 136102
rect 60058 136046 90598 136102
rect 90654 136046 90722 136102
rect 90778 136046 121318 136102
rect 121374 136046 121442 136102
rect 121498 136046 152038 136102
rect 152094 136046 152162 136102
rect 152218 136046 182758 136102
rect 182814 136046 182882 136102
rect 182938 136046 213478 136102
rect 213534 136046 213602 136102
rect 213658 136046 244198 136102
rect 244254 136046 244322 136102
rect 244378 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 479878 136102
rect 479934 136046 480002 136102
rect 480058 136046 510598 136102
rect 510654 136046 510722 136102
rect 510778 136046 541318 136102
rect 541374 136046 541442 136102
rect 541498 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 39954 135978
rect 40010 135922 40078 135978
rect 40134 135922 40202 135978
rect 40258 135922 40326 135978
rect 40382 135922 59878 135978
rect 59934 135922 60002 135978
rect 60058 135922 90598 135978
rect 90654 135922 90722 135978
rect 90778 135922 121318 135978
rect 121374 135922 121442 135978
rect 121498 135922 152038 135978
rect 152094 135922 152162 135978
rect 152218 135922 182758 135978
rect 182814 135922 182882 135978
rect 182938 135922 213478 135978
rect 213534 135922 213602 135978
rect 213658 135922 244198 135978
rect 244254 135922 244322 135978
rect 244378 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 479878 135978
rect 479934 135922 480002 135978
rect 480058 135922 510598 135978
rect 510654 135922 510722 135978
rect 510778 135922 541318 135978
rect 541374 135922 541442 135978
rect 541498 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect 268700 133498 411700 133514
rect 268700 133442 268716 133498
rect 268772 133442 411628 133498
rect 411684 133442 411700 133498
rect 268700 133426 411700 133442
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 44518 130350
rect 44574 130294 44642 130350
rect 44698 130294 75238 130350
rect 75294 130294 75362 130350
rect 75418 130294 105958 130350
rect 106014 130294 106082 130350
rect 106138 130294 136678 130350
rect 136734 130294 136802 130350
rect 136858 130294 167398 130350
rect 167454 130294 167522 130350
rect 167578 130294 198118 130350
rect 198174 130294 198242 130350
rect 198298 130294 228838 130350
rect 228894 130294 228962 130350
rect 229018 130294 259558 130350
rect 259614 130294 259682 130350
rect 259738 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 464518 130350
rect 464574 130294 464642 130350
rect 464698 130294 495238 130350
rect 495294 130294 495362 130350
rect 495418 130294 525958 130350
rect 526014 130294 526082 130350
rect 526138 130294 556678 130350
rect 556734 130294 556802 130350
rect 556858 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 44518 130226
rect 44574 130170 44642 130226
rect 44698 130170 75238 130226
rect 75294 130170 75362 130226
rect 75418 130170 105958 130226
rect 106014 130170 106082 130226
rect 106138 130170 136678 130226
rect 136734 130170 136802 130226
rect 136858 130170 167398 130226
rect 167454 130170 167522 130226
rect 167578 130170 198118 130226
rect 198174 130170 198242 130226
rect 198298 130170 228838 130226
rect 228894 130170 228962 130226
rect 229018 130170 259558 130226
rect 259614 130170 259682 130226
rect 259738 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 464518 130226
rect 464574 130170 464642 130226
rect 464698 130170 495238 130226
rect 495294 130170 495362 130226
rect 495418 130170 525958 130226
rect 526014 130170 526082 130226
rect 526138 130170 556678 130226
rect 556734 130170 556802 130226
rect 556858 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 44518 130102
rect 44574 130046 44642 130102
rect 44698 130046 75238 130102
rect 75294 130046 75362 130102
rect 75418 130046 105958 130102
rect 106014 130046 106082 130102
rect 106138 130046 136678 130102
rect 136734 130046 136802 130102
rect 136858 130046 167398 130102
rect 167454 130046 167522 130102
rect 167578 130046 198118 130102
rect 198174 130046 198242 130102
rect 198298 130046 228838 130102
rect 228894 130046 228962 130102
rect 229018 130046 259558 130102
rect 259614 130046 259682 130102
rect 259738 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 464518 130102
rect 464574 130046 464642 130102
rect 464698 130046 495238 130102
rect 495294 130046 495362 130102
rect 495418 130046 525958 130102
rect 526014 130046 526082 130102
rect 526138 130046 556678 130102
rect 556734 130046 556802 130102
rect 556858 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 44518 129978
rect 44574 129922 44642 129978
rect 44698 129922 75238 129978
rect 75294 129922 75362 129978
rect 75418 129922 105958 129978
rect 106014 129922 106082 129978
rect 106138 129922 136678 129978
rect 136734 129922 136802 129978
rect 136858 129922 167398 129978
rect 167454 129922 167522 129978
rect 167578 129922 198118 129978
rect 198174 129922 198242 129978
rect 198298 129922 228838 129978
rect 228894 129922 228962 129978
rect 229018 129922 259558 129978
rect 259614 129922 259682 129978
rect 259738 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 464518 129978
rect 464574 129922 464642 129978
rect 464698 129922 495238 129978
rect 495294 129922 495362 129978
rect 495418 129922 525958 129978
rect 526014 129922 526082 129978
rect 526138 129922 556678 129978
rect 556734 129922 556802 129978
rect 556858 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect 298156 124318 395012 124334
rect 298156 124262 298172 124318
rect 298228 124262 394940 124318
rect 394996 124262 395012 124318
rect 298156 124246 395012 124262
rect 304876 124138 388964 124154
rect 304876 124082 304892 124138
rect 304948 124082 388892 124138
rect 388948 124082 388964 124138
rect 304876 124066 388964 124082
rect 306556 123958 390980 123974
rect 306556 123902 306572 123958
rect 306628 123902 390908 123958
rect 390964 123902 390980 123958
rect 306556 123886 390980 123902
rect 308236 123778 386948 123794
rect 308236 123722 308252 123778
rect 308308 123722 386876 123778
rect 386932 123722 386948 123778
rect 308236 123706 386948 123722
rect 306780 123598 384932 123614
rect 306780 123542 306796 123598
rect 306852 123542 384860 123598
rect 384916 123542 384932 123598
rect 306780 123526 384932 123542
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 39954 118350
rect 40010 118294 40078 118350
rect 40134 118294 40202 118350
rect 40258 118294 40326 118350
rect 40382 118294 59878 118350
rect 59934 118294 60002 118350
rect 60058 118294 90598 118350
rect 90654 118294 90722 118350
rect 90778 118294 121318 118350
rect 121374 118294 121442 118350
rect 121498 118294 152038 118350
rect 152094 118294 152162 118350
rect 152218 118294 182758 118350
rect 182814 118294 182882 118350
rect 182938 118294 213478 118350
rect 213534 118294 213602 118350
rect 213658 118294 244198 118350
rect 244254 118294 244322 118350
rect 244378 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 479878 118350
rect 479934 118294 480002 118350
rect 480058 118294 510598 118350
rect 510654 118294 510722 118350
rect 510778 118294 541318 118350
rect 541374 118294 541442 118350
rect 541498 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 39954 118226
rect 40010 118170 40078 118226
rect 40134 118170 40202 118226
rect 40258 118170 40326 118226
rect 40382 118170 59878 118226
rect 59934 118170 60002 118226
rect 60058 118170 90598 118226
rect 90654 118170 90722 118226
rect 90778 118170 121318 118226
rect 121374 118170 121442 118226
rect 121498 118170 152038 118226
rect 152094 118170 152162 118226
rect 152218 118170 182758 118226
rect 182814 118170 182882 118226
rect 182938 118170 213478 118226
rect 213534 118170 213602 118226
rect 213658 118170 244198 118226
rect 244254 118170 244322 118226
rect 244378 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 479878 118226
rect 479934 118170 480002 118226
rect 480058 118170 510598 118226
rect 510654 118170 510722 118226
rect 510778 118170 541318 118226
rect 541374 118170 541442 118226
rect 541498 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 39954 118102
rect 40010 118046 40078 118102
rect 40134 118046 40202 118102
rect 40258 118046 40326 118102
rect 40382 118046 59878 118102
rect 59934 118046 60002 118102
rect 60058 118046 90598 118102
rect 90654 118046 90722 118102
rect 90778 118046 121318 118102
rect 121374 118046 121442 118102
rect 121498 118046 152038 118102
rect 152094 118046 152162 118102
rect 152218 118046 182758 118102
rect 182814 118046 182882 118102
rect 182938 118046 213478 118102
rect 213534 118046 213602 118102
rect 213658 118046 244198 118102
rect 244254 118046 244322 118102
rect 244378 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 479878 118102
rect 479934 118046 480002 118102
rect 480058 118046 510598 118102
rect 510654 118046 510722 118102
rect 510778 118046 541318 118102
rect 541374 118046 541442 118102
rect 541498 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 39954 117978
rect 40010 117922 40078 117978
rect 40134 117922 40202 117978
rect 40258 117922 40326 117978
rect 40382 117922 59878 117978
rect 59934 117922 60002 117978
rect 60058 117922 90598 117978
rect 90654 117922 90722 117978
rect 90778 117922 121318 117978
rect 121374 117922 121442 117978
rect 121498 117922 152038 117978
rect 152094 117922 152162 117978
rect 152218 117922 182758 117978
rect 182814 117922 182882 117978
rect 182938 117922 213478 117978
rect 213534 117922 213602 117978
rect 213658 117922 244198 117978
rect 244254 117922 244322 117978
rect 244378 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 479878 117978
rect 479934 117922 480002 117978
rect 480058 117922 510598 117978
rect 510654 117922 510722 117978
rect 510778 117922 541318 117978
rect 541374 117922 541442 117978
rect 541498 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect 359868 115858 457732 115874
rect 359868 115802 359884 115858
rect 359940 115802 457660 115858
rect 457716 115802 457732 115858
rect 359868 115786 457732 115802
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 44518 112350
rect 44574 112294 44642 112350
rect 44698 112294 75238 112350
rect 75294 112294 75362 112350
rect 75418 112294 105958 112350
rect 106014 112294 106082 112350
rect 106138 112294 136678 112350
rect 136734 112294 136802 112350
rect 136858 112294 167398 112350
rect 167454 112294 167522 112350
rect 167578 112294 198118 112350
rect 198174 112294 198242 112350
rect 198298 112294 228838 112350
rect 228894 112294 228962 112350
rect 229018 112294 259558 112350
rect 259614 112294 259682 112350
rect 259738 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 364518 112350
rect 364574 112294 364642 112350
rect 364698 112294 395238 112350
rect 395294 112294 395362 112350
rect 395418 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 464518 112350
rect 464574 112294 464642 112350
rect 464698 112294 495238 112350
rect 495294 112294 495362 112350
rect 495418 112294 525958 112350
rect 526014 112294 526082 112350
rect 526138 112294 556678 112350
rect 556734 112294 556802 112350
rect 556858 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 44518 112226
rect 44574 112170 44642 112226
rect 44698 112170 75238 112226
rect 75294 112170 75362 112226
rect 75418 112170 105958 112226
rect 106014 112170 106082 112226
rect 106138 112170 136678 112226
rect 136734 112170 136802 112226
rect 136858 112170 167398 112226
rect 167454 112170 167522 112226
rect 167578 112170 198118 112226
rect 198174 112170 198242 112226
rect 198298 112170 228838 112226
rect 228894 112170 228962 112226
rect 229018 112170 259558 112226
rect 259614 112170 259682 112226
rect 259738 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 364518 112226
rect 364574 112170 364642 112226
rect 364698 112170 395238 112226
rect 395294 112170 395362 112226
rect 395418 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 464518 112226
rect 464574 112170 464642 112226
rect 464698 112170 495238 112226
rect 495294 112170 495362 112226
rect 495418 112170 525958 112226
rect 526014 112170 526082 112226
rect 526138 112170 556678 112226
rect 556734 112170 556802 112226
rect 556858 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 44518 112102
rect 44574 112046 44642 112102
rect 44698 112046 75238 112102
rect 75294 112046 75362 112102
rect 75418 112046 105958 112102
rect 106014 112046 106082 112102
rect 106138 112046 136678 112102
rect 136734 112046 136802 112102
rect 136858 112046 167398 112102
rect 167454 112046 167522 112102
rect 167578 112046 198118 112102
rect 198174 112046 198242 112102
rect 198298 112046 228838 112102
rect 228894 112046 228962 112102
rect 229018 112046 259558 112102
rect 259614 112046 259682 112102
rect 259738 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 364518 112102
rect 364574 112046 364642 112102
rect 364698 112046 395238 112102
rect 395294 112046 395362 112102
rect 395418 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 464518 112102
rect 464574 112046 464642 112102
rect 464698 112046 495238 112102
rect 495294 112046 495362 112102
rect 495418 112046 525958 112102
rect 526014 112046 526082 112102
rect 526138 112046 556678 112102
rect 556734 112046 556802 112102
rect 556858 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 44518 111978
rect 44574 111922 44642 111978
rect 44698 111922 75238 111978
rect 75294 111922 75362 111978
rect 75418 111922 105958 111978
rect 106014 111922 106082 111978
rect 106138 111922 136678 111978
rect 136734 111922 136802 111978
rect 136858 111922 167398 111978
rect 167454 111922 167522 111978
rect 167578 111922 198118 111978
rect 198174 111922 198242 111978
rect 198298 111922 228838 111978
rect 228894 111922 228962 111978
rect 229018 111922 259558 111978
rect 259614 111922 259682 111978
rect 259738 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 364518 111978
rect 364574 111922 364642 111978
rect 364698 111922 395238 111978
rect 395294 111922 395362 111978
rect 395418 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 464518 111978
rect 464574 111922 464642 111978
rect 464698 111922 495238 111978
rect 495294 111922 495362 111978
rect 495418 111922 525958 111978
rect 526014 111922 526082 111978
rect 526138 111922 556678 111978
rect 556734 111922 556802 111978
rect 556858 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 59878 100350
rect 59934 100294 60002 100350
rect 60058 100294 90598 100350
rect 90654 100294 90722 100350
rect 90778 100294 121318 100350
rect 121374 100294 121442 100350
rect 121498 100294 152038 100350
rect 152094 100294 152162 100350
rect 152218 100294 182758 100350
rect 182814 100294 182882 100350
rect 182938 100294 213478 100350
rect 213534 100294 213602 100350
rect 213658 100294 244198 100350
rect 244254 100294 244322 100350
rect 244378 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 379878 100350
rect 379934 100294 380002 100350
rect 380058 100294 410598 100350
rect 410654 100294 410722 100350
rect 410778 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 479878 100350
rect 479934 100294 480002 100350
rect 480058 100294 510598 100350
rect 510654 100294 510722 100350
rect 510778 100294 541318 100350
rect 541374 100294 541442 100350
rect 541498 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 59878 100226
rect 59934 100170 60002 100226
rect 60058 100170 90598 100226
rect 90654 100170 90722 100226
rect 90778 100170 121318 100226
rect 121374 100170 121442 100226
rect 121498 100170 152038 100226
rect 152094 100170 152162 100226
rect 152218 100170 182758 100226
rect 182814 100170 182882 100226
rect 182938 100170 213478 100226
rect 213534 100170 213602 100226
rect 213658 100170 244198 100226
rect 244254 100170 244322 100226
rect 244378 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 379878 100226
rect 379934 100170 380002 100226
rect 380058 100170 410598 100226
rect 410654 100170 410722 100226
rect 410778 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 479878 100226
rect 479934 100170 480002 100226
rect 480058 100170 510598 100226
rect 510654 100170 510722 100226
rect 510778 100170 541318 100226
rect 541374 100170 541442 100226
rect 541498 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 59878 100102
rect 59934 100046 60002 100102
rect 60058 100046 90598 100102
rect 90654 100046 90722 100102
rect 90778 100046 121318 100102
rect 121374 100046 121442 100102
rect 121498 100046 152038 100102
rect 152094 100046 152162 100102
rect 152218 100046 182758 100102
rect 182814 100046 182882 100102
rect 182938 100046 213478 100102
rect 213534 100046 213602 100102
rect 213658 100046 244198 100102
rect 244254 100046 244322 100102
rect 244378 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 379878 100102
rect 379934 100046 380002 100102
rect 380058 100046 410598 100102
rect 410654 100046 410722 100102
rect 410778 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 479878 100102
rect 479934 100046 480002 100102
rect 480058 100046 510598 100102
rect 510654 100046 510722 100102
rect 510778 100046 541318 100102
rect 541374 100046 541442 100102
rect 541498 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 59878 99978
rect 59934 99922 60002 99978
rect 60058 99922 90598 99978
rect 90654 99922 90722 99978
rect 90778 99922 121318 99978
rect 121374 99922 121442 99978
rect 121498 99922 152038 99978
rect 152094 99922 152162 99978
rect 152218 99922 182758 99978
rect 182814 99922 182882 99978
rect 182938 99922 213478 99978
rect 213534 99922 213602 99978
rect 213658 99922 244198 99978
rect 244254 99922 244322 99978
rect 244378 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 379878 99978
rect 379934 99922 380002 99978
rect 380058 99922 410598 99978
rect 410654 99922 410722 99978
rect 410778 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 479878 99978
rect 479934 99922 480002 99978
rect 480058 99922 510598 99978
rect 510654 99922 510722 99978
rect 510778 99922 541318 99978
rect 541374 99922 541442 99978
rect 541498 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 44518 94350
rect 44574 94294 44642 94350
rect 44698 94294 75238 94350
rect 75294 94294 75362 94350
rect 75418 94294 105958 94350
rect 106014 94294 106082 94350
rect 106138 94294 136678 94350
rect 136734 94294 136802 94350
rect 136858 94294 167398 94350
rect 167454 94294 167522 94350
rect 167578 94294 198118 94350
rect 198174 94294 198242 94350
rect 198298 94294 228838 94350
rect 228894 94294 228962 94350
rect 229018 94294 259558 94350
rect 259614 94294 259682 94350
rect 259738 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 364518 94350
rect 364574 94294 364642 94350
rect 364698 94294 395238 94350
rect 395294 94294 395362 94350
rect 395418 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 464518 94350
rect 464574 94294 464642 94350
rect 464698 94294 495238 94350
rect 495294 94294 495362 94350
rect 495418 94294 525958 94350
rect 526014 94294 526082 94350
rect 526138 94294 556678 94350
rect 556734 94294 556802 94350
rect 556858 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 44518 94226
rect 44574 94170 44642 94226
rect 44698 94170 75238 94226
rect 75294 94170 75362 94226
rect 75418 94170 105958 94226
rect 106014 94170 106082 94226
rect 106138 94170 136678 94226
rect 136734 94170 136802 94226
rect 136858 94170 167398 94226
rect 167454 94170 167522 94226
rect 167578 94170 198118 94226
rect 198174 94170 198242 94226
rect 198298 94170 228838 94226
rect 228894 94170 228962 94226
rect 229018 94170 259558 94226
rect 259614 94170 259682 94226
rect 259738 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 364518 94226
rect 364574 94170 364642 94226
rect 364698 94170 395238 94226
rect 395294 94170 395362 94226
rect 395418 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 464518 94226
rect 464574 94170 464642 94226
rect 464698 94170 495238 94226
rect 495294 94170 495362 94226
rect 495418 94170 525958 94226
rect 526014 94170 526082 94226
rect 526138 94170 556678 94226
rect 556734 94170 556802 94226
rect 556858 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 44518 94102
rect 44574 94046 44642 94102
rect 44698 94046 75238 94102
rect 75294 94046 75362 94102
rect 75418 94046 105958 94102
rect 106014 94046 106082 94102
rect 106138 94046 136678 94102
rect 136734 94046 136802 94102
rect 136858 94046 167398 94102
rect 167454 94046 167522 94102
rect 167578 94046 198118 94102
rect 198174 94046 198242 94102
rect 198298 94046 228838 94102
rect 228894 94046 228962 94102
rect 229018 94046 259558 94102
rect 259614 94046 259682 94102
rect 259738 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 364518 94102
rect 364574 94046 364642 94102
rect 364698 94046 395238 94102
rect 395294 94046 395362 94102
rect 395418 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 464518 94102
rect 464574 94046 464642 94102
rect 464698 94046 495238 94102
rect 495294 94046 495362 94102
rect 495418 94046 525958 94102
rect 526014 94046 526082 94102
rect 526138 94046 556678 94102
rect 556734 94046 556802 94102
rect 556858 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 44518 93978
rect 44574 93922 44642 93978
rect 44698 93922 75238 93978
rect 75294 93922 75362 93978
rect 75418 93922 105958 93978
rect 106014 93922 106082 93978
rect 106138 93922 136678 93978
rect 136734 93922 136802 93978
rect 136858 93922 167398 93978
rect 167454 93922 167522 93978
rect 167578 93922 198118 93978
rect 198174 93922 198242 93978
rect 198298 93922 228838 93978
rect 228894 93922 228962 93978
rect 229018 93922 259558 93978
rect 259614 93922 259682 93978
rect 259738 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 364518 93978
rect 364574 93922 364642 93978
rect 364698 93922 395238 93978
rect 395294 93922 395362 93978
rect 395418 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 464518 93978
rect 464574 93922 464642 93978
rect 464698 93922 495238 93978
rect 495294 93922 495362 93978
rect 495418 93922 525958 93978
rect 526014 93922 526082 93978
rect 526138 93922 556678 93978
rect 556734 93922 556802 93978
rect 556858 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 59878 82350
rect 59934 82294 60002 82350
rect 60058 82294 90598 82350
rect 90654 82294 90722 82350
rect 90778 82294 121318 82350
rect 121374 82294 121442 82350
rect 121498 82294 152038 82350
rect 152094 82294 152162 82350
rect 152218 82294 182758 82350
rect 182814 82294 182882 82350
rect 182938 82294 213478 82350
rect 213534 82294 213602 82350
rect 213658 82294 244198 82350
rect 244254 82294 244322 82350
rect 244378 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 379878 82350
rect 379934 82294 380002 82350
rect 380058 82294 410598 82350
rect 410654 82294 410722 82350
rect 410778 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 479878 82350
rect 479934 82294 480002 82350
rect 480058 82294 510598 82350
rect 510654 82294 510722 82350
rect 510778 82294 541318 82350
rect 541374 82294 541442 82350
rect 541498 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 59878 82226
rect 59934 82170 60002 82226
rect 60058 82170 90598 82226
rect 90654 82170 90722 82226
rect 90778 82170 121318 82226
rect 121374 82170 121442 82226
rect 121498 82170 152038 82226
rect 152094 82170 152162 82226
rect 152218 82170 182758 82226
rect 182814 82170 182882 82226
rect 182938 82170 213478 82226
rect 213534 82170 213602 82226
rect 213658 82170 244198 82226
rect 244254 82170 244322 82226
rect 244378 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 379878 82226
rect 379934 82170 380002 82226
rect 380058 82170 410598 82226
rect 410654 82170 410722 82226
rect 410778 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 479878 82226
rect 479934 82170 480002 82226
rect 480058 82170 510598 82226
rect 510654 82170 510722 82226
rect 510778 82170 541318 82226
rect 541374 82170 541442 82226
rect 541498 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82147 597980 82170
rect -1916 82102 299528 82147
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 59878 82102
rect 59934 82046 60002 82102
rect 60058 82046 90598 82102
rect 90654 82046 90722 82102
rect 90778 82046 121318 82102
rect 121374 82046 121442 82102
rect 121498 82046 152038 82102
rect 152094 82046 152162 82102
rect 152218 82046 182758 82102
rect 182814 82046 182882 82102
rect 182938 82046 213478 82102
rect 213534 82046 213602 82102
rect 213658 82046 244198 82102
rect 244254 82046 244322 82102
rect 244378 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82091 299528 82102
rect 299584 82091 299632 82147
rect 299688 82091 299736 82147
rect 299792 82091 307844 82147
rect 307900 82091 307948 82147
rect 308004 82091 308052 82147
rect 308108 82091 316160 82147
rect 316216 82091 316264 82147
rect 316320 82091 316368 82147
rect 316424 82091 324476 82147
rect 324532 82091 324580 82147
rect 324636 82091 324684 82147
rect 324740 82102 597980 82147
rect 324740 82091 347154 82102
rect 286142 82046 347154 82091
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 379878 82102
rect 379934 82046 380002 82102
rect 380058 82046 410598 82102
rect 410654 82046 410722 82102
rect 410778 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 479878 82102
rect 479934 82046 480002 82102
rect 480058 82046 510598 82102
rect 510654 82046 510722 82102
rect 510778 82046 541318 82102
rect 541374 82046 541442 82102
rect 541498 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 82043 597980 82046
rect -1916 81987 299528 82043
rect 299584 81987 299632 82043
rect 299688 81987 299736 82043
rect 299792 81987 307844 82043
rect 307900 81987 307948 82043
rect 308004 81987 308052 82043
rect 308108 81987 316160 82043
rect 316216 81987 316264 82043
rect 316320 81987 316368 82043
rect 316424 81987 324476 82043
rect 324532 81987 324580 82043
rect 324636 81987 324684 82043
rect 324740 81987 597980 82043
rect -1916 81978 597980 81987
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 59878 81978
rect 59934 81922 60002 81978
rect 60058 81922 90598 81978
rect 90654 81922 90722 81978
rect 90778 81922 121318 81978
rect 121374 81922 121442 81978
rect 121498 81922 152038 81978
rect 152094 81922 152162 81978
rect 152218 81922 182758 81978
rect 182814 81922 182882 81978
rect 182938 81922 213478 81978
rect 213534 81922 213602 81978
rect 213658 81922 244198 81978
rect 244254 81922 244322 81978
rect 244378 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81939 347154 81978
rect 286142 81922 299528 81939
rect -1916 81883 299528 81922
rect 299584 81883 299632 81939
rect 299688 81883 299736 81939
rect 299792 81883 307844 81939
rect 307900 81883 307948 81939
rect 308004 81883 308052 81939
rect 308108 81883 316160 81939
rect 316216 81883 316264 81939
rect 316320 81883 316368 81939
rect 316424 81883 324476 81939
rect 324532 81883 324580 81939
rect 324636 81883 324684 81939
rect 324740 81922 347154 81939
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 379878 81978
rect 379934 81922 380002 81978
rect 380058 81922 410598 81978
rect 410654 81922 410722 81978
rect 410778 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 479878 81978
rect 479934 81922 480002 81978
rect 480058 81922 510598 81978
rect 510654 81922 510722 81978
rect 510778 81922 541318 81978
rect 541374 81922 541442 81978
rect 541498 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 324740 81883 597980 81922
rect -1916 81826 597980 81883
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 44518 76350
rect 44574 76294 44642 76350
rect 44698 76294 75238 76350
rect 75294 76294 75362 76350
rect 75418 76294 105958 76350
rect 106014 76294 106082 76350
rect 106138 76294 136678 76350
rect 136734 76294 136802 76350
rect 136858 76294 167398 76350
rect 167454 76294 167522 76350
rect 167578 76294 198118 76350
rect 198174 76294 198242 76350
rect 198298 76294 228838 76350
rect 228894 76294 228962 76350
rect 229018 76294 259558 76350
rect 259614 76294 259682 76350
rect 259738 76294 281994 76350
rect 282050 76294 282118 76350
rect 282174 76294 282242 76350
rect 282298 76294 282366 76350
rect 282422 76294 295412 76350
rect 295468 76294 295536 76350
rect 295592 76294 303728 76350
rect 303784 76294 303852 76350
rect 303908 76294 312044 76350
rect 312100 76294 312168 76350
rect 312224 76294 312714 76350
rect 312770 76294 312838 76350
rect 312894 76294 312962 76350
rect 313018 76294 313086 76350
rect 313142 76294 320360 76350
rect 320416 76294 320484 76350
rect 320540 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 364518 76350
rect 364574 76294 364642 76350
rect 364698 76294 395238 76350
rect 395294 76294 395362 76350
rect 395418 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 464518 76350
rect 464574 76294 464642 76350
rect 464698 76294 495238 76350
rect 495294 76294 495362 76350
rect 495418 76294 525958 76350
rect 526014 76294 526082 76350
rect 526138 76294 556678 76350
rect 556734 76294 556802 76350
rect 556858 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 44518 76226
rect 44574 76170 44642 76226
rect 44698 76170 75238 76226
rect 75294 76170 75362 76226
rect 75418 76170 105958 76226
rect 106014 76170 106082 76226
rect 106138 76170 136678 76226
rect 136734 76170 136802 76226
rect 136858 76170 167398 76226
rect 167454 76170 167522 76226
rect 167578 76170 198118 76226
rect 198174 76170 198242 76226
rect 198298 76170 228838 76226
rect 228894 76170 228962 76226
rect 229018 76170 259558 76226
rect 259614 76170 259682 76226
rect 259738 76170 281994 76226
rect 282050 76170 282118 76226
rect 282174 76170 282242 76226
rect 282298 76170 282366 76226
rect 282422 76170 295412 76226
rect 295468 76170 295536 76226
rect 295592 76170 303728 76226
rect 303784 76170 303852 76226
rect 303908 76170 312044 76226
rect 312100 76170 312168 76226
rect 312224 76170 312714 76226
rect 312770 76170 312838 76226
rect 312894 76170 312962 76226
rect 313018 76170 313086 76226
rect 313142 76170 320360 76226
rect 320416 76170 320484 76226
rect 320540 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 364518 76226
rect 364574 76170 364642 76226
rect 364698 76170 395238 76226
rect 395294 76170 395362 76226
rect 395418 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 464518 76226
rect 464574 76170 464642 76226
rect 464698 76170 495238 76226
rect 495294 76170 495362 76226
rect 495418 76170 525958 76226
rect 526014 76170 526082 76226
rect 526138 76170 556678 76226
rect 556734 76170 556802 76226
rect 556858 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 44518 76102
rect 44574 76046 44642 76102
rect 44698 76046 75238 76102
rect 75294 76046 75362 76102
rect 75418 76046 105958 76102
rect 106014 76046 106082 76102
rect 106138 76046 136678 76102
rect 136734 76046 136802 76102
rect 136858 76046 167398 76102
rect 167454 76046 167522 76102
rect 167578 76046 198118 76102
rect 198174 76046 198242 76102
rect 198298 76046 228838 76102
rect 228894 76046 228962 76102
rect 229018 76046 259558 76102
rect 259614 76046 259682 76102
rect 259738 76046 281994 76102
rect 282050 76046 282118 76102
rect 282174 76046 282242 76102
rect 282298 76046 282366 76102
rect 282422 76046 295412 76102
rect 295468 76046 295536 76102
rect 295592 76046 303728 76102
rect 303784 76046 303852 76102
rect 303908 76046 312044 76102
rect 312100 76046 312168 76102
rect 312224 76046 312714 76102
rect 312770 76046 312838 76102
rect 312894 76046 312962 76102
rect 313018 76046 313086 76102
rect 313142 76046 320360 76102
rect 320416 76046 320484 76102
rect 320540 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 364518 76102
rect 364574 76046 364642 76102
rect 364698 76046 395238 76102
rect 395294 76046 395362 76102
rect 395418 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 464518 76102
rect 464574 76046 464642 76102
rect 464698 76046 495238 76102
rect 495294 76046 495362 76102
rect 495418 76046 525958 76102
rect 526014 76046 526082 76102
rect 526138 76046 556678 76102
rect 556734 76046 556802 76102
rect 556858 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 44518 75978
rect 44574 75922 44642 75978
rect 44698 75922 75238 75978
rect 75294 75922 75362 75978
rect 75418 75922 105958 75978
rect 106014 75922 106082 75978
rect 106138 75922 136678 75978
rect 136734 75922 136802 75978
rect 136858 75922 167398 75978
rect 167454 75922 167522 75978
rect 167578 75922 198118 75978
rect 198174 75922 198242 75978
rect 198298 75922 228838 75978
rect 228894 75922 228962 75978
rect 229018 75922 259558 75978
rect 259614 75922 259682 75978
rect 259738 75922 281994 75978
rect 282050 75922 282118 75978
rect 282174 75922 282242 75978
rect 282298 75922 282366 75978
rect 282422 75922 295412 75978
rect 295468 75922 295536 75978
rect 295592 75922 303728 75978
rect 303784 75922 303852 75978
rect 303908 75922 312044 75978
rect 312100 75922 312168 75978
rect 312224 75922 312714 75978
rect 312770 75922 312838 75978
rect 312894 75922 312962 75978
rect 313018 75922 313086 75978
rect 313142 75922 320360 75978
rect 320416 75922 320484 75978
rect 320540 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 364518 75978
rect 364574 75922 364642 75978
rect 364698 75922 395238 75978
rect 395294 75922 395362 75978
rect 395418 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 464518 75978
rect 464574 75922 464642 75978
rect 464698 75922 495238 75978
rect 495294 75922 495362 75978
rect 495418 75922 525958 75978
rect 526014 75922 526082 75978
rect 526138 75922 556678 75978
rect 556734 75922 556802 75978
rect 556858 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 39954 64350
rect 40010 64294 40078 64350
rect 40134 64294 40202 64350
rect 40258 64294 40326 64350
rect 40382 64294 59878 64350
rect 59934 64294 60002 64350
rect 60058 64294 90598 64350
rect 90654 64294 90722 64350
rect 90778 64294 121318 64350
rect 121374 64294 121442 64350
rect 121498 64294 152038 64350
rect 152094 64294 152162 64350
rect 152218 64294 182758 64350
rect 182814 64294 182882 64350
rect 182938 64294 213478 64350
rect 213534 64294 213602 64350
rect 213658 64294 244198 64350
rect 244254 64294 244322 64350
rect 244378 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 299570 64350
rect 299626 64294 299694 64350
rect 299750 64294 307886 64350
rect 307942 64294 308010 64350
rect 308066 64294 316202 64350
rect 316258 64294 316326 64350
rect 316382 64294 324518 64350
rect 324574 64294 324642 64350
rect 324698 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 379878 64350
rect 379934 64294 380002 64350
rect 380058 64294 410598 64350
rect 410654 64294 410722 64350
rect 410778 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 479878 64350
rect 479934 64294 480002 64350
rect 480058 64294 510598 64350
rect 510654 64294 510722 64350
rect 510778 64294 541318 64350
rect 541374 64294 541442 64350
rect 541498 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 39954 64226
rect 40010 64170 40078 64226
rect 40134 64170 40202 64226
rect 40258 64170 40326 64226
rect 40382 64170 59878 64226
rect 59934 64170 60002 64226
rect 60058 64170 90598 64226
rect 90654 64170 90722 64226
rect 90778 64170 121318 64226
rect 121374 64170 121442 64226
rect 121498 64170 152038 64226
rect 152094 64170 152162 64226
rect 152218 64170 182758 64226
rect 182814 64170 182882 64226
rect 182938 64170 213478 64226
rect 213534 64170 213602 64226
rect 213658 64170 244198 64226
rect 244254 64170 244322 64226
rect 244378 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 299570 64226
rect 299626 64170 299694 64226
rect 299750 64170 307886 64226
rect 307942 64170 308010 64226
rect 308066 64170 316202 64226
rect 316258 64170 316326 64226
rect 316382 64170 324518 64226
rect 324574 64170 324642 64226
rect 324698 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 379878 64226
rect 379934 64170 380002 64226
rect 380058 64170 410598 64226
rect 410654 64170 410722 64226
rect 410778 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 479878 64226
rect 479934 64170 480002 64226
rect 480058 64170 510598 64226
rect 510654 64170 510722 64226
rect 510778 64170 541318 64226
rect 541374 64170 541442 64226
rect 541498 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 39954 64102
rect 40010 64046 40078 64102
rect 40134 64046 40202 64102
rect 40258 64046 40326 64102
rect 40382 64046 59878 64102
rect 59934 64046 60002 64102
rect 60058 64046 90598 64102
rect 90654 64046 90722 64102
rect 90778 64046 121318 64102
rect 121374 64046 121442 64102
rect 121498 64046 152038 64102
rect 152094 64046 152162 64102
rect 152218 64046 182758 64102
rect 182814 64046 182882 64102
rect 182938 64046 213478 64102
rect 213534 64046 213602 64102
rect 213658 64046 244198 64102
rect 244254 64046 244322 64102
rect 244378 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 299570 64102
rect 299626 64046 299694 64102
rect 299750 64046 307886 64102
rect 307942 64046 308010 64102
rect 308066 64046 316202 64102
rect 316258 64046 316326 64102
rect 316382 64046 324518 64102
rect 324574 64046 324642 64102
rect 324698 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 379878 64102
rect 379934 64046 380002 64102
rect 380058 64046 410598 64102
rect 410654 64046 410722 64102
rect 410778 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 479878 64102
rect 479934 64046 480002 64102
rect 480058 64046 510598 64102
rect 510654 64046 510722 64102
rect 510778 64046 541318 64102
rect 541374 64046 541442 64102
rect 541498 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 39954 63978
rect 40010 63922 40078 63978
rect 40134 63922 40202 63978
rect 40258 63922 40326 63978
rect 40382 63922 59878 63978
rect 59934 63922 60002 63978
rect 60058 63922 90598 63978
rect 90654 63922 90722 63978
rect 90778 63922 121318 63978
rect 121374 63922 121442 63978
rect 121498 63922 152038 63978
rect 152094 63922 152162 63978
rect 152218 63922 182758 63978
rect 182814 63922 182882 63978
rect 182938 63922 213478 63978
rect 213534 63922 213602 63978
rect 213658 63922 244198 63978
rect 244254 63922 244322 63978
rect 244378 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 299570 63978
rect 299626 63922 299694 63978
rect 299750 63922 307886 63978
rect 307942 63922 308010 63978
rect 308066 63922 316202 63978
rect 316258 63922 316326 63978
rect 316382 63922 324518 63978
rect 324574 63922 324642 63978
rect 324698 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 379878 63978
rect 379934 63922 380002 63978
rect 380058 63922 410598 63978
rect 410654 63922 410722 63978
rect 410778 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 479878 63978
rect 479934 63922 480002 63978
rect 480058 63922 510598 63978
rect 510654 63922 510722 63978
rect 510778 63922 541318 63978
rect 541374 63922 541442 63978
rect 541498 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 44518 58350
rect 44574 58294 44642 58350
rect 44698 58294 75238 58350
rect 75294 58294 75362 58350
rect 75418 58294 105958 58350
rect 106014 58294 106082 58350
rect 106138 58294 136678 58350
rect 136734 58294 136802 58350
rect 136858 58294 167398 58350
rect 167454 58294 167522 58350
rect 167578 58294 198118 58350
rect 198174 58294 198242 58350
rect 198298 58294 228838 58350
rect 228894 58294 228962 58350
rect 229018 58294 259558 58350
rect 259614 58294 259682 58350
rect 259738 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 295412 58350
rect 295468 58294 295536 58350
rect 295592 58294 303728 58350
rect 303784 58294 303852 58350
rect 303908 58294 312044 58350
rect 312100 58294 312168 58350
rect 312224 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 320360 58350
rect 320416 58294 320484 58350
rect 320540 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 364518 58350
rect 364574 58294 364642 58350
rect 364698 58294 395238 58350
rect 395294 58294 395362 58350
rect 395418 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 464518 58350
rect 464574 58294 464642 58350
rect 464698 58294 495238 58350
rect 495294 58294 495362 58350
rect 495418 58294 525958 58350
rect 526014 58294 526082 58350
rect 526138 58294 556678 58350
rect 556734 58294 556802 58350
rect 556858 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 44518 58226
rect 44574 58170 44642 58226
rect 44698 58170 75238 58226
rect 75294 58170 75362 58226
rect 75418 58170 105958 58226
rect 106014 58170 106082 58226
rect 106138 58170 136678 58226
rect 136734 58170 136802 58226
rect 136858 58170 167398 58226
rect 167454 58170 167522 58226
rect 167578 58170 198118 58226
rect 198174 58170 198242 58226
rect 198298 58170 228838 58226
rect 228894 58170 228962 58226
rect 229018 58170 259558 58226
rect 259614 58170 259682 58226
rect 259738 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 295412 58226
rect 295468 58170 295536 58226
rect 295592 58170 303728 58226
rect 303784 58170 303852 58226
rect 303908 58170 312044 58226
rect 312100 58170 312168 58226
rect 312224 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 320360 58226
rect 320416 58170 320484 58226
rect 320540 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 364518 58226
rect 364574 58170 364642 58226
rect 364698 58170 395238 58226
rect 395294 58170 395362 58226
rect 395418 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 464518 58226
rect 464574 58170 464642 58226
rect 464698 58170 495238 58226
rect 495294 58170 495362 58226
rect 495418 58170 525958 58226
rect 526014 58170 526082 58226
rect 526138 58170 556678 58226
rect 556734 58170 556802 58226
rect 556858 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 44518 58102
rect 44574 58046 44642 58102
rect 44698 58046 75238 58102
rect 75294 58046 75362 58102
rect 75418 58046 105958 58102
rect 106014 58046 106082 58102
rect 106138 58046 136678 58102
rect 136734 58046 136802 58102
rect 136858 58046 167398 58102
rect 167454 58046 167522 58102
rect 167578 58046 198118 58102
rect 198174 58046 198242 58102
rect 198298 58046 228838 58102
rect 228894 58046 228962 58102
rect 229018 58046 259558 58102
rect 259614 58046 259682 58102
rect 259738 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 295412 58102
rect 295468 58046 295536 58102
rect 295592 58046 303728 58102
rect 303784 58046 303852 58102
rect 303908 58046 312044 58102
rect 312100 58046 312168 58102
rect 312224 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 320360 58102
rect 320416 58046 320484 58102
rect 320540 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 364518 58102
rect 364574 58046 364642 58102
rect 364698 58046 395238 58102
rect 395294 58046 395362 58102
rect 395418 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 464518 58102
rect 464574 58046 464642 58102
rect 464698 58046 495238 58102
rect 495294 58046 495362 58102
rect 495418 58046 525958 58102
rect 526014 58046 526082 58102
rect 526138 58046 556678 58102
rect 556734 58046 556802 58102
rect 556858 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 44518 57978
rect 44574 57922 44642 57978
rect 44698 57922 75238 57978
rect 75294 57922 75362 57978
rect 75418 57922 105958 57978
rect 106014 57922 106082 57978
rect 106138 57922 136678 57978
rect 136734 57922 136802 57978
rect 136858 57922 167398 57978
rect 167454 57922 167522 57978
rect 167578 57922 198118 57978
rect 198174 57922 198242 57978
rect 198298 57922 228838 57978
rect 228894 57922 228962 57978
rect 229018 57922 259558 57978
rect 259614 57922 259682 57978
rect 259738 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 295412 57978
rect 295468 57922 295536 57978
rect 295592 57922 303728 57978
rect 303784 57922 303852 57978
rect 303908 57922 312044 57978
rect 312100 57922 312168 57978
rect 312224 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 320360 57978
rect 320416 57922 320484 57978
rect 320540 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 364518 57978
rect 364574 57922 364642 57978
rect 364698 57922 395238 57978
rect 395294 57922 395362 57978
rect 395418 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 464518 57978
rect 464574 57922 464642 57978
rect 464698 57922 495238 57978
rect 495294 57922 495362 57978
rect 495418 57922 525958 57978
rect 526014 57922 526082 57978
rect 526138 57922 556678 57978
rect 556734 57922 556802 57978
rect 556858 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect 209116 47998 312468 48014
rect 209116 47942 209132 47998
rect 209188 47942 312396 47998
rect 312452 47942 312468 47998
rect 209116 47926 312468 47942
rect 172940 47818 311796 47834
rect 172940 47762 172956 47818
rect 173012 47762 311724 47818
rect 311780 47762 311796 47818
rect 172940 47746 311796 47762
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 39954 46350
rect 40010 46294 40078 46350
rect 40134 46294 40202 46350
rect 40258 46294 40326 46350
rect 40382 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 101394 46350
rect 101450 46294 101518 46350
rect 101574 46294 101642 46350
rect 101698 46294 101766 46350
rect 101822 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 39954 46226
rect 40010 46170 40078 46226
rect 40134 46170 40202 46226
rect 40258 46170 40326 46226
rect 40382 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 101394 46226
rect 101450 46170 101518 46226
rect 101574 46170 101642 46226
rect 101698 46170 101766 46226
rect 101822 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 39954 46102
rect 40010 46046 40078 46102
rect 40134 46046 40202 46102
rect 40258 46046 40326 46102
rect 40382 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 101394 46102
rect 101450 46046 101518 46102
rect 101574 46046 101642 46102
rect 101698 46046 101766 46102
rect 101822 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 39954 45978
rect 40010 45922 40078 45978
rect 40134 45922 40202 45978
rect 40258 45922 40326 45978
rect 40382 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 101394 45978
rect 101450 45922 101518 45978
rect 101574 45922 101642 45978
rect 101698 45922 101766 45978
rect 101822 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect 39660 4978 60916 4994
rect 39660 4922 39676 4978
rect 39732 4922 60844 4978
rect 60900 4922 60916 4978
rect 39660 4906 60916 4922
rect 91516 4978 315044 4994
rect 91516 4922 91532 4978
rect 91588 4922 314972 4978
rect 315028 4922 315044 4978
rect 91516 4906 315044 4922
rect 34956 4798 55204 4814
rect 34956 4742 34972 4798
rect 35028 4742 55132 4798
rect 55188 4742 55204 4798
rect 34956 4726 55204 4742
rect 142924 4798 284804 4814
rect 142924 4742 142940 4798
rect 142996 4742 284732 4798
rect 284788 4742 284804 4798
rect 142924 4726 284804 4742
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use avali_logo  avali_logo
timestamp 0
transform 1 0 60000 0 1 475000
box 0 0 80000 93920
use wrapped_ay8913  ay8913
timestamp 0
transform 1 0 40000 0 1 240000
box 1258 0 60000 60000
use blinker  blinker
timestamp 0
transform 1 0 290000 0 1 50000
box 1258 0 34768 32230
use hellorld  hellorld
timestamp 0
transform 1 0 140000 0 1 260000
box 1258 1792 26000 26000
use wrapped_mc14500  mc14500
timestamp 0
transform 1 0 310000 0 1 160000
box 1258 0 37000 37000
use multiplexer  multiplexer
timestamp 0
transform 1 0 190000 0 1 240000
box 0 0 150000 140000
use wrapped_sid  sid
timestamp 0
transform 1 0 40000 0 1 50000
box 1258 0 230000 160000
use tholin_avalonsemi_tbb1143  tbb1143
timestamp 0
transform 1 0 130000 0 1 320000
box 1258 2688 46000 43120
use wrapped_pdp11  wrapped_pdp11
timestamp 0
transform 1 0 190000 0 1 410000
box 0 0 360000 156860
use wrapped_qcpu  wrapped_qcpu
timestamp 0
transform 1 0 460000 0 1 50000
box 0 802 100000 100000
use wrapped_sn76489  wrapped_sn76489
timestamp 0
transform 1 0 360000 0 1 50000
box 0 3076 60000 70000
use wrapped_tholin_riscv  wrapped_tholin_riscv
timestamp 0
transform 1 0 360000 0 1 175000
box 0 0 198782 220000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 210462 67478 245074 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 298094 67478 484408 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 530232 67478 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 210462 98198 473048 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 541432 98198 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 210462 128918 491128 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 539352 128918 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 210462 159638 260964 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 284908 159638 323954 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 364206 159638 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 210462 190358 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 210462 221078 241154 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 367758 221078 410034 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 568670 221078 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 48802 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 210462 251798 241154 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 367758 251798 410034 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 568670 251798 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 241154 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 367758 282518 410034 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 568670 282518 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 241154 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 367758 313238 410034 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 568670 313238 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 163170 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 193230 343958 410034 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 568670 343958 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 53730 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 115262 374678 173466 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 568670 374678 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 53730 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 115262 405398 173466 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 568670 405398 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 173466 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 568670 436118 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 48690 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 568670 466838 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 48690 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 568670 497558 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 48690 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 394038 528278 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 48690 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 394038 558998 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 -1644 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 -1644 40478 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 -1644 71198 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 210462 71198 245074 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 298094 71198 480728 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 533912 71198 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 -1644 101918 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 210462 101918 473528 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 542872 101918 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 -1644 132638 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 210462 132638 493368 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 542072 132638 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 -1644 163358 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 210462 163358 265522 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 282254 163358 323954 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 364206 163358 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 -1644 194078 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 210462 194078 410034 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 568670 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 -1644 224798 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 367758 224798 410034 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 568670 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 -1644 255518 48802 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 367758 255518 410034 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 568670 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 -1644 286238 241154 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 367758 286238 410034 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 568670 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 -1644 316958 50964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 84316 316958 163170 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 193230 316958 241154 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 367758 316958 410034 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 568670 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 -1644 347678 163170 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 193230 347678 410034 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 568670 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 -1644 378398 53730 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 115262 378398 173466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 568670 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 -1644 409118 53730 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 115262 409118 173466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 568670 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 -1644 439838 173466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 568670 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 -1644 470558 48690 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 149870 470558 173466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 568670 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 -1644 501278 48690 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 149870 501278 173466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 568670 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 -1644 531998 48690 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 149870 531998 173466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 394038 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 -1644 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 548990 382322 548990 382322 0 vdd
rlabel via4 533630 388322 533630 388322 0 vss
rlabel metal2 42210 240520 42210 240520 0 ay8913_do\[0\]
rlabel metal2 259098 379960 259098 379960 0 ay8913_do\[10\]
rlabel metal2 259994 379960 259994 379960 0 ay8913_do\[11\]
rlabel metal2 260890 379960 260890 379960 0 ay8913_do\[12\]
rlabel metal2 262206 379960 262206 379960 0 ay8913_do\[13\]
rlabel metal2 70952 237594 70952 237594 0 ay8913_do\[14\]
rlabel metal4 72968 238007 72968 238007 0 ay8913_do\[15\]
rlabel metal2 264474 379960 264474 379960 0 ay8913_do\[16\]
rlabel metal4 77000 238097 77000 238097 0 ay8913_do\[17\]
rlabel metal2 266266 379960 266266 379960 0 ay8913_do\[18\]
rlabel metal2 125160 310632 125160 310632 0 ay8913_do\[19\]
rlabel metal2 44450 240520 44450 240520 0 ay8913_do\[1\]
rlabel metal2 100408 311416 100408 311416 0 ay8913_do\[20\]
rlabel metal2 118440 310800 118440 310800 0 ay8913_do\[21\]
rlabel metal2 96600 237888 96600 237888 0 ay8913_do\[22\]
rlabel metal2 100184 311248 100184 311248 0 ay8913_do\[23\]
rlabel metal3 96824 238280 96824 238280 0 ay8913_do\[24\]
rlabel via3 97048 238255 97048 238255 0 ay8913_do\[25\]
rlabel metal2 95144 239274 95144 239274 0 ay8913_do\[26\]
rlabel metal2 97160 239218 97160 239218 0 ay8913_do\[27\]
rlabel metal2 46760 239274 46760 239274 0 ay8913_do\[2\]
rlabel metal2 48776 239106 48776 239106 0 ay8913_do\[3\]
rlabel metal2 50792 239162 50792 239162 0 ay8913_do\[4\]
rlabel metal2 52808 239218 52808 239218 0 ay8913_do\[5\]
rlabel metal2 54824 238994 54824 238994 0 ay8913_do\[6\]
rlabel metal2 256410 379960 256410 379960 0 ay8913_do\[7\]
rlabel metal2 257362 379960 257362 379960 0 ay8913_do\[8\]
rlabel metal2 258202 379960 258202 379960 0 ay8913_do\[9\]
rlabel metal2 233114 379960 233114 379960 0 blinker_do\[0\]
rlabel metal2 234766 379960 234766 379960 0 blinker_do\[1\]
rlabel metal4 235256 374065 235256 374065 0 blinker_do\[2\]
rlabel metal3 167006 261800 167006 261800 0 custom_settings\[0\]
rlabel metal4 359352 255777 359352 255777 0 custom_settings\[10\]
rlabel metal3 167566 283976 167566 283976 0 custom_settings\[11\]
rlabel metal3 188650 514920 188650 514920 0 custom_settings\[12\]
rlabel metal4 355544 204120 355544 204120 0 custom_settings\[13\]
rlabel metal3 188258 529256 188258 529256 0 custom_settings\[14\]
rlabel metal3 188930 536424 188930 536424 0 custom_settings\[15\]
rlabel metal3 188090 543592 188090 543592 0 custom_settings\[16\]
rlabel metal3 355376 280504 355376 280504 0 custom_settings\[17\]
rlabel metal3 188986 557928 188986 557928 0 custom_settings\[18\]
rlabel metal3 188202 565096 188202 565096 0 custom_settings\[19\]
rlabel metal3 167062 263816 167062 263816 0 custom_settings\[1\]
rlabel via4 457688 115847 457688 115847 0 custom_settings\[20\]
rlabel metal4 457688 120400 457688 120400 0 custom_settings\[21\]
rlabel metal3 459368 121772 459368 121772 0 custom_settings\[22\]
rlabel metal4 352632 160664 352632 160664 0 custom_settings\[23\]
rlabel metal3 344666 299656 344666 299656 0 custom_settings\[24\]
rlabel metal4 355768 216216 355768 216216 0 custom_settings\[25\]
rlabel metal4 352184 217448 352184 217448 0 custom_settings\[26\]
rlabel metal4 354200 219352 354200 219352 0 custom_settings\[27\]
rlabel metal4 356104 168168 356104 168168 0 custom_settings\[28\]
rlabel metal4 354312 223160 354312 223160 0 custom_settings\[29\]
rlabel metal3 187264 282184 187264 282184 0 custom_settings\[2\]
rlabel metal5 337204 304830 337204 304830 0 custom_settings\[30\]
rlabel metal4 352520 234192 352520 234192 0 custom_settings\[31\]
rlabel metal3 188818 450408 188818 450408 0 custom_settings\[3\]
rlabel metal3 168238 269864 168238 269864 0 custom_settings\[4\]
rlabel metal3 188874 464744 188874 464744 0 custom_settings\[5\]
rlabel metal3 186536 283864 186536 283864 0 custom_settings\[6\]
rlabel metal3 189224 285768 189224 285768 0 custom_settings\[7\]
rlabel metal4 188104 286207 188104 286207 0 custom_settings\[8\]
rlabel metal4 190736 234990 190736 234990 0 custom_settings\[9\]
rlabel metal2 161336 292894 161336 292894 0 hellorld_do
rlabel metal3 195832 379400 195832 379400 0 io_in[0]
rlabel metal3 358344 232344 358344 232344 0 io_in[10]
rlabel metal3 358232 238168 358232 238168 0 io_in[11]
rlabel metal3 351344 188104 351344 188104 0 io_in[12]
rlabel metal3 357336 406616 357336 406616 0 io_in[13]
rlabel metal4 243544 407785 243544 407785 0 io_in[14]
rlabel metal3 357280 164584 357280 164584 0 io_in[15]
rlabel metal3 357560 406728 357560 406728 0 io_in[16]
rlabel metal3 357672 235144 357672 235144 0 io_in[17]
rlabel metal3 265664 406616 265664 406616 0 io_in[18]
rlabel metal3 78176 304024 78176 304024 0 io_in[19]
rlabel metal3 93240 304024 93240 304024 0 io_in[20]
rlabel metal3 188216 487256 188216 487256 0 io_in[21]
rlabel metal2 121352 583002 121352 583002 0 io_in[22]
rlabel metal2 55160 502418 55160 502418 0 io_in[23]
rlabel metal3 358736 240296 358736 240296 0 io_in[24]
rlabel metal2 302974 410088 302974 410088 0 io_in[25]
rlabel metal4 312088 172169 312088 172169 0 io_in[26]
rlabel metal3 355992 331016 355992 331016 0 io_in[27]
rlabel metal3 359786 337232 359786 337232 0 io_in[28]
rlabel metal3 2310 375704 2310 375704 0 io_in[29]
rlabel metal3 2310 333368 2310 333368 0 io_in[30]
rlabel metal4 307384 145751 307384 145751 0 io_in[31]
rlabel metal3 359464 360500 359464 360500 0 io_in[32]
rlabel metal3 2310 206360 2310 206360 0 io_in[33]
rlabel metal3 2310 164024 2310 164024 0 io_in[34]
rlabel metal3 2310 121688 2310 121688 0 io_in[35]
rlabel metal3 351736 305704 351736 305704 0 io_in[36]
rlabel metal2 350728 147420 350728 147420 0 io_in[37]
rlabel metal2 195160 402122 195160 402122 0 io_in[5]
rlabel metal2 289016 53032 289016 53032 0 io_in[6]
rlabel metal3 422408 68824 422408 68824 0 io_in[7]
rlabel metal4 210392 379288 210392 379288 0 io_in[8]
rlabel metal2 471912 398720 471912 398720 0 io_in[9]
rlabel metal3 233912 236264 233912 236264 0 io_oeb[0]
rlabel metal3 188090 255528 188090 255528 0 io_oeb[10]
rlabel metal3 188034 256872 188034 256872 0 io_oeb[11]
rlabel metal3 188146 258216 188146 258216 0 io_oeb[12]
rlabel metal3 593082 549192 593082 549192 0 io_oeb[13]
rlabel metal3 593082 588616 593082 588616 0 io_oeb[14]
rlabel metal2 540568 586362 540568 586362 0 io_oeb[15]
rlabel metal2 474376 587202 474376 587202 0 io_oeb[16]
rlabel metal3 189938 264936 189938 264936 0 io_oeb[17]
rlabel metal3 189770 266280 189770 266280 0 io_oeb[18]
rlabel metal3 189826 267624 189826 267624 0 io_oeb[19]
rlabel metal3 593082 73416 593082 73416 0 io_oeb[1]
rlabel metal2 209608 593474 209608 593474 0 io_oeb[20]
rlabel metal2 143416 503202 143416 503202 0 io_oeb[21]
rlabel metal2 77336 583842 77336 583842 0 io_oeb[22]
rlabel metal2 11032 448602 11032 448602 0 io_oeb[23]
rlabel metal3 2310 558936 2310 558936 0 io_oeb[24]
rlabel metal3 2366 516600 2366 516600 0 io_oeb[25]
rlabel metal3 2422 474264 2422 474264 0 io_oeb[26]
rlabel metal3 183722 278376 183722 278376 0 io_oeb[27]
rlabel metal3 2422 389592 2422 389592 0 io_oeb[28]
rlabel metal3 2310 347256 2310 347256 0 io_oeb[29]
rlabel metal4 190736 231840 190736 231840 0 io_oeb[2]
rlabel metal4 167272 293664 167272 293664 0 io_oeb[30]
rlabel metal3 2310 262808 2310 262808 0 io_oeb[31]
rlabel metal3 190120 285278 190120 285278 0 io_oeb[32]
rlabel metal3 2478 178024 2478 178024 0 io_oeb[33]
rlabel metal3 2534 135800 2534 135800 0 io_oeb[34]
rlabel metal3 2422 93464 2422 93464 0 io_oeb[35]
rlabel metal3 2366 51128 2366 51128 0 io_oeb[36]
rlabel metal3 2310 8792 2310 8792 0 io_oeb[37]
rlabel metal4 304920 240072 304920 240072 0 io_oeb[3]
rlabel metal3 593250 192136 593250 192136 0 io_oeb[4]
rlabel metal3 593194 231896 593194 231896 0 io_oeb[5]
rlabel metal4 355208 192207 355208 192207 0 io_oeb[6]
rlabel metal3 593082 311080 593082 311080 0 io_oeb[7]
rlabel metal2 187208 283080 187208 283080 0 io_oeb[8]
rlabel metal3 593306 390600 593306 390600 0 io_oeb[9]
rlabel metal2 196182 379960 196182 379960 0 io_out[0]
rlabel metal2 204722 379960 204722 379960 0 io_out[10]
rlabel metal4 570360 430323 570360 430323 0 io_out[11]
rlabel metal2 563640 449288 563640 449288 0 io_out[12]
rlabel metal4 565320 470061 565320 470061 0 io_out[13]
rlabel metal2 208446 379960 208446 379960 0 io_out[14]
rlabel metal2 209622 379960 209622 379960 0 io_out[15]
rlabel metal2 210098 379960 210098 379960 0 io_out[16]
rlabel metal2 210994 379960 210994 379960 0 io_out[17]
rlabel metal2 211890 379960 211890 379960 0 io_out[18]
rlabel metal2 212786 379960 212786 379960 0 io_out[19]
rlabel metal2 197078 379960 197078 379960 0 io_out[1]
rlabel metal2 213682 379960 213682 379960 0 io_out[20]
rlabel metal2 214578 379960 214578 379960 0 io_out[21]
rlabel metal2 99512 593082 99512 593082 0 io_out[22]
rlabel metal2 216370 379960 216370 379960 0 io_out[23]
rlabel metal2 217266 379960 217266 379960 0 io_out[24]
rlabel metal2 218162 379960 218162 379960 0 io_out[25]
rlabel metal2 219058 379960 219058 379960 0 io_out[26]
rlabel metal2 219954 379960 219954 379960 0 io_out[27]
rlabel metal3 89838 403704 89838 403704 0 io_out[28]
rlabel metal3 220080 378784 220080 378784 0 io_out[29]
rlabel metal3 590562 99848 590562 99848 0 io_out[2]
rlabel metal2 125272 348992 125272 348992 0 io_out[30]
rlabel metal2 223538 379960 223538 379960 0 io_out[31]
rlabel metal3 65310 234360 65310 234360 0 io_out[32]
rlabel metal3 7350 192024 7350 192024 0 io_out[33]
rlabel metal2 225946 379960 225946 379960 0 io_out[34]
rlabel metal2 29400 243712 29400 243712 0 io_out[35]
rlabel metal2 21000 222432 21000 222432 0 io_out[36]
rlabel metal2 27720 201320 27720 201320 0 io_out[37]
rlabel metal2 198870 379960 198870 379960 0 io_out[3]
rlabel metal4 570360 286245 570360 286245 0 io_out[4]
rlabel metal2 200606 379960 200606 379960 0 io_out[5]
rlabel metal3 593082 258440 593082 258440 0 io_out[6]
rlabel metal2 202034 379960 202034 379960 0 io_out[7]
rlabel metal2 567000 366128 567000 366128 0 io_out[8]
rlabel metal3 593082 377384 593082 377384 0 io_out[9]
rlabel metal3 189434 326760 189434 326760 0 mc14500_do\[0\]
rlabel metal3 188146 340200 188146 340200 0 mc14500_do\[10\]
rlabel metal3 253456 217672 253456 217672 0 mc14500_do\[11\]
rlabel metal3 189602 342888 189602 342888 0 mc14500_do\[12\]
rlabel metal2 326200 214942 326200 214942 0 mc14500_do\[13\]
rlabel metal2 327320 210910 327320 210910 0 mc14500_do\[14\]
rlabel metal3 188202 346920 188202 346920 0 mc14500_do\[15\]
rlabel metal2 329560 212422 329560 212422 0 mc14500_do\[16\]
rlabel metal2 330680 215894 330680 215894 0 mc14500_do\[17\]
rlabel metal2 331800 210014 331800 210014 0 mc14500_do\[18\]
rlabel metal2 332920 213318 332920 213318 0 mc14500_do\[19\]
rlabel metal2 312760 207438 312760 207438 0 mc14500_do\[1\]
rlabel metal2 334040 208166 334040 208166 0 mc14500_do\[20\]
rlabel metal3 189658 354984 189658 354984 0 mc14500_do\[21\]
rlabel metal2 336280 214886 336280 214886 0 mc14500_do\[22\]
rlabel metal2 337400 210798 337400 210798 0 mc14500_do\[23\]
rlabel metal3 188258 359016 188258 359016 0 mc14500_do\[24\]
rlabel metal3 183218 360360 183218 360360 0 mc14500_do\[25\]
rlabel metal3 185682 361704 185682 361704 0 mc14500_do\[26\]
rlabel metal3 260736 234696 260736 234696 0 mc14500_do\[27\]
rlabel metal3 187810 364392 187810 364392 0 mc14500_do\[28\]
rlabel metal3 187362 365736 187362 365736 0 mc14500_do\[29\]
rlabel metal2 313880 207382 313880 207382 0 mc14500_do\[2\]
rlabel metal3 189714 367080 189714 367080 0 mc14500_do\[30\]
rlabel metal3 186410 330792 186410 330792 0 mc14500_do\[3\]
rlabel metal3 187250 332136 187250 332136 0 mc14500_do\[4\]
rlabel metal3 183106 333480 183106 333480 0 mc14500_do\[5\]
rlabel metal3 186354 334824 186354 334824 0 mc14500_do\[6\]
rlabel metal3 189490 336168 189490 336168 0 mc14500_do\[7\]
rlabel metal3 183050 337512 183050 337512 0 mc14500_do\[8\]
rlabel metal3 249816 234136 249816 234136 0 mc14500_do\[9\]
rlabel metal4 237048 376585 237048 376585 0 mc14500_sram_addr\[0\]
rlabel metal2 238238 379400 238238 379400 0 mc14500_sram_addr\[1\]
rlabel metal2 239190 379960 239190 379960 0 mc14500_sram_addr\[2\]
rlabel metal2 239974 379960 239974 379960 0 mc14500_sram_addr\[3\]
rlabel metal2 351176 268408 351176 268408 0 mc14500_sram_addr\[4\]
rlabel metal2 241178 379960 241178 379960 0 mc14500_sram_addr\[5\]
rlabel metal3 261240 379400 261240 379400 0 mc14500_sram_gwe
rlabel metal3 294448 379736 294448 379736 0 mc14500_sram_in\[0\]
rlabel metal2 352856 268128 352856 268128 0 mc14500_sram_in\[1\]
rlabel metal4 349496 270433 349496 270433 0 mc14500_sram_in\[2\]
rlabel metal2 325976 158802 325976 158802 0 mc14500_sram_in\[3\]
rlabel metal2 327544 158914 327544 158914 0 mc14500_sram_in\[4\]
rlabel metal2 246834 379960 246834 379960 0 mc14500_sram_in\[5\]
rlabel metal4 330680 157727 330680 157727 0 mc14500_sram_in\[6\]
rlabel metal4 332248 157637 332248 157637 0 mc14500_sram_in\[7\]
rlabel metal2 275646 379960 275646 379960 0 pdp11_do\[0\]
rlabel metal2 405720 408968 405720 408968 0 pdp11_do\[10\]
rlabel metal2 431704 406434 431704 406434 0 pdp11_do\[11\]
rlabel metal2 297010 379960 297010 379960 0 pdp11_do\[12\]
rlabel metal2 298802 379960 298802 379960 0 pdp11_do\[13\]
rlabel metal2 447832 407274 447832 407274 0 pdp11_do\[14\]
rlabel metal2 302526 379960 302526 379960 0 pdp11_do\[15\]
rlabel metal2 304178 379960 304178 379960 0 pdp11_do\[16\]
rlabel metal2 305970 379960 305970 379960 0 pdp11_do\[17\]
rlabel metal2 307762 379960 307762 379960 0 pdp11_do\[18\]
rlabel metal2 309554 379960 309554 379960 0 pdp11_do\[19\]
rlabel metal2 377944 402290 377944 402290 0 pdp11_do\[1\]
rlabel metal2 311346 379960 311346 379960 0 pdp11_do\[20\]
rlabel metal2 313138 379960 313138 379960 0 pdp11_do\[21\]
rlabel metal2 490840 408898 490840 408898 0 pdp11_do\[22\]
rlabel metal3 493808 406616 493808 406616 0 pdp11_do\[23\]
rlabel metal2 501592 403074 501592 403074 0 pdp11_do\[24\]
rlabel metal2 320306 379960 320306 379960 0 pdp11_do\[25\]
rlabel metal2 322098 379960 322098 379960 0 pdp11_do\[26\]
rlabel metal2 517720 408842 517720 408842 0 pdp11_do\[27\]
rlabel metal2 523096 402906 523096 402906 0 pdp11_do\[28\]
rlabel metal2 327474 379960 327474 379960 0 pdp11_do\[29\]
rlabel metal2 279090 379960 279090 379960 0 pdp11_do\[2\]
rlabel metal2 329406 379960 329406 379960 0 pdp11_do\[30\]
rlabel metal2 331058 379960 331058 379960 0 pdp11_do\[31\]
rlabel metal2 332850 379960 332850 379960 0 pdp11_do\[32\]
rlabel metal2 280882 379960 280882 379960 0 pdp11_do\[3\]
rlabel metal2 282674 379960 282674 379960 0 pdp11_do\[4\]
rlabel metal2 284466 379960 284466 379960 0 pdp11_do\[5\]
rlabel metal2 286678 379960 286678 379960 0 pdp11_do\[6\]
rlabel metal2 288050 379960 288050 379960 0 pdp11_do\[7\]
rlabel metal2 290262 379960 290262 379960 0 pdp11_do\[8\]
rlabel metal2 352184 402584 352184 402584 0 pdp11_do\[9\]
rlabel metal2 276822 379960 276822 379960 0 pdp11_oeb\[0\]
rlabel metal2 294322 379960 294322 379960 0 pdp11_oeb\[10\]
rlabel metal2 296114 379960 296114 379960 0 pdp11_oeb\[11\]
rlabel metal2 297906 379960 297906 379960 0 pdp11_oeb\[12\]
rlabel metal2 299698 379960 299698 379960 0 pdp11_oeb\[13\]
rlabel metal2 301490 379960 301490 379960 0 pdp11_oeb\[14\]
rlabel metal2 303422 379960 303422 379960 0 pdp11_oeb\[15\]
rlabel metal2 305438 379960 305438 379960 0 pdp11_oeb\[16\]
rlabel metal2 307174 379960 307174 379960 0 pdp11_oeb\[17\]
rlabel metal2 308658 379960 308658 379960 0 pdp11_oeb\[18\]
rlabel metal2 310450 379960 310450 379960 0 pdp11_oeb\[19\]
rlabel metal2 278194 379960 278194 379960 0 pdp11_oeb\[1\]
rlabel metal2 312242 379960 312242 379960 0 pdp11_oeb\[20\]
rlabel metal2 314034 379960 314034 379960 0 pdp11_oeb\[21\]
rlabel metal2 315966 379960 315966 379960 0 pdp11_oeb\[22\]
rlabel metal2 318038 379960 318038 379960 0 pdp11_oeb\[23\]
rlabel metal2 319830 379960 319830 379960 0 pdp11_oeb\[24\]
rlabel metal2 321202 379960 321202 379960 0 pdp11_oeb\[25\]
rlabel metal2 323358 379960 323358 379960 0 pdp11_oeb\[26\]
rlabel metal2 324786 379960 324786 379960 0 pdp11_oeb\[27\]
rlabel metal2 326578 379960 326578 379960 0 pdp11_oeb\[28\]
rlabel metal2 328846 379960 328846 379960 0 pdp11_oeb\[29\]
rlabel metal2 279986 379960 279986 379960 0 pdp11_oeb\[2\]
rlabel metal2 330582 379960 330582 379960 0 pdp11_oeb\[30\]
rlabel metal2 332318 379960 332318 379960 0 pdp11_oeb\[31\]
rlabel metal2 334054 379960 334054 379960 0 pdp11_oeb\[32\]
rlabel metal2 281778 379960 281778 379960 0 pdp11_oeb\[3\]
rlabel metal2 283570 379960 283570 379960 0 pdp11_oeb\[4\]
rlabel metal2 285362 379960 285362 379960 0 pdp11_oeb\[5\]
rlabel metal2 287154 379960 287154 379960 0 pdp11_oeb\[6\]
rlabel metal2 289086 379960 289086 379960 0 pdp11_oeb\[7\]
rlabel metal2 290738 379960 290738 379960 0 pdp11_oeb\[8\]
rlabel metal2 292530 379960 292530 379960 0 pdp11_oeb\[9\]
rlabel metal2 350728 180824 350728 180824 0 qcpu_do\[0\]
rlabel metal2 352296 180656 352296 180656 0 qcpu_do\[10\]
rlabel metal2 525448 151606 525448 151606 0 qcpu_do\[11\]
rlabel metal2 305032 197008 305032 197008 0 qcpu_do\[12\]
rlabel metal2 304024 196952 304024 196952 0 qcpu_do\[13\]
rlabel metal2 278936 239106 278936 239106 0 qcpu_do\[14\]
rlabel metal2 279608 238882 279608 238882 0 qcpu_do\[15\]
rlabel metal2 503944 154952 503944 154952 0 qcpu_do\[16\]
rlabel metal2 280952 239162 280952 239162 0 qcpu_do\[17\]
rlabel metal2 505624 152992 505624 152992 0 qcpu_do\[18\]
rlabel metal2 282296 238994 282296 238994 0 qcpu_do\[19\]
rlabel metal2 270424 238504 270424 238504 0 qcpu_do\[1\]
rlabel metal2 537544 152726 537544 152726 0 qcpu_do\[20\]
rlabel metal2 538888 151046 538888 151046 0 qcpu_do\[21\]
rlabel metal2 540232 151494 540232 151494 0 qcpu_do\[22\]
rlabel metal2 541576 151438 541576 151438 0 qcpu_do\[23\]
rlabel via3 501032 149129 501032 149129 0 qcpu_do\[24\]
rlabel metal2 286328 239274 286328 239274 0 qcpu_do\[25\]
rlabel metal2 287000 199738 287000 199738 0 qcpu_do\[26\]
rlabel metal2 287672 199570 287672 199570 0 qcpu_do\[27\]
rlabel metal2 288344 199458 288344 199458 0 qcpu_do\[28\]
rlabel metal2 289016 239218 289016 239218 0 qcpu_do\[29\]
rlabel metal2 513352 154630 513352 154630 0 qcpu_do\[2\]
rlabel metal2 289688 199514 289688 199514 0 qcpu_do\[30\]
rlabel metal2 290360 200970 290360 200970 0 qcpu_do\[31\]
rlabel metal2 291032 195370 291032 195370 0 qcpu_do\[32\]
rlabel metal2 514696 151102 514696 151102 0 qcpu_do\[3\]
rlabel metal2 355544 189952 355544 189952 0 qcpu_do\[4\]
rlabel metal2 310632 185416 310632 185416 0 qcpu_do\[5\]
rlabel metal2 310408 185640 310408 185640 0 qcpu_do\[6\]
rlabel metal2 520072 155134 520072 155134 0 qcpu_do\[7\]
rlabel metal2 521416 155302 521416 155302 0 qcpu_do\[8\]
rlabel metal2 522760 155246 522760 155246 0 qcpu_do\[9\]
rlabel metal3 350392 209944 350392 209944 0 qcpu_oeb\[0\]
rlabel metal2 563416 60480 563416 60480 0 qcpu_oeb\[10\]
rlabel metal4 353752 183344 353752 183344 0 qcpu_oeb\[11\]
rlabel metal4 559496 123872 559496 123872 0 qcpu_oeb\[12\]
rlabel metal5 342832 193230 342832 193230 0 qcpu_oeb\[13\]
rlabel metal4 350840 183600 350840 183600 0 qcpu_oeb\[14\]
rlabel metal2 562968 114576 562968 114576 0 qcpu_oeb\[15\]
rlabel metal2 563528 63560 563528 63560 0 qcpu_oeb\[16\]
rlabel metal4 353640 183624 353640 183624 0 qcpu_oeb\[17\]
rlabel metal4 350728 250488 350728 250488 0 qcpu_oeb\[18\]
rlabel metal2 563080 117656 563080 117656 0 qcpu_oeb\[19\]
rlabel metal3 355376 280392 355376 280392 0 qcpu_oeb\[1\]
rlabel metal2 563192 119336 563192 119336 0 qcpu_oeb\[20\]
rlabel metal4 352408 247296 352408 247296 0 qcpu_oeb\[21\]
rlabel metal4 563528 120848 563528 120848 0 qcpu_oeb\[22\]
rlabel metal4 350504 247352 350504 247352 0 qcpu_oeb\[23\]
rlabel metal4 353976 240520 353976 240520 0 qcpu_oeb\[24\]
rlabel metal3 348068 167048 348068 167048 0 qcpu_oeb\[25\]
rlabel metal4 562968 130648 562968 130648 0 qcpu_oeb\[26\]
rlabel metal4 563752 125832 563752 125832 0 qcpu_oeb\[27\]
rlabel metal4 352296 248752 352296 248752 0 qcpu_oeb\[28\]
rlabel metal4 350392 247520 350392 247520 0 qcpu_oeb\[29\]
rlabel metal3 351960 191688 351960 191688 0 qcpu_oeb\[2\]
rlabel metal4 355656 248864 355656 248864 0 qcpu_oeb\[30\]
rlabel metal4 561176 139563 561176 139563 0 qcpu_oeb\[31\]
rlabel metal4 354088 252168 354088 252168 0 qcpu_oeb\[32\]
rlabel metal2 563640 54712 563640 54712 0 qcpu_oeb\[3\]
rlabel metal2 563304 56672 563304 56672 0 qcpu_oeb\[4\]
rlabel metal4 355320 179704 355320 179704 0 qcpu_oeb\[5\]
rlabel metal4 351960 181160 351960 181160 0 qcpu_oeb\[6\]
rlabel metal3 353640 282184 353640 282184 0 qcpu_oeb\[7\]
rlabel metal3 350280 193256 350280 193256 0 qcpu_oeb\[8\]
rlabel metal4 352968 150857 352968 150857 0 qcpu_oeb\[9\]
rlabel metal2 561512 129416 561512 129416 0 qcpu_sram_addr\[0\]
rlabel metal4 564536 134355 564536 134355 0 qcpu_sram_addr\[1\]
rlabel metal3 426720 162120 426720 162120 0 qcpu_sram_addr\[2\]
rlabel metal4 564648 136823 564648 136823 0 qcpu_sram_addr\[3\]
rlabel metal2 561624 133392 561624 133392 0 qcpu_sram_addr\[4\]
rlabel metal4 564760 135871 564760 135871 0 qcpu_sram_addr\[5\]
rlabel metal2 561288 146216 561288 146216 0 qcpu_sram_gwe
rlabel metal3 387604 149240 387604 149240 0 qcpu_sram_in\[0\]
rlabel metal2 564648 137424 564648 137424 0 qcpu_sram_in\[1\]
rlabel metal4 566216 140833 566216 140833 0 qcpu_sram_in\[2\]
rlabel metal2 564536 142296 564536 142296 0 qcpu_sram_in\[3\]
rlabel metal3 559608 124278 559608 124278 0 qcpu_sram_in\[4\]
rlabel metal4 561288 142285 561288 142285 0 qcpu_sram_in\[5\]
rlabel metal2 561400 143024 561400 143024 0 qcpu_sram_in\[6\]
rlabel metal2 566216 144648 566216 144648 0 qcpu_sram_in\[7\]
rlabel metal2 333816 158690 333816 158690 0 qcpu_sram_out\[0\]
rlabel metal2 335384 158970 335384 158970 0 qcpu_sram_out\[1\]
rlabel metal2 336952 158802 336952 158802 0 qcpu_sram_out\[2\]
rlabel metal2 357896 158256 357896 158256 0 qcpu_sram_out\[3\]
rlabel metal2 352520 158592 352520 158592 0 qcpu_sram_out\[4\]
rlabel metal2 354536 176792 354536 176792 0 qcpu_sram_out\[5\]
rlabel metal5 345184 191610 345184 191610 0 qcpu_sram_out\[6\]
rlabel metal2 350728 158648 350728 158648 0 qcpu_sram_out\[7\]
rlabel metal3 63112 304024 63112 304024 0 rst_ay8913
rlabel metal2 232386 379960 232386 379960 0 rst_blinker
rlabel metal2 152824 303926 152824 303926 0 rst_hellorld
rlabel metal4 349720 180796 349720 180796 0 rst_mc14500
rlabel metal3 190680 421806 190680 421806 0 rst_pdp11
rlabel metal3 190680 323722 190680 323722 0 rst_qcpu
rlabel metal2 212296 48874 212296 48874 0 rst_sid
rlabel via4 236152 379723 236152 379723 0 rst_sn76489
rlabel metal3 182280 358680 182280 358680 0 rst_tbb1143
rlabel metal2 335118 379960 335118 379960 0 rst_tholin_riscv
rlabel metal3 188818 294504 188818 294504 0 sid_do\[0\]
rlabel metal3 187922 307944 187922 307944 0 sid_do\[10\]
rlabel metal3 271334 180824 271334 180824 0 sid_do\[11\]
rlabel metal3 187978 310632 187978 310632 0 sid_do\[12\]
rlabel metal3 182210 311976 182210 311976 0 sid_do\[13\]
rlabel metal3 184058 313320 184058 313320 0 sid_do\[14\]
rlabel metal3 271334 192472 271334 192472 0 sid_do\[15\]
rlabel metal3 271446 195384 271446 195384 0 sid_do\[16\]
rlabel metal3 225400 219688 225400 219688 0 sid_do\[17\]
rlabel metal4 174440 265720 174440 265720 0 sid_do\[18\]
rlabel metal4 174664 264824 174664 264824 0 sid_do\[19\]
rlabel metal3 188762 295848 188762 295848 0 sid_do\[1\]
rlabel metal4 174552 267120 174552 267120 0 sid_do\[20\]
rlabel metal3 188874 297192 188874 297192 0 sid_do\[2\]
rlabel metal3 188594 298536 188594 298536 0 sid_do\[3\]
rlabel metal3 186522 299880 186522 299880 0 sid_do\[4\]
rlabel metal3 188482 301224 188482 301224 0 sid_do\[5\]
rlabel metal3 188538 302568 188538 302568 0 sid_do\[6\]
rlabel metal3 188930 303912 188930 303912 0 sid_do\[7\]
rlabel metal3 187306 305256 187306 305256 0 sid_do\[8\]
rlabel metal3 185682 306600 185682 306600 0 sid_do\[9\]
rlabel metal4 187432 322689 187432 322689 0 sid_oeb
rlabel metal2 250712 238098 250712 238098 0 sn76489_do\[0\]
rlabel metal2 382872 121870 382872 121870 0 sn76489_do\[10\]
rlabel metal2 258104 234738 258104 234738 0 sn76489_do\[11\]
rlabel metal2 258776 225722 258776 225722 0 sn76489_do\[12\]
rlabel metal2 259448 233282 259448 233282 0 sn76489_do\[13\]
rlabel metal2 260120 238322 260120 238322 0 sn76489_do\[14\]
rlabel metal2 260792 225778 260792 225778 0 sn76489_do\[15\]
rlabel metal2 261464 227066 261464 227066 0 sn76489_do\[16\]
rlabel metal2 306936 170744 306936 170744 0 sn76489_do\[17\]
rlabel metal2 306712 170744 306712 170744 0 sn76489_do\[18\]
rlabel metal2 307160 172592 307160 172592 0 sn76489_do\[19\]
rlabel metal2 251384 238210 251384 238210 0 sn76489_do\[1\]
rlabel metal2 264152 228802 264152 228802 0 sn76489_do\[20\]
rlabel metal2 264824 229138 264824 229138 0 sn76489_do\[21\]
rlabel metal2 303128 173432 303128 173432 0 sn76489_do\[22\]
rlabel metal2 266168 229194 266168 229194 0 sn76489_do\[23\]
rlabel metal2 266840 228746 266840 228746 0 sn76489_do\[24\]
rlabel metal3 268128 237048 268128 237048 0 sn76489_do\[25\]
rlabel metal2 268632 238504 268632 238504 0 sn76489_do\[26\]
rlabel metal2 269094 240072 269094 240072 0 sn76489_do\[27\]
rlabel metal2 308280 168784 308280 168784 0 sn76489_do\[2\]
rlabel metal2 303352 170016 303352 170016 0 sn76489_do\[3\]
rlabel metal2 306600 173712 306600 173712 0 sn76489_do\[4\]
rlabel metal2 372792 121758 372792 121758 0 sn76489_do\[5\]
rlabel metal2 374808 121814 374808 121814 0 sn76489_do\[6\]
rlabel metal2 255416 230650 255416 230650 0 sn76489_do\[7\]
rlabel metal2 256088 230706 256088 230706 0 sn76489_do\[8\]
rlabel metal2 380856 121702 380856 121702 0 sn76489_do\[9\]
rlabel metal3 175896 349958 175896 349958 0 tbb1143_do\[0\]
rlabel metal3 178318 352968 178318 352968 0 tbb1143_do\[1\]
rlabel metal3 180054 356328 180054 356328 0 tbb1143_do\[2\]
rlabel metal3 181678 359688 181678 359688 0 tbb1143_do\[3\]
rlabel metal3 179214 363048 179214 363048 0 tbb1143_do\[4\]
rlabel metal2 355880 189000 355880 189000 0 tholin_riscv_do\[0\]
rlabel metal2 423640 173866 423640 173866 0 tholin_riscv_do\[10\]
rlabel metal2 429688 173810 429688 173810 0 tholin_riscv_do\[11\]
rlabel metal2 350392 264432 350392 264432 0 tholin_riscv_do\[12\]
rlabel metal2 353752 263928 353752 263928 0 tholin_riscv_do\[13\]
rlabel metal2 355432 265384 355432 265384 0 tholin_riscv_do\[14\]
rlabel metal2 354200 185136 354200 185136 0 tholin_riscv_do\[15\]
rlabel metal2 352072 265328 352072 265328 0 tholin_riscv_do\[16\]
rlabel metal3 342678 360584 342678 360584 0 tholin_riscv_do\[17\]
rlabel metal2 472024 173082 472024 173082 0 tholin_riscv_do\[18\]
rlabel metal2 478072 172242 478072 172242 0 tholin_riscv_do\[19\]
rlabel metal2 354088 260736 354088 260736 0 tholin_riscv_do\[1\]
rlabel metal5 351960 192330 351960 192330 0 tholin_riscv_do\[20\]
rlabel metal4 359800 193979 359800 193979 0 tholin_riscv_do\[21\]
rlabel metal2 350280 267288 350280 267288 0 tholin_riscv_do\[22\]
rlabel metal2 353640 266784 353640 266784 0 tholin_riscv_do\[23\]
rlabel metal2 355320 267288 355320 267288 0 tholin_riscv_do\[24\]
rlabel metal2 351960 268688 351960 268688 0 tholin_riscv_do\[25\]
rlabel metal2 520408 174818 520408 174818 0 tholin_riscv_do\[26\]
rlabel metal2 346976 167832 346976 167832 0 tholin_riscv_do\[27\]
rlabel metal3 344246 370440 344246 370440 0 tholin_riscv_do\[28\]
rlabel metal2 538552 174034 538552 174034 0 tholin_riscv_do\[29\]
rlabel via4 375256 175227 375256 175227 0 tholin_riscv_do\[2\]
rlabel metal2 544600 173978 544600 173978 0 tholin_riscv_do\[30\]
rlabel metal3 342006 373128 342006 373128 0 tholin_riscv_do\[31\]
rlabel metal2 562856 283192 562856 283192 0 tholin_riscv_do\[32\]
rlabel metal2 355656 260176 355656 260176 0 tholin_riscv_do\[3\]
rlabel metal2 352184 261296 352184 261296 0 tholin_riscv_do\[4\]
rlabel metal3 344470 349832 344470 349832 0 tholin_riscv_do\[5\]
rlabel metal4 352744 183811 352744 183811 0 tholin_riscv_do\[6\]
rlabel metal2 405496 173754 405496 173754 0 tholin_riscv_do\[7\]
rlabel metal3 344414 352520 344414 352520 0 tholin_riscv_do\[8\]
rlabel metal3 342566 353416 342566 353416 0 tholin_riscv_do\[9\]
rlabel metal2 301784 236754 301784 236754 0 tholin_riscv_oeb\[0\]
rlabel metal2 312536 236264 312536 236264 0 tholin_riscv_oeb\[10\]
rlabel metal3 359912 389256 359912 389256 0 tholin_riscv_oeb\[11\]
rlabel metal4 359912 389545 359912 389545 0 tholin_riscv_oeb\[12\]
rlabel metal3 326256 237720 326256 237720 0 tholin_riscv_oeb\[13\]
rlabel metal2 350728 316120 350728 316120 0 tholin_riscv_oeb\[14\]
rlabel metal3 328608 237832 328608 237832 0 tholin_riscv_oeb\[15\]
rlabel metal2 354200 321664 354200 321664 0 tholin_riscv_oeb\[16\]
rlabel metal3 334992 238392 334992 238392 0 tholin_riscv_oeb\[17\]
rlabel metal2 472024 401646 472024 401646 0 tholin_riscv_oeb\[18\]
rlabel metal2 350504 320656 350504 320656 0 tholin_riscv_oeb\[19\]
rlabel metal2 302456 234234 302456 234234 0 tholin_riscv_oeb\[1\]
rlabel metal4 359576 398888 359576 398888 0 tholin_riscv_oeb\[20\]
rlabel metal2 352296 319928 352296 319928 0 tholin_riscv_oeb\[21\]
rlabel via3 359912 388905 359912 388905 0 tholin_riscv_oeb\[22\]
rlabel metal2 502264 399966 502264 399966 0 tholin_riscv_oeb\[23\]
rlabel metal2 508312 395822 508312 395822 0 tholin_riscv_oeb\[24\]
rlabel metal2 514360 396270 514360 396270 0 tholin_riscv_oeb\[25\]
rlabel metal3 519792 398104 519792 398104 0 tholin_riscv_oeb\[26\]
rlabel metal4 526456 397021 526456 397021 0 tholin_riscv_oeb\[27\]
rlabel metal4 353528 318600 353528 318600 0 tholin_riscv_oeb\[28\]
rlabel metal4 354424 316260 354424 316260 0 tholin_riscv_oeb\[29\]
rlabel metal2 375256 396158 375256 396158 0 tholin_riscv_oeb\[2\]
rlabel metal2 544600 398342 544600 398342 0 tholin_riscv_oeb\[30\]
rlabel metal4 550648 396583 550648 396583 0 tholin_riscv_oeb\[31\]
rlabel metal4 355880 319770 355880 319770 0 tholin_riscv_oeb\[32\]
rlabel metal2 303800 238154 303800 238154 0 tholin_riscv_oeb\[3\]
rlabel metal2 304472 238266 304472 238266 0 tholin_riscv_oeb\[4\]
rlabel metal2 305144 238378 305144 238378 0 tholin_riscv_oeb\[5\]
rlabel metal2 305816 238210 305816 238210 0 tholin_riscv_oeb\[6\]
rlabel metal2 306488 238826 306488 238826 0 tholin_riscv_oeb\[7\]
rlabel metal2 307160 238098 307160 238098 0 tholin_riscv_oeb\[8\]
rlabel metal2 307832 238042 307832 238042 0 tholin_riscv_oeb\[9\]
rlabel metal2 230006 379960 230006 379960 0 user_irq[0]
rlabel metal2 231182 379960 231182 379960 0 user_irq[1]
rlabel metal2 231742 379960 231742 379960 0 user_irq[2]
rlabel metal2 97384 48986 97384 48986 0 wb_clk_i
rlabel metal2 13272 114926 13272 114926 0 wb_rst_i
rlabel metal2 15400 2310 15400 2310 0 wbs_ack_o
rlabel metal2 22792 116550 22792 116550 0 wbs_adr_i[0]
rlabel metal4 48552 144200 48552 144200 0 wbs_adr_i[10]
rlabel metal2 215096 237314 215096 237314 0 wbs_adr_i[11]
rlabel metal2 215768 237258 215768 237258 0 wbs_adr_i[12]
rlabel metal2 216440 237258 216440 237258 0 wbs_adr_i[13]
rlabel metal2 217112 237314 217112 237314 0 wbs_adr_i[14]
rlabel metal2 218344 238504 218344 238504 0 wbs_adr_i[15]
rlabel metal3 219240 237048 219240 237048 0 wbs_adr_i[16]
rlabel metal2 219128 235746 219128 235746 0 wbs_adr_i[17]
rlabel metal2 219800 235858 219800 235858 0 wbs_adr_i[18]
rlabel metal2 138936 24318 138936 24318 0 wbs_adr_i[19]
rlabel metal2 30408 114030 30408 114030 0 wbs_adr_i[1]
rlabel metal2 144648 22694 144648 22694 0 wbs_adr_i[20]
rlabel metal2 150360 20958 150360 20958 0 wbs_adr_i[21]
rlabel metal2 156072 21014 156072 21014 0 wbs_adr_i[22]
rlabel metal2 161784 21070 161784 21070 0 wbs_adr_i[23]
rlabel metal2 167496 22750 167496 22750 0 wbs_adr_i[24]
rlabel metal2 173208 21126 173208 21126 0 wbs_adr_i[25]
rlabel metal2 225176 237594 225176 237594 0 wbs_adr_i[26]
rlabel metal2 225848 237146 225848 237146 0 wbs_adr_i[27]
rlabel metal2 190344 24430 190344 24430 0 wbs_adr_i[28]
rlabel metal2 196056 20734 196056 20734 0 wbs_adr_i[29]
rlabel metal2 209048 231434 209048 231434 0 wbs_adr_i[2]
rlabel metal2 227864 238266 227864 238266 0 wbs_adr_i[30]
rlabel metal3 239400 47768 239400 47768 0 wbs_adr_i[31]
rlabel metal2 45640 2702 45640 2702 0 wbs_adr_i[3]
rlabel metal3 50120 49560 50120 49560 0 wbs_adr_i[4]
rlabel metal2 211064 229642 211064 229642 0 wbs_adr_i[5]
rlabel metal2 211736 225442 211736 225442 0 wbs_adr_i[6]
rlabel metal2 70392 2534 70392 2534 0 wbs_adr_i[7]
rlabel metal2 76104 2702 76104 2702 0 wbs_adr_i[8]
rlabel metal4 48664 114352 48664 114352 0 wbs_adr_i[9]
rlabel metal2 17304 2310 17304 2310 0 wbs_cyc_i
rlabel metal2 24920 2310 24920 2310 0 wbs_dat_i[0]
rlabel metal4 235928 235861 235928 235861 0 wbs_dat_i[10]
rlabel metal2 236824 238504 236824 238504 0 wbs_dat_i[11]
rlabel metal2 100856 20846 100856 20846 0 wbs_dat_i[12]
rlabel metal2 237944 233786 237944 233786 0 wbs_dat_i[13]
rlabel metal2 238616 224994 238616 224994 0 wbs_dat_i[14]
rlabel metal2 117992 19278 117992 19278 0 wbs_dat_i[15]
rlabel metal2 123704 25046 123704 25046 0 wbs_dat_i[16]
rlabel metal2 240632 236362 240632 236362 0 wbs_dat_i[17]
rlabel metal2 241304 232162 241304 232162 0 wbs_dat_i[18]
rlabel metal4 241976 237737 241976 237737 0 wbs_dat_i[19]
rlabel metal3 131096 214200 131096 214200 0 wbs_dat_i[1]
rlabel metal2 146776 3990 146776 3990 0 wbs_dat_i[20]
rlabel metal2 243320 239218 243320 239218 0 wbs_dat_i[21]
rlabel metal2 158200 3150 158200 3150 0 wbs_dat_i[22]
rlabel metal2 163688 6510 163688 6510 0 wbs_dat_i[23]
rlabel metal2 169400 14910 169400 14910 0 wbs_dat_i[24]
rlabel metal2 246008 238994 246008 238994 0 wbs_dat_i[25]
rlabel metal2 181048 2646 181048 2646 0 wbs_dat_i[26]
rlabel metal2 186536 24374 186536 24374 0 wbs_dat_i[27]
rlabel metal2 192248 12558 192248 12558 0 wbs_dat_i[28]
rlabel metal2 248696 239050 248696 239050 0 wbs_dat_i[29]
rlabel metal2 39928 111566 39928 111566 0 wbs_dat_i[2]
rlabel metal2 249368 239106 249368 239106 0 wbs_dat_i[30]
rlabel metal2 209608 2254 209608 2254 0 wbs_dat_i[31]
rlabel metal2 47544 2310 47544 2310 0 wbs_dat_i[3]
rlabel metal4 55160 4093 55160 4093 0 wbs_dat_i[4]
rlabel metal2 232568 226282 232568 226282 0 wbs_dat_i[5]
rlabel metal4 233240 235861 233240 235861 0 wbs_dat_i[6]
rlabel metal2 72296 2478 72296 2478 0 wbs_dat_i[7]
rlabel metal2 78008 2590 78008 2590 0 wbs_dat_i[8]
rlabel metal4 52024 114296 52024 114296 0 wbs_dat_i[9]
rlabel metal2 26600 111510 26600 111510 0 wbs_dat_o[0]
rlabel metal2 91560 1918 91560 1918 0 wbs_dat_o[10]
rlabel metal2 97048 17430 97048 17430 0 wbs_dat_o[11]
rlabel metal2 286888 130256 286888 130256 0 wbs_dat_o[12]
rlabel metal2 286440 130368 286440 130368 0 wbs_dat_o[13]
rlabel metal2 114408 2534 114408 2534 0 wbs_dat_o[14]
rlabel metal2 119896 15750 119896 15750 0 wbs_dat_o[15]
rlabel metal2 125608 17598 125608 17598 0 wbs_dat_o[16]
rlabel metal3 207200 31192 207200 31192 0 wbs_dat_o[17]
rlabel metal2 137032 19334 137032 19334 0 wbs_dat_o[18]
rlabel metal2 142968 1918 142968 1918 0 wbs_dat_o[19]
rlabel metal4 329224 230711 329224 230711 0 wbs_dat_o[1]
rlabel metal2 148456 22638 148456 22638 0 wbs_dat_o[20]
rlabel metal2 154392 2366 154392 2366 0 wbs_dat_o[21]
rlabel metal2 354648 246624 354648 246624 0 wbs_dat_o[22]
rlabel metal2 165816 2422 165816 2422 0 wbs_dat_o[23]
rlabel metal2 171528 2254 171528 2254 0 wbs_dat_o[24]
rlabel metal2 351400 254520 351400 254520 0 wbs_dat_o[25]
rlabel metal2 182952 2478 182952 2478 0 wbs_dat_o[26]
rlabel metal2 188440 15918 188440 15918 0 wbs_dat_o[27]
rlabel metal2 194376 2590 194376 2590 0 wbs_dat_o[28]
rlabel metal2 349608 256368 349608 256368 0 wbs_dat_o[29]
rlabel metal3 309344 219800 309344 219800 0 wbs_dat_o[2]
rlabel metal4 288232 240240 288232 240240 0 wbs_dat_o[30]
rlabel metal2 211512 2534 211512 2534 0 wbs_dat_o[31]
rlabel metal2 49448 2366 49448 2366 0 wbs_dat_o[3]
rlabel metal4 311864 134235 311864 134235 0 wbs_dat_o[4]
rlabel metal4 309960 128632 309960 128632 0 wbs_dat_o[5]
rlabel metal2 68488 12446 68488 12446 0 wbs_dat_o[6]
rlabel metal2 74200 12390 74200 12390 0 wbs_dat_o[7]
rlabel metal3 177296 24584 177296 24584 0 wbs_dat_o[8]
rlabel metal4 311640 134471 311640 134471 0 wbs_dat_o[9]
rlabel metal2 19208 2310 19208 2310 0 wbs_stb_i
rlabel metal2 20888 114870 20888 114870 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
