magic
tech gf180mcuD
magscale 1 10
timestamp 1712517911
<< metal1 >>
rect 5506 47966 5518 48018
rect 5570 48015 5582 48018
rect 6514 48015 6526 48018
rect 5570 47969 6526 48015
rect 5570 47966 5582 47969
rect 6514 47966 6526 47969
rect 6578 47966 6590 48018
rect 30818 47966 30830 48018
rect 30882 48015 30894 48018
rect 31602 48015 31614 48018
rect 30882 47969 31614 48015
rect 30882 47966 30894 47969
rect 31602 47966 31614 47969
rect 31666 47966 31678 48018
rect 34066 47966 34078 48018
rect 34130 48015 34142 48018
rect 35074 48015 35086 48018
rect 34130 47969 35086 48015
rect 34130 47966 34142 47969
rect 35074 47966 35086 47969
rect 35138 47966 35150 48018
rect 1344 47850 49616 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 49616 47850
rect 1344 47764 49616 47798
rect 6526 47682 6578 47694
rect 6526 47618 6578 47630
rect 42366 47682 42418 47694
rect 42366 47618 42418 47630
rect 45390 47682 45442 47694
rect 45390 47618 45442 47630
rect 19070 47570 19122 47582
rect 19070 47506 19122 47518
rect 30830 47570 30882 47582
rect 40574 47570 40626 47582
rect 35074 47518 35086 47570
rect 35138 47518 35150 47570
rect 44482 47518 44494 47570
rect 44546 47518 44558 47570
rect 48738 47518 48750 47570
rect 48802 47518 48814 47570
rect 30830 47506 30882 47518
rect 40574 47506 40626 47518
rect 19294 47458 19346 47470
rect 19294 47394 19346 47406
rect 31614 47458 31666 47470
rect 40014 47458 40066 47470
rect 42142 47458 42194 47470
rect 32162 47406 32174 47458
rect 32226 47406 32238 47458
rect 41906 47406 41918 47458
rect 41970 47406 41982 47458
rect 31614 47394 31666 47406
rect 40014 47394 40066 47406
rect 42142 47394 42194 47406
rect 42814 47458 42866 47470
rect 45614 47458 45666 47470
rect 47742 47458 47794 47470
rect 43698 47406 43710 47458
rect 43762 47406 43774 47458
rect 44818 47406 44830 47458
rect 44882 47406 44894 47458
rect 45826 47406 45838 47458
rect 45890 47406 45902 47458
rect 46386 47406 46398 47458
rect 46450 47406 46462 47458
rect 48178 47406 48190 47458
rect 48242 47406 48254 47458
rect 49074 47406 49086 47458
rect 49138 47406 49150 47458
rect 42814 47394 42866 47406
rect 45614 47394 45666 47406
rect 47742 47394 47794 47406
rect 6862 47346 6914 47358
rect 6862 47282 6914 47294
rect 19854 47346 19906 47358
rect 19854 47282 19906 47294
rect 26574 47346 26626 47358
rect 26574 47282 26626 47294
rect 29710 47346 29762 47358
rect 29710 47282 29762 47294
rect 31054 47346 31106 47358
rect 36318 47346 36370 47358
rect 32946 47294 32958 47346
rect 33010 47294 33022 47346
rect 31054 47282 31106 47294
rect 36318 47282 36370 47294
rect 38782 47346 38834 47358
rect 38782 47282 38834 47294
rect 41582 47346 41634 47358
rect 41582 47282 41634 47294
rect 45278 47346 45330 47358
rect 45278 47282 45330 47294
rect 6638 47234 6690 47246
rect 6638 47170 6690 47182
rect 26238 47234 26290 47246
rect 26238 47170 26290 47182
rect 29374 47234 29426 47246
rect 29374 47170 29426 47182
rect 35982 47234 36034 47246
rect 35982 47170 36034 47182
rect 36878 47234 36930 47246
rect 36878 47170 36930 47182
rect 37438 47234 37490 47246
rect 37438 47170 37490 47182
rect 37774 47234 37826 47246
rect 37774 47170 37826 47182
rect 38334 47234 38386 47246
rect 38334 47170 38386 47182
rect 39230 47234 39282 47246
rect 39230 47170 39282 47182
rect 41022 47234 41074 47246
rect 41022 47170 41074 47182
rect 41358 47234 41410 47246
rect 41358 47170 41410 47182
rect 41470 47234 41522 47246
rect 41470 47170 41522 47182
rect 42030 47234 42082 47246
rect 42030 47170 42082 47182
rect 42926 47234 42978 47246
rect 46174 47234 46226 47246
rect 43922 47182 43934 47234
rect 43986 47182 43998 47234
rect 42926 47170 42978 47182
rect 46174 47170 46226 47182
rect 1344 47066 49616 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 49616 47066
rect 1344 46980 49616 47014
rect 32398 46898 32450 46910
rect 32398 46834 32450 46846
rect 33742 46898 33794 46910
rect 33742 46834 33794 46846
rect 34190 46898 34242 46910
rect 34190 46834 34242 46846
rect 8430 46786 8482 46798
rect 47518 46786 47570 46798
rect 5506 46734 5518 46786
rect 5570 46734 5582 46786
rect 26002 46734 26014 46786
rect 26066 46734 26078 46786
rect 29586 46734 29598 46786
rect 29650 46734 29662 46786
rect 35186 46734 35198 46786
rect 35250 46734 35262 46786
rect 41682 46734 41694 46786
rect 41746 46734 41758 46786
rect 45042 46734 45054 46786
rect 45106 46734 45118 46786
rect 8430 46722 8482 46734
rect 47518 46722 47570 46734
rect 48750 46786 48802 46798
rect 48750 46722 48802 46734
rect 32062 46674 32114 46686
rect 47854 46674 47906 46686
rect 6290 46622 6302 46674
rect 6354 46622 6366 46674
rect 7074 46622 7086 46674
rect 7138 46622 7150 46674
rect 8082 46622 8094 46674
rect 8146 46622 8158 46674
rect 21634 46622 21646 46674
rect 21698 46622 21710 46674
rect 25218 46622 25230 46674
rect 25282 46622 25294 46674
rect 28914 46622 28926 46674
rect 28978 46622 28990 46674
rect 34402 46622 34414 46674
rect 34466 46622 34478 46674
rect 41010 46622 41022 46674
rect 41074 46622 41086 46674
rect 44370 46622 44382 46674
rect 44434 46622 44446 46674
rect 48962 46622 48974 46674
rect 49026 46622 49038 46674
rect 32062 46610 32114 46622
rect 47854 46610 47906 46622
rect 6750 46562 6802 46574
rect 37886 46562 37938 46574
rect 3378 46510 3390 46562
rect 3442 46510 3454 46562
rect 7298 46510 7310 46562
rect 7362 46510 7374 46562
rect 8194 46510 8206 46562
rect 8258 46510 8270 46562
rect 18834 46510 18846 46562
rect 18898 46510 18910 46562
rect 20962 46510 20974 46562
rect 21026 46510 21038 46562
rect 28130 46510 28142 46562
rect 28194 46510 28206 46562
rect 31714 46510 31726 46562
rect 31778 46510 31790 46562
rect 37314 46510 37326 46562
rect 37378 46510 37390 46562
rect 6750 46498 6802 46510
rect 37886 46498 37938 46510
rect 38334 46562 38386 46574
rect 38334 46498 38386 46510
rect 38894 46562 38946 46574
rect 38894 46498 38946 46510
rect 39342 46562 39394 46574
rect 39342 46498 39394 46510
rect 39790 46562 39842 46574
rect 39790 46498 39842 46510
rect 40462 46562 40514 46574
rect 43810 46510 43822 46562
rect 43874 46510 43886 46562
rect 47170 46510 47182 46562
rect 47234 46510 47246 46562
rect 40462 46498 40514 46510
rect 37998 46450 38050 46462
rect 37998 46386 38050 46398
rect 38446 46450 38498 46462
rect 38658 46398 38670 46450
rect 38722 46447 38734 46450
rect 38882 46447 38894 46450
rect 38722 46401 38894 46447
rect 38722 46398 38734 46401
rect 38882 46398 38894 46401
rect 38946 46398 38958 46450
rect 38446 46386 38498 46398
rect 1344 46282 49616 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 49616 46282
rect 1344 46196 49616 46230
rect 44270 46114 44322 46126
rect 27010 46062 27022 46114
rect 27074 46062 27086 46114
rect 29698 46062 29710 46114
rect 29762 46062 29774 46114
rect 30258 46062 30270 46114
rect 30322 46062 30334 46114
rect 41234 46062 41246 46114
rect 41298 46062 41310 46114
rect 44270 46050 44322 46062
rect 44158 46002 44210 46014
rect 10546 45950 10558 46002
rect 10610 45950 10622 46002
rect 31938 45950 31950 46002
rect 32002 45950 32014 46002
rect 38434 45950 38446 46002
rect 38498 45950 38510 46002
rect 40562 45950 40574 46002
rect 40626 45950 40638 46002
rect 46274 45950 46286 46002
rect 46338 45950 46350 46002
rect 44158 45938 44210 45950
rect 4510 45890 4562 45902
rect 4510 45826 4562 45838
rect 4734 45890 4786 45902
rect 7086 45890 7138 45902
rect 26574 45890 26626 45902
rect 4946 45838 4958 45890
rect 5010 45838 5022 45890
rect 5842 45838 5854 45890
rect 5906 45838 5918 45890
rect 7746 45838 7758 45890
rect 7810 45838 7822 45890
rect 4734 45826 4786 45838
rect 7086 45826 7138 45838
rect 26574 45826 26626 45838
rect 27358 45890 27410 45902
rect 27358 45826 27410 45838
rect 27582 45890 27634 45902
rect 27582 45826 27634 45838
rect 29150 45890 29202 45902
rect 29150 45826 29202 45838
rect 29374 45890 29426 45902
rect 29374 45826 29426 45838
rect 30606 45890 30658 45902
rect 30606 45826 30658 45838
rect 30830 45890 30882 45902
rect 41582 45890 41634 45902
rect 36418 45838 36430 45890
rect 36482 45838 36494 45890
rect 37314 45838 37326 45890
rect 37378 45838 37390 45890
rect 37650 45838 37662 45890
rect 37714 45838 37726 45890
rect 30830 45826 30882 45838
rect 41582 45826 41634 45838
rect 41806 45890 41858 45902
rect 45390 45890 45442 45902
rect 42690 45838 42702 45890
rect 42754 45838 42766 45890
rect 43026 45838 43038 45890
rect 43090 45838 43102 45890
rect 43922 45838 43934 45890
rect 43986 45838 43998 45890
rect 41806 45826 41858 45838
rect 45390 45826 45442 45838
rect 45726 45890 45778 45902
rect 45726 45826 45778 45838
rect 45838 45890 45890 45902
rect 49074 45838 49086 45890
rect 49138 45838 49150 45890
rect 45838 45826 45890 45838
rect 4398 45778 4450 45790
rect 4398 45714 4450 45726
rect 6750 45778 6802 45790
rect 6750 45714 6802 45726
rect 7198 45778 7250 45790
rect 7198 45714 7250 45726
rect 7310 45778 7362 45790
rect 26686 45778 26738 45790
rect 8418 45726 8430 45778
rect 8482 45726 8494 45778
rect 7310 45714 7362 45726
rect 26686 45714 26738 45726
rect 27918 45778 27970 45790
rect 27918 45714 27970 45726
rect 28030 45778 28082 45790
rect 28030 45714 28082 45726
rect 28254 45778 28306 45790
rect 28254 45714 28306 45726
rect 28478 45778 28530 45790
rect 28478 45714 28530 45726
rect 36990 45778 37042 45790
rect 44942 45778 44994 45790
rect 42578 45726 42590 45778
rect 42642 45726 42654 45778
rect 48402 45726 48414 45778
rect 48466 45726 48478 45778
rect 36990 45714 37042 45726
rect 44942 45714 44994 45726
rect 26462 45666 26514 45678
rect 6066 45614 6078 45666
rect 6130 45614 6142 45666
rect 26462 45602 26514 45614
rect 37102 45666 37154 45678
rect 44830 45666 44882 45678
rect 43250 45614 43262 45666
rect 43314 45614 43326 45666
rect 43474 45614 43486 45666
rect 43538 45614 43550 45666
rect 37102 45602 37154 45614
rect 44830 45602 44882 45614
rect 45614 45666 45666 45678
rect 45614 45602 45666 45614
rect 1344 45498 49616 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 49616 45498
rect 1344 45412 49616 45446
rect 9662 45330 9714 45342
rect 30046 45330 30098 45342
rect 28130 45278 28142 45330
rect 28194 45278 28206 45330
rect 9662 45266 9714 45278
rect 30046 45266 30098 45278
rect 30718 45330 30770 45342
rect 41806 45330 41858 45342
rect 36418 45278 36430 45330
rect 36482 45278 36494 45330
rect 30718 45266 30770 45278
rect 41806 45266 41858 45278
rect 25230 45218 25282 45230
rect 3042 45166 3054 45218
rect 3106 45166 3118 45218
rect 8194 45166 8206 45218
rect 8258 45166 8270 45218
rect 21634 45166 21646 45218
rect 21698 45166 21710 45218
rect 25230 45154 25282 45166
rect 29934 45218 29986 45230
rect 29934 45154 29986 45166
rect 31502 45218 31554 45230
rect 31502 45154 31554 45166
rect 32958 45218 33010 45230
rect 32958 45154 33010 45166
rect 35534 45218 35586 45230
rect 41246 45218 41298 45230
rect 38098 45166 38110 45218
rect 38162 45166 38174 45218
rect 35534 45154 35586 45166
rect 41246 45154 41298 45166
rect 41694 45218 41746 45230
rect 41694 45154 41746 45166
rect 42366 45218 42418 45230
rect 48750 45218 48802 45230
rect 45266 45166 45278 45218
rect 45330 45166 45342 45218
rect 42366 45154 42418 45166
rect 48750 45154 48802 45166
rect 25566 45106 25618 45118
rect 2258 45054 2270 45106
rect 2322 45054 2334 45106
rect 8978 45054 8990 45106
rect 9042 45054 9054 45106
rect 23538 45054 23550 45106
rect 23602 45054 23614 45106
rect 25566 45042 25618 45054
rect 26910 45106 26962 45118
rect 28590 45106 28642 45118
rect 27122 45054 27134 45106
rect 27186 45054 27198 45106
rect 26910 45042 26962 45054
rect 28590 45042 28642 45054
rect 28702 45106 28754 45118
rect 28702 45042 28754 45054
rect 28814 45106 28866 45118
rect 30606 45106 30658 45118
rect 30258 45054 30270 45106
rect 30322 45054 30334 45106
rect 28814 45042 28866 45054
rect 30606 45042 30658 45054
rect 30942 45106 30994 45118
rect 30942 45042 30994 45054
rect 31166 45106 31218 45118
rect 33630 45106 33682 45118
rect 32162 45054 32174 45106
rect 32226 45054 32238 45106
rect 33394 45054 33406 45106
rect 33458 45054 33470 45106
rect 31166 45042 31218 45054
rect 33630 45042 33682 45054
rect 33742 45106 33794 45118
rect 33742 45042 33794 45054
rect 33854 45106 33906 45118
rect 36094 45106 36146 45118
rect 49086 45106 49138 45118
rect 35074 45054 35086 45106
rect 35138 45054 35150 45106
rect 37426 45054 37438 45106
rect 37490 45054 37502 45106
rect 47058 45054 47070 45106
rect 47122 45054 47134 45106
rect 33854 45042 33906 45054
rect 36094 45042 36146 45054
rect 49086 45042 49138 45054
rect 18734 44994 18786 45006
rect 5170 44942 5182 44994
rect 5234 44942 5246 44994
rect 6066 44942 6078 44994
rect 6130 44942 6142 44994
rect 9538 44942 9550 44994
rect 9602 44942 9614 44994
rect 18734 44930 18786 44942
rect 27806 44994 27858 45006
rect 35870 44994 35922 45006
rect 32386 44942 32398 44994
rect 32450 44942 32462 44994
rect 35186 44942 35198 44994
rect 35250 44942 35262 44994
rect 27806 44930 27858 44942
rect 35870 44930 35922 44942
rect 37102 44994 37154 45006
rect 41358 44994 41410 45006
rect 40226 44942 40238 44994
rect 40290 44942 40302 44994
rect 37102 44930 37154 44942
rect 41358 44930 41410 44942
rect 42478 44994 42530 45006
rect 42478 44930 42530 44942
rect 9886 44882 9938 44894
rect 9886 44818 9938 44830
rect 41806 44882 41858 44894
rect 41806 44818 41858 44830
rect 42590 44882 42642 44894
rect 42590 44818 42642 44830
rect 1344 44714 49616 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 49616 44714
rect 1344 44628 49616 44662
rect 20414 44546 20466 44558
rect 27358 44546 27410 44558
rect 27010 44494 27022 44546
rect 27074 44494 27086 44546
rect 20414 44482 20466 44494
rect 27358 44482 27410 44494
rect 48078 44546 48130 44558
rect 48078 44482 48130 44494
rect 48414 44546 48466 44558
rect 48850 44494 48862 44546
rect 48914 44543 48926 44546
rect 49298 44543 49310 44546
rect 48914 44497 49310 44543
rect 48914 44494 48926 44497
rect 49298 44494 49310 44497
rect 49362 44494 49374 44546
rect 48414 44482 48466 44494
rect 32510 44434 32562 44446
rect 37214 44434 37266 44446
rect 41134 44434 41186 44446
rect 4610 44382 4622 44434
rect 4674 44382 4686 44434
rect 8978 44382 8990 44434
rect 9042 44382 9054 44434
rect 19282 44382 19294 44434
rect 19346 44382 19358 44434
rect 24546 44382 24558 44434
rect 24610 44382 24622 44434
rect 26674 44382 26686 44434
rect 26738 44382 26750 44434
rect 32050 44382 32062 44434
rect 32114 44382 32126 44434
rect 33394 44382 33406 44434
rect 33458 44382 33470 44434
rect 34738 44382 34750 44434
rect 34802 44382 34814 44434
rect 38322 44382 38334 44434
rect 38386 44382 38398 44434
rect 40450 44382 40462 44434
rect 40514 44382 40526 44434
rect 32510 44370 32562 44382
rect 37214 44370 37266 44382
rect 41134 44370 41186 44382
rect 45614 44434 45666 44446
rect 45614 44370 45666 44382
rect 47182 44434 47234 44446
rect 47182 44370 47234 44382
rect 5742 44322 5794 44334
rect 1810 44270 1822 44322
rect 1874 44270 1886 44322
rect 5742 44258 5794 44270
rect 5854 44322 5906 44334
rect 27582 44322 27634 44334
rect 6178 44270 6190 44322
rect 6242 44270 6254 44322
rect 12226 44270 12238 44322
rect 12290 44270 12302 44322
rect 16482 44270 16494 44322
rect 16546 44270 16558 44322
rect 21970 44270 21982 44322
rect 22034 44270 22046 44322
rect 23874 44270 23886 44322
rect 23938 44270 23950 44322
rect 5854 44258 5906 44270
rect 27582 44258 27634 44270
rect 27918 44322 27970 44334
rect 33518 44322 33570 44334
rect 34190 44322 34242 44334
rect 35086 44322 35138 44334
rect 41022 44322 41074 44334
rect 29138 44270 29150 44322
rect 29202 44270 29214 44322
rect 33954 44270 33966 44322
rect 34018 44270 34030 44322
rect 34850 44270 34862 44322
rect 34914 44270 34926 44322
rect 37538 44270 37550 44322
rect 37602 44270 37614 44322
rect 27918 44258 27970 44270
rect 33518 44258 33570 44270
rect 34190 44258 34242 44270
rect 35086 44258 35138 44270
rect 41022 44258 41074 44270
rect 41358 44322 41410 44334
rect 41358 44258 41410 44270
rect 42478 44322 42530 44334
rect 43038 44322 43090 44334
rect 42690 44270 42702 44322
rect 42754 44270 42766 44322
rect 42478 44258 42530 44270
rect 43038 44258 43090 44270
rect 43262 44322 43314 44334
rect 43822 44322 43874 44334
rect 43586 44270 43598 44322
rect 43650 44270 43662 44322
rect 43262 44258 43314 44270
rect 43822 44258 43874 44270
rect 45838 44322 45890 44334
rect 45838 44258 45890 44270
rect 46062 44322 46114 44334
rect 46062 44258 46114 44270
rect 46510 44322 46562 44334
rect 46510 44258 46562 44270
rect 46622 44322 46674 44334
rect 46622 44258 46674 44270
rect 46734 44322 46786 44334
rect 46734 44258 46786 44270
rect 47406 44322 47458 44334
rect 47406 44258 47458 44270
rect 48190 44322 48242 44334
rect 48190 44258 48242 44270
rect 48526 44322 48578 44334
rect 48526 44258 48578 44270
rect 20302 44210 20354 44222
rect 2482 44158 2494 44210
rect 2546 44158 2558 44210
rect 6066 44158 6078 44210
rect 6130 44158 6142 44210
rect 17154 44158 17166 44210
rect 17218 44158 17230 44210
rect 20302 44146 20354 44158
rect 22318 44210 22370 44222
rect 22318 44146 22370 44158
rect 22990 44210 23042 44222
rect 35870 44210 35922 44222
rect 29922 44158 29934 44210
rect 29986 44158 29998 44210
rect 22990 44146 23042 44158
rect 35870 44146 35922 44158
rect 37102 44210 37154 44222
rect 37102 44146 37154 44158
rect 42142 44210 42194 44222
rect 42142 44146 42194 44158
rect 44270 44210 44322 44222
rect 44270 44146 44322 44158
rect 44830 44210 44882 44222
rect 44830 44146 44882 44158
rect 45054 44210 45106 44222
rect 45054 44146 45106 44158
rect 6638 44098 6690 44110
rect 6638 44034 6690 44046
rect 12686 44098 12738 44110
rect 12686 44034 12738 44046
rect 21646 44098 21698 44110
rect 21646 44034 21698 44046
rect 22206 44098 22258 44110
rect 22206 44034 22258 44046
rect 22430 44098 22482 44110
rect 22430 44034 22482 44046
rect 22542 44098 22594 44110
rect 22542 44034 22594 44046
rect 23102 44098 23154 44110
rect 32398 44098 32450 44110
rect 28242 44046 28254 44098
rect 28306 44046 28318 44098
rect 23102 44034 23154 44046
rect 32398 44034 32450 44046
rect 32958 44098 33010 44110
rect 32958 44034 33010 44046
rect 33406 44098 33458 44110
rect 33406 44034 33458 44046
rect 33742 44098 33794 44110
rect 33742 44034 33794 44046
rect 36206 44098 36258 44110
rect 36206 44034 36258 44046
rect 40910 44098 40962 44110
rect 40910 44034 40962 44046
rect 41246 44098 41298 44110
rect 41246 44034 41298 44046
rect 42254 44098 42306 44110
rect 42254 44034 42306 44046
rect 43150 44098 43202 44110
rect 43150 44034 43202 44046
rect 43934 44098 43986 44110
rect 43934 44034 43986 44046
rect 44046 44098 44098 44110
rect 44046 44034 44098 44046
rect 44942 44098 44994 44110
rect 44942 44034 44994 44046
rect 45502 44098 45554 44110
rect 49198 44098 49250 44110
rect 47730 44046 47742 44098
rect 47794 44046 47806 44098
rect 45502 44034 45554 44046
rect 49198 44034 49250 44046
rect 1344 43930 49616 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 49616 43930
rect 1344 43844 49616 43878
rect 7646 43762 7698 43774
rect 7646 43698 7698 43710
rect 17390 43762 17442 43774
rect 17390 43698 17442 43710
rect 30046 43762 30098 43774
rect 33954 43710 33966 43762
rect 34018 43710 34030 43762
rect 30046 43698 30098 43710
rect 2942 43650 2994 43662
rect 6078 43650 6130 43662
rect 5618 43598 5630 43650
rect 5682 43598 5694 43650
rect 2942 43586 2994 43598
rect 6078 43586 6130 43598
rect 6190 43650 6242 43662
rect 6190 43586 6242 43598
rect 6302 43650 6354 43662
rect 7422 43650 7474 43662
rect 7074 43598 7086 43650
rect 7138 43598 7150 43650
rect 6302 43586 6354 43598
rect 7422 43586 7474 43598
rect 8206 43650 8258 43662
rect 8206 43586 8258 43598
rect 8878 43650 8930 43662
rect 8878 43586 8930 43598
rect 11454 43650 11506 43662
rect 28254 43650 28306 43662
rect 23650 43598 23662 43650
rect 23714 43598 23726 43650
rect 11454 43586 11506 43598
rect 28254 43586 28306 43598
rect 33182 43650 33234 43662
rect 33182 43586 33234 43598
rect 33630 43650 33682 43662
rect 33630 43586 33682 43598
rect 35982 43650 36034 43662
rect 35982 43586 36034 43598
rect 36094 43650 36146 43662
rect 36094 43586 36146 43598
rect 36766 43650 36818 43662
rect 36766 43586 36818 43598
rect 37102 43650 37154 43662
rect 48974 43650 49026 43662
rect 46162 43598 46174 43650
rect 46226 43598 46238 43650
rect 37102 43586 37154 43598
rect 48974 43586 49026 43598
rect 3054 43538 3106 43550
rect 6750 43538 6802 43550
rect 3490 43486 3502 43538
rect 3554 43486 3566 43538
rect 3054 43474 3106 43486
rect 6750 43474 6802 43486
rect 8766 43538 8818 43550
rect 10894 43538 10946 43550
rect 17726 43538 17778 43550
rect 27470 43538 27522 43550
rect 10434 43486 10446 43538
rect 10498 43486 10510 43538
rect 11218 43486 11230 43538
rect 11282 43486 11294 43538
rect 13906 43486 13918 43538
rect 13970 43486 13982 43538
rect 18386 43486 18398 43538
rect 18450 43486 18462 43538
rect 24322 43486 24334 43538
rect 24386 43486 24398 43538
rect 27234 43486 27246 43538
rect 27298 43486 27310 43538
rect 8766 43474 8818 43486
rect 10894 43474 10946 43486
rect 17726 43474 17778 43486
rect 27470 43474 27522 43486
rect 27694 43538 27746 43550
rect 27694 43474 27746 43486
rect 27806 43538 27858 43550
rect 27806 43474 27858 43486
rect 31166 43538 31218 43550
rect 31166 43474 31218 43486
rect 31614 43538 31666 43550
rect 31614 43474 31666 43486
rect 31838 43538 31890 43550
rect 36542 43538 36594 43550
rect 34178 43486 34190 43538
rect 34242 43486 34254 43538
rect 35186 43486 35198 43538
rect 35250 43486 35262 43538
rect 31838 43474 31890 43486
rect 36542 43474 36594 43486
rect 36654 43538 36706 43550
rect 36654 43474 36706 43486
rect 36878 43538 36930 43550
rect 44830 43538 44882 43550
rect 37538 43486 37550 43538
rect 37602 43486 37614 43538
rect 41010 43486 41022 43538
rect 41074 43486 41086 43538
rect 44482 43486 44494 43538
rect 44546 43486 44558 43538
rect 36878 43474 36930 43486
rect 44830 43474 44882 43486
rect 46734 43538 46786 43550
rect 46734 43474 46786 43486
rect 47294 43538 47346 43550
rect 47294 43474 47346 43486
rect 47518 43538 47570 43550
rect 47518 43474 47570 43486
rect 3278 43426 3330 43438
rect 3278 43362 3330 43374
rect 5294 43426 5346 43438
rect 5294 43362 5346 43374
rect 7534 43426 7586 43438
rect 25902 43426 25954 43438
rect 9762 43374 9774 43426
rect 9826 43374 9838 43426
rect 14690 43374 14702 43426
rect 14754 43374 14766 43426
rect 16818 43374 16830 43426
rect 16882 43374 16894 43426
rect 19058 43374 19070 43426
rect 19122 43374 19134 43426
rect 21186 43374 21198 43426
rect 21250 43374 21262 43426
rect 21522 43374 21534 43426
rect 21586 43374 21598 43426
rect 7534 43362 7586 43374
rect 25902 43362 25954 43374
rect 26350 43426 26402 43438
rect 26350 43362 26402 43374
rect 26910 43426 26962 43438
rect 26910 43362 26962 43374
rect 27582 43426 27634 43438
rect 27582 43362 27634 43374
rect 29150 43426 29202 43438
rect 29150 43362 29202 43374
rect 30158 43426 30210 43438
rect 30158 43362 30210 43374
rect 30830 43426 30882 43438
rect 30830 43362 30882 43374
rect 31726 43426 31778 43438
rect 31726 43362 31778 43374
rect 32174 43426 32226 43438
rect 32174 43362 32226 43374
rect 33070 43426 33122 43438
rect 33070 43362 33122 43374
rect 33518 43426 33570 43438
rect 35646 43426 35698 43438
rect 45838 43426 45890 43438
rect 34738 43374 34750 43426
rect 34802 43374 34814 43426
rect 38210 43374 38222 43426
rect 38274 43374 38286 43426
rect 40338 43374 40350 43426
rect 40402 43374 40414 43426
rect 41682 43374 41694 43426
rect 41746 43374 41758 43426
rect 43810 43374 43822 43426
rect 43874 43374 43886 43426
rect 44370 43374 44382 43426
rect 44434 43374 44446 43426
rect 33518 43362 33570 43374
rect 35646 43362 35698 43374
rect 45838 43362 45890 43374
rect 47182 43426 47234 43438
rect 47182 43362 47234 43374
rect 48078 43426 48130 43438
rect 48078 43362 48130 43374
rect 48862 43426 48914 43438
rect 48862 43362 48914 43374
rect 3838 43314 3890 43326
rect 3838 43250 3890 43262
rect 3950 43314 4002 43326
rect 3950 43250 4002 43262
rect 4174 43314 4226 43326
rect 4174 43250 4226 43262
rect 4286 43314 4338 43326
rect 5070 43314 5122 43326
rect 4722 43262 4734 43314
rect 4786 43262 4798 43314
rect 4286 43250 4338 43262
rect 5070 43250 5122 43262
rect 8094 43314 8146 43326
rect 8094 43250 8146 43262
rect 8430 43314 8482 43326
rect 8430 43250 8482 43262
rect 8878 43314 8930 43326
rect 11118 43314 11170 43326
rect 9874 43262 9886 43314
rect 9938 43262 9950 43314
rect 8878 43250 8930 43262
rect 11118 43250 11170 43262
rect 26238 43314 26290 43326
rect 26238 43250 26290 43262
rect 28478 43314 28530 43326
rect 28478 43250 28530 43262
rect 28814 43314 28866 43326
rect 28814 43250 28866 43262
rect 29374 43314 29426 43326
rect 29374 43250 29426 43262
rect 29710 43314 29762 43326
rect 29710 43250 29762 43262
rect 32286 43314 32338 43326
rect 32286 43250 32338 43262
rect 44158 43314 44210 43326
rect 44158 43250 44210 43262
rect 45054 43314 45106 43326
rect 46510 43314 46562 43326
rect 45378 43262 45390 43314
rect 45442 43262 45454 43314
rect 45054 43250 45106 43262
rect 46510 43250 46562 43262
rect 47630 43314 47682 43326
rect 47630 43250 47682 43262
rect 48750 43314 48802 43326
rect 48750 43250 48802 43262
rect 1344 43146 49616 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 49616 43146
rect 1344 43060 49616 43094
rect 6414 42978 6466 42990
rect 19966 42978 20018 42990
rect 11554 42926 11566 42978
rect 11618 42926 11630 42978
rect 6414 42914 6466 42926
rect 19966 42914 20018 42926
rect 27358 42978 27410 42990
rect 27358 42914 27410 42926
rect 29150 42978 29202 42990
rect 29150 42914 29202 42926
rect 37214 42978 37266 42990
rect 43374 42978 43426 42990
rect 37538 42926 37550 42978
rect 37602 42926 37614 42978
rect 37214 42914 37266 42926
rect 43374 42914 43426 42926
rect 44830 42978 44882 42990
rect 44830 42914 44882 42926
rect 44942 42978 44994 42990
rect 44942 42914 44994 42926
rect 45390 42978 45442 42990
rect 45390 42914 45442 42926
rect 45614 42978 45666 42990
rect 45614 42914 45666 42926
rect 18398 42866 18450 42878
rect 2482 42814 2494 42866
rect 2546 42814 2558 42866
rect 4610 42814 4622 42866
rect 4674 42814 4686 42866
rect 6066 42814 6078 42866
rect 6130 42814 6142 42866
rect 9874 42814 9886 42866
rect 9938 42814 9950 42866
rect 18398 42802 18450 42814
rect 19182 42866 19234 42878
rect 19182 42802 19234 42814
rect 23214 42866 23266 42878
rect 29262 42866 29314 42878
rect 36990 42866 37042 42878
rect 42590 42866 42642 42878
rect 26898 42814 26910 42866
rect 26962 42814 26974 42866
rect 28242 42814 28254 42866
rect 28306 42814 28318 42866
rect 30146 42814 30158 42866
rect 30210 42814 30222 42866
rect 32722 42814 32734 42866
rect 32786 42814 32798 42866
rect 35298 42814 35310 42866
rect 35362 42814 35374 42866
rect 42130 42814 42142 42866
rect 42194 42814 42206 42866
rect 23214 42802 23266 42814
rect 29262 42802 29314 42814
rect 36990 42802 37042 42814
rect 42590 42802 42642 42814
rect 44158 42866 44210 42878
rect 47058 42814 47070 42866
rect 47122 42814 47134 42866
rect 49186 42814 49198 42866
rect 49250 42814 49262 42866
rect 44158 42802 44210 42814
rect 6638 42754 6690 42766
rect 10334 42754 10386 42766
rect 12014 42754 12066 42766
rect 1810 42702 1822 42754
rect 1874 42702 1886 42754
rect 7074 42702 7086 42754
rect 7138 42702 7150 42754
rect 10770 42702 10782 42754
rect 10834 42702 10846 42754
rect 6638 42690 6690 42702
rect 10334 42690 10386 42702
rect 12014 42690 12066 42702
rect 12126 42754 12178 42766
rect 16830 42754 16882 42766
rect 12338 42702 12350 42754
rect 12402 42702 12414 42754
rect 12126 42690 12178 42702
rect 16830 42690 16882 42702
rect 17054 42754 17106 42766
rect 27806 42754 27858 42766
rect 21858 42702 21870 42754
rect 21922 42702 21934 42754
rect 22530 42702 22542 42754
rect 22594 42702 22606 42754
rect 22866 42702 22878 42754
rect 22930 42702 22942 42754
rect 24098 42702 24110 42754
rect 24162 42702 24174 42754
rect 17054 42690 17106 42702
rect 27806 42690 27858 42702
rect 27918 42754 27970 42766
rect 27918 42690 27970 42702
rect 28142 42754 28194 42766
rect 31950 42754 32002 42766
rect 28354 42702 28366 42754
rect 28418 42702 28430 42754
rect 29922 42702 29934 42754
rect 29986 42702 29998 42754
rect 30594 42702 30606 42754
rect 30658 42702 30670 42754
rect 28142 42690 28194 42702
rect 31950 42690 32002 42702
rect 32062 42754 32114 42766
rect 32062 42690 32114 42702
rect 32622 42754 32674 42766
rect 32622 42690 32674 42702
rect 33854 42754 33906 42766
rect 35422 42754 35474 42766
rect 34850 42702 34862 42754
rect 34914 42702 34926 42754
rect 35186 42702 35198 42754
rect 35250 42702 35262 42754
rect 33854 42690 33906 42702
rect 35422 42690 35474 42702
rect 35758 42754 35810 42766
rect 35758 42690 35810 42702
rect 38334 42754 38386 42766
rect 38334 42690 38386 42702
rect 38782 42754 38834 42766
rect 42478 42754 42530 42766
rect 39218 42702 39230 42754
rect 39282 42702 39294 42754
rect 38782 42690 38834 42702
rect 42478 42690 42530 42702
rect 42814 42754 42866 42766
rect 42814 42690 42866 42702
rect 42926 42754 42978 42766
rect 46274 42702 46286 42754
rect 46338 42702 46350 42754
rect 42926 42690 42978 42702
rect 10222 42642 10274 42654
rect 7746 42590 7758 42642
rect 7810 42590 7822 42642
rect 10222 42578 10274 42590
rect 14814 42642 14866 42654
rect 14814 42578 14866 42590
rect 15150 42642 15202 42654
rect 20078 42642 20130 42654
rect 16482 42590 16494 42642
rect 16546 42590 16558 42642
rect 15150 42578 15202 42590
rect 20078 42578 20130 42590
rect 22206 42642 22258 42654
rect 22206 42578 22258 42590
rect 23438 42642 23490 42654
rect 27246 42642 27298 42654
rect 24770 42590 24782 42642
rect 24834 42590 24846 42642
rect 23438 42578 23490 42590
rect 27246 42578 27298 42590
rect 30158 42642 30210 42654
rect 30158 42578 30210 42590
rect 31054 42642 31106 42654
rect 31054 42578 31106 42590
rect 33182 42642 33234 42654
rect 33182 42578 33234 42590
rect 34190 42642 34242 42654
rect 43598 42642 43650 42654
rect 40002 42590 40014 42642
rect 40066 42590 40078 42642
rect 34190 42578 34242 42590
rect 43598 42578 43650 42590
rect 44046 42642 44098 42654
rect 44046 42578 44098 42590
rect 45054 42642 45106 42654
rect 45054 42578 45106 42590
rect 18286 42530 18338 42542
rect 18286 42466 18338 42478
rect 19070 42530 19122 42542
rect 19070 42466 19122 42478
rect 21646 42530 21698 42542
rect 21646 42466 21698 42478
rect 22094 42530 22146 42542
rect 22094 42466 22146 42478
rect 22318 42530 22370 42542
rect 22318 42466 22370 42478
rect 23102 42530 23154 42542
rect 23102 42466 23154 42478
rect 23326 42530 23378 42542
rect 23326 42466 23378 42478
rect 30382 42530 30434 42542
rect 30382 42466 30434 42478
rect 31166 42530 31218 42542
rect 31166 42466 31218 42478
rect 31614 42530 31666 42542
rect 31614 42466 31666 42478
rect 31726 42530 31778 42542
rect 31726 42466 31778 42478
rect 31838 42530 31890 42542
rect 31838 42466 31890 42478
rect 32734 42530 32786 42542
rect 32734 42466 32786 42478
rect 32958 42530 33010 42542
rect 32958 42466 33010 42478
rect 33742 42530 33794 42542
rect 33742 42466 33794 42478
rect 34414 42530 34466 42542
rect 34414 42466 34466 42478
rect 34526 42530 34578 42542
rect 34526 42466 34578 42478
rect 34638 42530 34690 42542
rect 34638 42466 34690 42478
rect 35646 42530 35698 42542
rect 35646 42466 35698 42478
rect 36430 42530 36482 42542
rect 36430 42466 36482 42478
rect 38446 42530 38498 42542
rect 38446 42466 38498 42478
rect 38558 42530 38610 42542
rect 38558 42466 38610 42478
rect 38670 42530 38722 42542
rect 38670 42466 38722 42478
rect 43486 42530 43538 42542
rect 43486 42466 43538 42478
rect 1344 42362 49616 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 49616 42362
rect 1344 42276 49616 42310
rect 7982 42194 8034 42206
rect 22318 42194 22370 42206
rect 17938 42142 17950 42194
rect 18002 42142 18014 42194
rect 7982 42130 8034 42142
rect 22318 42130 22370 42142
rect 24670 42194 24722 42206
rect 24670 42130 24722 42142
rect 32398 42194 32450 42206
rect 39454 42194 39506 42206
rect 38546 42142 38558 42194
rect 38610 42142 38622 42194
rect 32398 42130 32450 42142
rect 39454 42130 39506 42142
rect 39678 42194 39730 42206
rect 39678 42130 39730 42142
rect 47182 42194 47234 42206
rect 47182 42130 47234 42142
rect 13806 42082 13858 42094
rect 13806 42018 13858 42030
rect 16830 42082 16882 42094
rect 39902 42082 39954 42094
rect 18946 42030 18958 42082
rect 19010 42030 19022 42082
rect 31490 42030 31502 42082
rect 31554 42030 31566 42082
rect 34402 42030 34414 42082
rect 34466 42030 34478 42082
rect 16830 42018 16882 42030
rect 39902 42018 39954 42030
rect 42702 42082 42754 42094
rect 42702 42018 42754 42030
rect 43262 42082 43314 42094
rect 43262 42018 43314 42030
rect 48862 42082 48914 42094
rect 48862 42018 48914 42030
rect 8206 41970 8258 41982
rect 6626 41918 6638 41970
rect 6690 41918 6702 41970
rect 8206 41906 8258 41918
rect 8654 41970 8706 41982
rect 13470 41970 13522 41982
rect 16718 41970 16770 41982
rect 23102 41970 23154 41982
rect 9986 41918 9998 41970
rect 10050 41918 10062 41970
rect 16370 41918 16382 41970
rect 16434 41918 16446 41970
rect 19170 41918 19182 41970
rect 19234 41918 19246 41970
rect 8654 41906 8706 41918
rect 13470 41906 13522 41918
rect 16718 41906 16770 41918
rect 23102 41906 23154 41918
rect 24558 41970 24610 41982
rect 32510 41970 32562 41982
rect 25218 41918 25230 41970
rect 25282 41918 25294 41970
rect 30818 41918 30830 41970
rect 30882 41918 30894 41970
rect 31378 41918 31390 41970
rect 31442 41918 31454 41970
rect 24558 41906 24610 41918
rect 32510 41906 32562 41918
rect 33070 41970 33122 41982
rect 38894 41970 38946 41982
rect 37426 41918 37438 41970
rect 37490 41918 37502 41970
rect 38098 41918 38110 41970
rect 38162 41918 38174 41970
rect 33070 41906 33122 41918
rect 38894 41906 38946 41918
rect 39342 41970 39394 41982
rect 39342 41906 39394 41918
rect 40350 41970 40402 41982
rect 40350 41906 40402 41918
rect 41694 41970 41746 41982
rect 41694 41906 41746 41918
rect 43038 41970 43090 41982
rect 43038 41906 43090 41918
rect 43598 41970 43650 41982
rect 43598 41906 43650 41918
rect 44494 41970 44546 41982
rect 44494 41906 44546 41918
rect 44718 41970 44770 41982
rect 44718 41906 44770 41918
rect 45726 41970 45778 41982
rect 45726 41906 45778 41918
rect 47182 41970 47234 41982
rect 47182 41906 47234 41918
rect 47518 41970 47570 41982
rect 47518 41906 47570 41918
rect 49198 41970 49250 41982
rect 49198 41906 49250 41918
rect 17390 41858 17442 41870
rect 2258 41806 2270 41858
rect 2322 41806 2334 41858
rect 7858 41806 7870 41858
rect 7922 41806 7934 41858
rect 10658 41806 10670 41858
rect 10722 41806 10734 41858
rect 12786 41806 12798 41858
rect 12850 41806 12862 41858
rect 17390 41794 17442 41806
rect 18510 41858 18562 41870
rect 18510 41794 18562 41806
rect 20078 41858 20130 41870
rect 20078 41794 20130 41806
rect 22542 41858 22594 41870
rect 22542 41794 22594 41806
rect 23550 41858 23602 41870
rect 23550 41794 23602 41806
rect 24334 41858 24386 41870
rect 33518 41858 33570 41870
rect 27234 41806 27246 41858
rect 27298 41806 27310 41858
rect 31490 41806 31502 41858
rect 31554 41806 31566 41858
rect 24334 41794 24386 41806
rect 33518 41794 33570 41806
rect 34750 41858 34802 41870
rect 39566 41858 39618 41870
rect 35186 41806 35198 41858
rect 35250 41806 35262 41858
rect 34750 41794 34802 41806
rect 39566 41794 39618 41806
rect 40238 41858 40290 41870
rect 40238 41794 40290 41806
rect 41470 41858 41522 41870
rect 41470 41794 41522 41806
rect 41806 41858 41858 41870
rect 41806 41794 41858 41806
rect 43486 41858 43538 41870
rect 43486 41794 43538 41806
rect 44942 41858 44994 41870
rect 44942 41794 44994 41806
rect 45278 41858 45330 41870
rect 45278 41794 45330 41806
rect 46734 41858 46786 41870
rect 46734 41794 46786 41806
rect 48190 41858 48242 41870
rect 48190 41794 48242 41806
rect 17614 41746 17666 41758
rect 17614 41682 17666 41694
rect 18622 41746 18674 41758
rect 18622 41682 18674 41694
rect 19966 41746 20018 41758
rect 19966 41682 20018 41694
rect 22654 41746 22706 41758
rect 32398 41746 32450 41758
rect 22866 41694 22878 41746
rect 22930 41743 22942 41746
rect 23426 41743 23438 41746
rect 22930 41697 23438 41743
rect 22930 41694 22942 41697
rect 23426 41694 23438 41697
rect 23490 41694 23502 41746
rect 22654 41682 22706 41694
rect 32398 41682 32450 41694
rect 33294 41746 33346 41758
rect 33294 41682 33346 41694
rect 33966 41746 34018 41758
rect 33966 41682 34018 41694
rect 42254 41746 42306 41758
rect 42254 41682 42306 41694
rect 42366 41746 42418 41758
rect 42366 41682 42418 41694
rect 42590 41746 42642 41758
rect 42590 41682 42642 41694
rect 43822 41746 43874 41758
rect 43822 41682 43874 41694
rect 44270 41746 44322 41758
rect 44270 41682 44322 41694
rect 45502 41746 45554 41758
rect 45502 41682 45554 41694
rect 45950 41746 46002 41758
rect 45950 41682 46002 41694
rect 46398 41746 46450 41758
rect 46398 41682 46450 41694
rect 47294 41746 47346 41758
rect 47294 41682 47346 41694
rect 1344 41578 49616 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 49616 41578
rect 1344 41492 49616 41526
rect 36206 41410 36258 41422
rect 30706 41358 30718 41410
rect 30770 41358 30782 41410
rect 36206 41346 36258 41358
rect 37102 41410 37154 41422
rect 37102 41346 37154 41358
rect 6414 41298 6466 41310
rect 12910 41298 12962 41310
rect 17726 41298 17778 41310
rect 20638 41298 20690 41310
rect 28478 41298 28530 41310
rect 44046 41298 44098 41310
rect 4610 41246 4622 41298
rect 4674 41246 4686 41298
rect 9538 41246 9550 41298
rect 9602 41246 9614 41298
rect 14242 41246 14254 41298
rect 14306 41246 14318 41298
rect 16370 41246 16382 41298
rect 16434 41246 16446 41298
rect 20066 41246 20078 41298
rect 20130 41246 20142 41298
rect 21298 41246 21310 41298
rect 21362 41246 21374 41298
rect 23426 41246 23438 41298
rect 23490 41246 23502 41298
rect 25554 41246 25566 41298
rect 25618 41246 25630 41298
rect 27682 41246 27694 41298
rect 27746 41246 27758 41298
rect 30370 41246 30382 41298
rect 30434 41246 30446 41298
rect 33954 41246 33966 41298
rect 34018 41246 34030 41298
rect 38546 41246 38558 41298
rect 38610 41246 38622 41298
rect 47058 41246 47070 41298
rect 47122 41246 47134 41298
rect 49186 41246 49198 41298
rect 49250 41246 49262 41298
rect 6414 41234 6466 41246
rect 12910 41234 12962 41246
rect 17726 41234 17778 41246
rect 20638 41234 20690 41246
rect 28478 41234 28530 41246
rect 44046 41234 44098 41246
rect 6750 41186 6802 41198
rect 17614 41186 17666 41198
rect 1810 41134 1822 41186
rect 1874 41134 1886 41186
rect 6962 41134 6974 41186
rect 7026 41134 7038 41186
rect 12450 41134 12462 41186
rect 12514 41134 12526 41186
rect 13570 41134 13582 41186
rect 13634 41134 13646 41186
rect 17042 41134 17054 41186
rect 17106 41134 17118 41186
rect 6750 41122 6802 41134
rect 17614 41122 17666 41134
rect 18174 41186 18226 41198
rect 18174 41122 18226 41134
rect 18846 41186 18898 41198
rect 29374 41186 29426 41198
rect 19506 41134 19518 41186
rect 19570 41134 19582 41186
rect 20178 41134 20190 41186
rect 20242 41134 20254 41186
rect 24098 41134 24110 41186
rect 24162 41134 24174 41186
rect 24770 41134 24782 41186
rect 24834 41134 24846 41186
rect 29138 41134 29150 41186
rect 29202 41134 29214 41186
rect 18846 41122 18898 41134
rect 29374 41122 29426 41134
rect 29486 41186 29538 41198
rect 35198 41186 35250 41198
rect 31490 41134 31502 41186
rect 31554 41134 31566 41186
rect 32274 41134 32286 41186
rect 32338 41134 32350 41186
rect 33618 41134 33630 41186
rect 33682 41134 33694 41186
rect 29486 41122 29538 41134
rect 35198 41122 35250 41134
rect 35534 41186 35586 41198
rect 44830 41186 44882 41198
rect 42130 41134 42142 41186
rect 42194 41134 42206 41186
rect 44258 41134 44270 41186
rect 44322 41134 44334 41186
rect 35534 41122 35586 41134
rect 44830 41122 44882 41134
rect 45390 41186 45442 41198
rect 46386 41134 46398 41186
rect 46450 41134 46462 41186
rect 45390 41122 45442 41134
rect 18734 41074 18786 41086
rect 2482 41022 2494 41074
rect 2546 41022 2558 41074
rect 6514 41022 6526 41074
rect 6578 41022 6590 41074
rect 8306 41022 8318 41074
rect 8370 41022 8382 41074
rect 11666 41022 11678 41074
rect 11730 41022 11742 41074
rect 18498 41022 18510 41074
rect 18562 41022 18574 41074
rect 18734 41010 18786 41022
rect 19742 41074 19794 41086
rect 19742 41010 19794 41022
rect 20526 41074 20578 41086
rect 20526 41010 20578 41022
rect 28590 41074 28642 41086
rect 28590 41010 28642 41022
rect 36318 41074 36370 41086
rect 36318 41010 36370 41022
rect 36990 41074 37042 41086
rect 43934 41074 43986 41086
rect 37650 41022 37662 41074
rect 37714 41022 37726 41074
rect 36990 41010 37042 41022
rect 43934 41010 43986 41022
rect 5742 40962 5794 40974
rect 7422 40962 7474 40974
rect 6066 40910 6078 40962
rect 6130 40910 6142 40962
rect 5742 40898 5794 40910
rect 7422 40898 7474 40910
rect 7646 40962 7698 40974
rect 8654 40962 8706 40974
rect 7970 40910 7982 40962
rect 8034 40910 8046 40962
rect 7646 40898 7698 40910
rect 8654 40898 8706 40910
rect 9102 40962 9154 40974
rect 9102 40898 9154 40910
rect 12798 40962 12850 40974
rect 12798 40898 12850 40910
rect 17950 40962 18002 40974
rect 17950 40898 18002 40910
rect 19966 40962 20018 40974
rect 19966 40898 20018 40910
rect 28142 40962 28194 40974
rect 35310 40962 35362 40974
rect 29922 40910 29934 40962
rect 29986 40910 29998 40962
rect 28142 40898 28194 40910
rect 35310 40898 35362 40910
rect 35422 40962 35474 40974
rect 35422 40898 35474 40910
rect 35646 40962 35698 40974
rect 35646 40898 35698 40910
rect 36206 40962 36258 40974
rect 36206 40898 36258 40910
rect 37998 40962 38050 40974
rect 37998 40898 38050 40910
rect 44718 40962 44770 40974
rect 44718 40898 44770 40910
rect 45054 40962 45106 40974
rect 45054 40898 45106 40910
rect 45278 40962 45330 40974
rect 45278 40898 45330 40910
rect 45950 40962 46002 40974
rect 45950 40898 46002 40910
rect 1344 40794 49616 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 49616 40794
rect 1344 40708 49616 40742
rect 17502 40626 17554 40638
rect 6626 40574 6638 40626
rect 6690 40574 6702 40626
rect 10658 40574 10670 40626
rect 10722 40574 10734 40626
rect 17502 40562 17554 40574
rect 19854 40626 19906 40638
rect 19854 40562 19906 40574
rect 20078 40626 20130 40638
rect 20078 40562 20130 40574
rect 20974 40626 21026 40638
rect 20974 40562 21026 40574
rect 21534 40626 21586 40638
rect 21534 40562 21586 40574
rect 22990 40626 23042 40638
rect 22990 40562 23042 40574
rect 23102 40626 23154 40638
rect 23102 40562 23154 40574
rect 23214 40626 23266 40638
rect 23998 40626 24050 40638
rect 23650 40574 23662 40626
rect 23714 40574 23726 40626
rect 23214 40562 23266 40574
rect 23998 40562 24050 40574
rect 25902 40626 25954 40638
rect 25902 40562 25954 40574
rect 27470 40626 27522 40638
rect 27470 40562 27522 40574
rect 27582 40626 27634 40638
rect 27582 40562 27634 40574
rect 27694 40626 27746 40638
rect 27694 40562 27746 40574
rect 33630 40626 33682 40638
rect 33630 40562 33682 40574
rect 34526 40626 34578 40638
rect 34526 40562 34578 40574
rect 39006 40626 39058 40638
rect 39006 40562 39058 40574
rect 39902 40626 39954 40638
rect 39902 40562 39954 40574
rect 40350 40626 40402 40638
rect 40350 40562 40402 40574
rect 41022 40626 41074 40638
rect 41022 40562 41074 40574
rect 42366 40626 42418 40638
rect 42366 40562 42418 40574
rect 48974 40626 49026 40638
rect 48974 40562 49026 40574
rect 2718 40514 2770 40526
rect 2718 40450 2770 40462
rect 7758 40514 7810 40526
rect 7758 40450 7810 40462
rect 8766 40514 8818 40526
rect 8766 40450 8818 40462
rect 10894 40514 10946 40526
rect 22094 40514 22146 40526
rect 13570 40462 13582 40514
rect 13634 40462 13646 40514
rect 10894 40450 10946 40462
rect 22094 40450 22146 40462
rect 22654 40514 22706 40526
rect 22654 40450 22706 40462
rect 25454 40514 25506 40526
rect 39454 40514 39506 40526
rect 29810 40462 29822 40514
rect 29874 40462 29886 40514
rect 25454 40450 25506 40462
rect 39454 40450 39506 40462
rect 41806 40514 41858 40526
rect 41806 40450 41858 40462
rect 3726 40402 3778 40414
rect 5070 40402 5122 40414
rect 4610 40350 4622 40402
rect 4674 40350 4686 40402
rect 3726 40338 3778 40350
rect 5070 40338 5122 40350
rect 5406 40402 5458 40414
rect 5406 40338 5458 40350
rect 5742 40402 5794 40414
rect 5742 40338 5794 40350
rect 6302 40402 6354 40414
rect 6302 40338 6354 40350
rect 7646 40402 7698 40414
rect 7646 40338 7698 40350
rect 8094 40402 8146 40414
rect 10446 40402 10498 40414
rect 10322 40350 10334 40402
rect 10386 40350 10398 40402
rect 8094 40338 8146 40350
rect 10446 40338 10498 40350
rect 10558 40402 10610 40414
rect 17726 40402 17778 40414
rect 20526 40402 20578 40414
rect 16594 40350 16606 40402
rect 16658 40350 16670 40402
rect 18162 40350 18174 40402
rect 18226 40350 18238 40402
rect 18386 40350 18398 40402
rect 18450 40350 18462 40402
rect 19618 40350 19630 40402
rect 19682 40350 19694 40402
rect 20290 40350 20302 40402
rect 20354 40350 20366 40402
rect 10558 40338 10610 40350
rect 17726 40338 17778 40350
rect 20526 40338 20578 40350
rect 21198 40402 21250 40414
rect 21198 40338 21250 40350
rect 21982 40402 22034 40414
rect 21982 40338 22034 40350
rect 22878 40402 22930 40414
rect 22878 40338 22930 40350
rect 24446 40402 24498 40414
rect 24446 40338 24498 40350
rect 25678 40402 25730 40414
rect 27358 40402 27410 40414
rect 32958 40402 33010 40414
rect 26114 40350 26126 40402
rect 26178 40350 26190 40402
rect 27906 40350 27918 40402
rect 27970 40350 27982 40402
rect 30146 40350 30158 40402
rect 30210 40350 30222 40402
rect 31042 40350 31054 40402
rect 31106 40350 31118 40402
rect 32162 40350 32174 40402
rect 32226 40350 32238 40402
rect 25678 40338 25730 40350
rect 27358 40338 27410 40350
rect 32958 40338 33010 40350
rect 33406 40402 33458 40414
rect 33406 40338 33458 40350
rect 34414 40402 34466 40414
rect 34414 40338 34466 40350
rect 34638 40402 34690 40414
rect 38894 40402 38946 40414
rect 37314 40350 37326 40402
rect 37378 40350 37390 40402
rect 38098 40350 38110 40402
rect 38162 40350 38174 40402
rect 34638 40338 34690 40350
rect 38894 40338 38946 40350
rect 39230 40402 39282 40414
rect 42914 40350 42926 40402
rect 42978 40350 42990 40402
rect 46386 40350 46398 40402
rect 46450 40350 46462 40402
rect 39230 40338 39282 40350
rect 2942 40290 2994 40302
rect 5294 40290 5346 40302
rect 2594 40238 2606 40290
rect 2658 40238 2670 40290
rect 4498 40238 4510 40290
rect 4562 40238 4574 40290
rect 2942 40226 2994 40238
rect 5294 40226 5346 40238
rect 6078 40290 6130 40302
rect 6078 40226 6130 40238
rect 7982 40290 8034 40302
rect 19966 40290 20018 40302
rect 18050 40238 18062 40290
rect 18114 40238 18126 40290
rect 7982 40226 8034 40238
rect 19966 40226 20018 40238
rect 21086 40290 21138 40302
rect 21086 40226 21138 40238
rect 21646 40290 21698 40302
rect 21646 40226 21698 40238
rect 25790 40290 25842 40302
rect 25790 40226 25842 40238
rect 26686 40290 26738 40302
rect 26686 40226 26738 40238
rect 28478 40290 28530 40302
rect 28478 40226 28530 40238
rect 33518 40290 33570 40302
rect 33518 40226 33570 40238
rect 33966 40290 34018 40302
rect 33966 40226 34018 40238
rect 34190 40290 34242 40302
rect 39118 40290 39170 40302
rect 35186 40238 35198 40290
rect 35250 40238 35262 40290
rect 34190 40226 34242 40238
rect 39118 40226 39170 40238
rect 39790 40290 39842 40302
rect 39790 40226 39842 40238
rect 41470 40290 41522 40302
rect 41470 40226 41522 40238
rect 42590 40290 42642 40302
rect 48962 40238 48974 40290
rect 49026 40238 49038 40290
rect 42590 40226 42642 40238
rect 8542 40178 8594 40190
rect 8542 40114 8594 40126
rect 8878 40178 8930 40190
rect 8878 40114 8930 40126
rect 24558 40178 24610 40190
rect 24558 40114 24610 40126
rect 26798 40178 26850 40190
rect 26798 40114 26850 40126
rect 28590 40178 28642 40190
rect 41918 40178 41970 40190
rect 31826 40126 31838 40178
rect 31890 40126 31902 40178
rect 28590 40114 28642 40126
rect 41918 40114 41970 40126
rect 42254 40178 42306 40190
rect 42254 40114 42306 40126
rect 48750 40178 48802 40190
rect 48750 40114 48802 40126
rect 1344 40010 49616 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 49616 40010
rect 1344 39924 49616 39958
rect 36430 39842 36482 39854
rect 8978 39790 8990 39842
rect 9042 39790 9054 39842
rect 13682 39790 13694 39842
rect 13746 39790 13758 39842
rect 46498 39790 46510 39842
rect 46562 39790 46574 39842
rect 36430 39778 36482 39790
rect 18734 39730 18786 39742
rect 21646 39730 21698 39742
rect 43374 39730 43426 39742
rect 5058 39678 5070 39730
rect 5122 39678 5134 39730
rect 9314 39678 9326 39730
rect 9378 39678 9390 39730
rect 19618 39678 19630 39730
rect 19682 39678 19694 39730
rect 22418 39678 22430 39730
rect 22482 39678 22494 39730
rect 24546 39678 24558 39730
rect 24610 39678 24622 39730
rect 25666 39678 25678 39730
rect 25730 39678 25742 39730
rect 27794 39678 27806 39730
rect 27858 39678 27870 39730
rect 42690 39678 42702 39730
rect 42754 39678 42766 39730
rect 18734 39666 18786 39678
rect 21646 39666 21698 39678
rect 43374 39666 43426 39678
rect 44158 39730 44210 39742
rect 44158 39666 44210 39678
rect 47742 39730 47794 39742
rect 48738 39678 48750 39730
rect 48802 39678 48814 39730
rect 47742 39666 47794 39678
rect 5854 39618 5906 39630
rect 2146 39566 2158 39618
rect 2210 39566 2222 39618
rect 5618 39566 5630 39618
rect 5682 39566 5694 39618
rect 5854 39554 5906 39566
rect 6078 39618 6130 39630
rect 7534 39618 7586 39630
rect 7298 39566 7310 39618
rect 7362 39566 7374 39618
rect 6078 39554 6130 39566
rect 7534 39554 7586 39566
rect 7646 39618 7698 39630
rect 7646 39554 7698 39566
rect 7758 39618 7810 39630
rect 14030 39618 14082 39630
rect 8194 39566 8206 39618
rect 8258 39566 8270 39618
rect 12226 39566 12238 39618
rect 12290 39566 12302 39618
rect 12674 39566 12686 39618
rect 12738 39566 12750 39618
rect 7758 39554 7810 39566
rect 14030 39554 14082 39566
rect 14254 39618 14306 39630
rect 14254 39554 14306 39566
rect 15038 39618 15090 39630
rect 15038 39554 15090 39566
rect 16382 39618 16434 39630
rect 16382 39554 16434 39566
rect 16494 39618 16546 39630
rect 16494 39554 16546 39566
rect 16942 39618 16994 39630
rect 16942 39554 16994 39566
rect 19182 39618 19234 39630
rect 19742 39618 19794 39630
rect 19506 39566 19518 39618
rect 19570 39566 19582 39618
rect 19182 39554 19234 39566
rect 19742 39554 19794 39566
rect 19966 39618 20018 39630
rect 20526 39618 20578 39630
rect 20178 39566 20190 39618
rect 20242 39566 20254 39618
rect 19966 39554 20018 39566
rect 20526 39554 20578 39566
rect 21422 39618 21474 39630
rect 21422 39554 21474 39566
rect 21870 39618 21922 39630
rect 34862 39618 34914 39630
rect 25218 39566 25230 39618
rect 25282 39566 25294 39618
rect 28578 39566 28590 39618
rect 28642 39566 28654 39618
rect 34402 39566 34414 39618
rect 34466 39566 34478 39618
rect 21870 39554 21922 39566
rect 34862 39554 34914 39566
rect 35310 39618 35362 39630
rect 35310 39554 35362 39566
rect 35422 39618 35474 39630
rect 37214 39618 37266 39630
rect 36978 39566 36990 39618
rect 37042 39566 37054 39618
rect 35422 39554 35474 39566
rect 37214 39554 37266 39566
rect 37438 39618 37490 39630
rect 37998 39618 38050 39630
rect 37650 39566 37662 39618
rect 37714 39566 37726 39618
rect 37438 39554 37490 39566
rect 37998 39554 38050 39566
rect 38670 39618 38722 39630
rect 43150 39618 43202 39630
rect 39778 39566 39790 39618
rect 39842 39566 39854 39618
rect 38670 39554 38722 39566
rect 43150 39554 43202 39566
rect 43486 39618 43538 39630
rect 45054 39618 45106 39630
rect 43698 39566 43710 39618
rect 43762 39566 43774 39618
rect 43486 39554 43538 39566
rect 45054 39554 45106 39566
rect 45278 39618 45330 39630
rect 45278 39554 45330 39566
rect 45390 39618 45442 39630
rect 47070 39618 47122 39630
rect 45714 39566 45726 39618
rect 45778 39566 45790 39618
rect 45390 39554 45442 39566
rect 47070 39554 47122 39566
rect 47182 39618 47234 39630
rect 47182 39554 47234 39566
rect 47966 39618 48018 39630
rect 47966 39554 48018 39566
rect 48190 39618 48242 39630
rect 48190 39554 48242 39566
rect 8430 39506 8482 39518
rect 2930 39454 2942 39506
rect 2994 39454 3006 39506
rect 8430 39442 8482 39454
rect 8542 39506 8594 39518
rect 14926 39506 14978 39518
rect 11442 39454 11454 39506
rect 11506 39454 11518 39506
rect 8542 39442 8594 39454
rect 14926 39442 14978 39454
rect 17726 39506 17778 39518
rect 17726 39442 17778 39454
rect 18622 39506 18674 39518
rect 18622 39442 18674 39454
rect 19070 39506 19122 39518
rect 19070 39442 19122 39454
rect 20638 39506 20690 39518
rect 20638 39442 20690 39454
rect 21758 39506 21810 39518
rect 36318 39506 36370 39518
rect 29362 39454 29374 39506
rect 29426 39454 29438 39506
rect 21758 39442 21810 39454
rect 36318 39442 36370 39454
rect 37326 39506 37378 39518
rect 43262 39506 43314 39518
rect 40562 39454 40574 39506
rect 40626 39454 40638 39506
rect 37326 39442 37378 39454
rect 43262 39442 43314 39454
rect 44830 39506 44882 39518
rect 44830 39442 44882 39454
rect 46958 39506 47010 39518
rect 46958 39442 47010 39454
rect 47630 39506 47682 39518
rect 47630 39442 47682 39454
rect 48862 39506 48914 39518
rect 48862 39442 48914 39454
rect 49086 39506 49138 39518
rect 49086 39442 49138 39454
rect 5742 39394 5794 39406
rect 5742 39330 5794 39342
rect 6862 39394 6914 39406
rect 6862 39330 6914 39342
rect 12910 39394 12962 39406
rect 12910 39330 12962 39342
rect 15150 39394 15202 39406
rect 15934 39394 15986 39406
rect 15586 39342 15598 39394
rect 15650 39342 15662 39394
rect 15150 39330 15202 39342
rect 15934 39330 15986 39342
rect 16718 39394 16770 39406
rect 16718 39330 16770 39342
rect 17502 39394 17554 39406
rect 17502 39330 17554 39342
rect 17614 39394 17666 39406
rect 17614 39330 17666 39342
rect 20862 39394 20914 39406
rect 20862 39330 20914 39342
rect 21534 39394 21586 39406
rect 21534 39330 21586 39342
rect 35534 39394 35586 39406
rect 35534 39330 35586 39342
rect 35646 39394 35698 39406
rect 35646 39330 35698 39342
rect 35758 39394 35810 39406
rect 39454 39394 39506 39406
rect 38322 39342 38334 39394
rect 38386 39342 38398 39394
rect 38994 39342 39006 39394
rect 39058 39342 39070 39394
rect 35758 39330 35810 39342
rect 39454 39330 39506 39342
rect 44718 39394 44770 39406
rect 44718 39330 44770 39342
rect 46286 39394 46338 39406
rect 46286 39330 46338 39342
rect 1344 39226 49616 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 49616 39226
rect 1344 39140 49616 39174
rect 26574 39058 26626 39070
rect 22978 39006 22990 39058
rect 23042 39006 23054 39058
rect 24658 39006 24670 39058
rect 24722 39006 24734 39058
rect 26574 38994 26626 39006
rect 26686 39058 26738 39070
rect 26686 38994 26738 39006
rect 26910 39058 26962 39070
rect 40350 39058 40402 39070
rect 27346 39006 27358 39058
rect 27410 39006 27422 39058
rect 28466 39006 28478 39058
rect 28530 39006 28542 39058
rect 32162 39006 32174 39058
rect 32226 39006 32238 39058
rect 26910 38994 26962 39006
rect 40350 38994 40402 39006
rect 41022 39058 41074 39070
rect 41022 38994 41074 39006
rect 41134 39058 41186 39070
rect 41134 38994 41186 39006
rect 41246 39058 41298 39070
rect 41246 38994 41298 39006
rect 41358 39058 41410 39070
rect 41358 38994 41410 39006
rect 42478 39058 42530 39070
rect 42478 38994 42530 39006
rect 43598 39058 43650 39070
rect 43598 38994 43650 39006
rect 44270 39058 44322 39070
rect 44270 38994 44322 39006
rect 7646 38946 7698 38958
rect 7646 38882 7698 38894
rect 8878 38946 8930 38958
rect 8878 38882 8930 38894
rect 10110 38946 10162 38958
rect 22654 38946 22706 38958
rect 13234 38894 13246 38946
rect 13298 38894 13310 38946
rect 10110 38882 10162 38894
rect 22654 38882 22706 38894
rect 23774 38946 23826 38958
rect 23774 38882 23826 38894
rect 25790 38946 25842 38958
rect 25790 38882 25842 38894
rect 26350 38946 26402 38958
rect 33070 38946 33122 38958
rect 41582 38946 41634 38958
rect 29922 38894 29934 38946
rect 29986 38894 29998 38946
rect 35410 38894 35422 38946
rect 35474 38894 35486 38946
rect 36306 38894 36318 38946
rect 36370 38894 36382 38946
rect 26350 38882 26402 38894
rect 33070 38882 33122 38894
rect 41582 38882 41634 38894
rect 45166 38946 45218 38958
rect 45166 38882 45218 38894
rect 47630 38946 47682 38958
rect 48738 38894 48750 38946
rect 48802 38894 48814 38946
rect 47630 38882 47682 38894
rect 6862 38834 6914 38846
rect 1810 38782 1822 38834
rect 1874 38782 1886 38834
rect 5954 38782 5966 38834
rect 6018 38782 6030 38834
rect 6862 38770 6914 38782
rect 7086 38834 7138 38846
rect 7086 38770 7138 38782
rect 7534 38834 7586 38846
rect 7534 38770 7586 38782
rect 8542 38834 8594 38846
rect 9774 38834 9826 38846
rect 18062 38834 18114 38846
rect 9538 38782 9550 38834
rect 9602 38782 9614 38834
rect 12450 38782 12462 38834
rect 12514 38782 12526 38834
rect 16370 38782 16382 38834
rect 16434 38782 16446 38834
rect 8542 38770 8594 38782
rect 9774 38770 9826 38782
rect 18062 38770 18114 38782
rect 20750 38834 20802 38846
rect 20750 38770 20802 38782
rect 20974 38834 21026 38846
rect 20974 38770 21026 38782
rect 21198 38834 21250 38846
rect 21198 38770 21250 38782
rect 21646 38834 21698 38846
rect 21646 38770 21698 38782
rect 21758 38834 21810 38846
rect 21758 38770 21810 38782
rect 21982 38834 22034 38846
rect 23326 38834 23378 38846
rect 22194 38782 22206 38834
rect 22258 38782 22270 38834
rect 21982 38770 22034 38782
rect 23326 38770 23378 38782
rect 23886 38834 23938 38846
rect 23886 38770 23938 38782
rect 24334 38834 24386 38846
rect 24334 38770 24386 38782
rect 25342 38834 25394 38846
rect 25342 38770 25394 38782
rect 26798 38834 26850 38846
rect 26798 38770 26850 38782
rect 27694 38834 27746 38846
rect 27694 38770 27746 38782
rect 28142 38834 28194 38846
rect 43486 38834 43538 38846
rect 44158 38834 44210 38846
rect 28690 38782 28702 38834
rect 28754 38782 28766 38834
rect 29250 38782 29262 38834
rect 29314 38782 29326 38834
rect 34850 38782 34862 38834
rect 34914 38782 34926 38834
rect 36642 38782 36654 38834
rect 36706 38782 36718 38834
rect 38098 38782 38110 38834
rect 38162 38782 38174 38834
rect 38770 38782 38782 38834
rect 38834 38782 38846 38834
rect 43922 38782 43934 38834
rect 43986 38782 43998 38834
rect 28142 38770 28194 38782
rect 43486 38770 43538 38782
rect 44158 38770 44210 38782
rect 44382 38834 44434 38846
rect 45838 38834 45890 38846
rect 48078 38834 48130 38846
rect 44594 38782 44606 38834
rect 44658 38782 44670 38834
rect 46274 38782 46286 38834
rect 46338 38782 46350 38834
rect 47058 38782 47070 38834
rect 47122 38782 47134 38834
rect 47394 38782 47406 38834
rect 47458 38782 47470 38834
rect 44382 38770 44434 38782
rect 45838 38770 45890 38782
rect 48078 38770 48130 38782
rect 49086 38834 49138 38846
rect 49086 38770 49138 38782
rect 5294 38722 5346 38734
rect 8430 38722 8482 38734
rect 15710 38722 15762 38734
rect 17838 38722 17890 38734
rect 2482 38670 2494 38722
rect 2546 38670 2558 38722
rect 4610 38670 4622 38722
rect 4674 38670 4686 38722
rect 5842 38670 5854 38722
rect 5906 38670 5918 38722
rect 15362 38670 15374 38722
rect 15426 38670 15438 38722
rect 16146 38670 16158 38722
rect 16210 38670 16222 38722
rect 5294 38658 5346 38670
rect 8430 38658 8482 38670
rect 15710 38658 15762 38670
rect 17838 38658 17890 38670
rect 18734 38722 18786 38734
rect 22542 38722 22594 38734
rect 22082 38670 22094 38722
rect 22146 38670 22158 38722
rect 18734 38658 18786 38670
rect 22542 38658 22594 38670
rect 33742 38722 33794 38734
rect 33742 38658 33794 38670
rect 34302 38722 34354 38734
rect 34302 38658 34354 38670
rect 36206 38722 36258 38734
rect 36206 38658 36258 38670
rect 39902 38722 39954 38734
rect 39902 38658 39954 38670
rect 40238 38722 40290 38734
rect 40238 38658 40290 38670
rect 42030 38722 42082 38734
rect 42030 38658 42082 38670
rect 42926 38722 42978 38734
rect 45726 38722 45778 38734
rect 45266 38670 45278 38722
rect 45330 38670 45342 38722
rect 42926 38658 42978 38670
rect 45726 38658 45778 38670
rect 48190 38722 48242 38734
rect 48190 38658 48242 38670
rect 7534 38610 7586 38622
rect 7534 38546 7586 38558
rect 8766 38610 8818 38622
rect 8766 38546 8818 38558
rect 9998 38610 10050 38622
rect 9998 38546 10050 38558
rect 18398 38610 18450 38622
rect 18398 38546 18450 38558
rect 18846 38610 18898 38622
rect 18846 38546 18898 38558
rect 20302 38610 20354 38622
rect 20302 38546 20354 38558
rect 23998 38610 24050 38622
rect 23998 38546 24050 38558
rect 33182 38610 33234 38622
rect 33182 38546 33234 38558
rect 39790 38610 39842 38622
rect 39790 38546 39842 38558
rect 44942 38610 44994 38622
rect 44942 38546 44994 38558
rect 46062 38610 46114 38622
rect 46062 38546 46114 38558
rect 1344 38442 49616 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 49616 38442
rect 1344 38356 49616 38390
rect 2606 38274 2658 38286
rect 2606 38210 2658 38222
rect 2942 38274 2994 38286
rect 13918 38274 13970 38286
rect 13570 38222 13582 38274
rect 13634 38222 13646 38274
rect 2942 38210 2994 38222
rect 13918 38210 13970 38222
rect 21758 38274 21810 38286
rect 21758 38210 21810 38222
rect 44942 38274 44994 38286
rect 45938 38222 45950 38274
rect 46002 38222 46014 38274
rect 44942 38210 44994 38222
rect 22766 38162 22818 38174
rect 27134 38162 27186 38174
rect 20290 38110 20302 38162
rect 20354 38110 20366 38162
rect 23314 38110 23326 38162
rect 23378 38110 23390 38162
rect 22766 38098 22818 38110
rect 27134 38098 27186 38110
rect 28590 38162 28642 38174
rect 36990 38162 37042 38174
rect 44158 38162 44210 38174
rect 29474 38110 29486 38162
rect 29538 38110 29550 38162
rect 33954 38110 33966 38162
rect 34018 38110 34030 38162
rect 37538 38110 37550 38162
rect 37602 38110 37614 38162
rect 39666 38110 39678 38162
rect 39730 38110 39742 38162
rect 43698 38110 43710 38162
rect 43762 38110 43774 38162
rect 28590 38098 28642 38110
rect 36990 38098 37042 38110
rect 44158 38098 44210 38110
rect 45390 38162 45442 38174
rect 47058 38110 47070 38162
rect 47122 38110 47134 38162
rect 49186 38110 49198 38162
rect 49250 38110 49262 38162
rect 45390 38098 45442 38110
rect 14142 38050 14194 38062
rect 10546 37998 10558 38050
rect 10610 37998 10622 38050
rect 14142 37986 14194 37998
rect 14814 38050 14866 38062
rect 14814 37986 14866 37998
rect 15150 38050 15202 38062
rect 15150 37986 15202 37998
rect 15934 38050 15986 38062
rect 15934 37986 15986 37998
rect 16046 38050 16098 38062
rect 17166 38050 17218 38062
rect 18174 38050 18226 38062
rect 21870 38050 21922 38062
rect 16930 37998 16942 38050
rect 16994 37998 17006 38050
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 17938 37998 17950 38050
rect 18002 37998 18014 38050
rect 19506 37998 19518 38050
rect 19570 37998 19582 38050
rect 20402 37998 20414 38050
rect 20466 37998 20478 38050
rect 16046 37986 16098 37998
rect 17166 37986 17218 37998
rect 18174 37986 18226 37998
rect 21870 37986 21922 37998
rect 22206 38050 22258 38062
rect 22206 37986 22258 37998
rect 22430 38050 22482 38062
rect 29598 38050 29650 38062
rect 30606 38050 30658 38062
rect 35646 38050 35698 38062
rect 45614 38050 45666 38062
rect 26226 37998 26238 38050
rect 26290 37998 26302 38050
rect 29362 37998 29374 38050
rect 29426 37998 29438 38050
rect 30034 37998 30046 38050
rect 30098 37998 30110 38050
rect 30930 37998 30942 38050
rect 30994 37998 31006 38050
rect 36194 37998 36206 38050
rect 36258 37998 36270 38050
rect 40338 37998 40350 38050
rect 40402 37998 40414 38050
rect 40898 37998 40910 38050
rect 40962 37998 40974 38050
rect 46274 37998 46286 38050
rect 46338 37998 46350 38050
rect 22430 37986 22482 37998
rect 29598 37986 29650 37998
rect 30606 37986 30658 37998
rect 35646 37986 35698 37998
rect 45614 37986 45666 37998
rect 2718 37938 2770 37950
rect 10894 37938 10946 37950
rect 5618 37886 5630 37938
rect 5682 37886 5694 37938
rect 2718 37874 2770 37886
rect 10894 37874 10946 37886
rect 15374 37938 15426 37950
rect 15374 37874 15426 37886
rect 15822 37938 15874 37950
rect 15822 37874 15874 37886
rect 18286 37938 18338 37950
rect 19070 37938 19122 37950
rect 26574 37938 26626 37950
rect 34862 37938 34914 37950
rect 18722 37886 18734 37938
rect 18786 37886 18798 37938
rect 20066 37886 20078 37938
rect 20130 37886 20142 37938
rect 25442 37886 25454 37938
rect 25506 37886 25518 37938
rect 31714 37886 31726 37938
rect 31778 37886 31790 37938
rect 18286 37874 18338 37886
rect 19070 37874 19122 37886
rect 26574 37874 26626 37886
rect 34862 37874 34914 37886
rect 34974 37938 35026 37950
rect 34974 37874 35026 37886
rect 35086 37938 35138 37950
rect 35086 37874 35138 37886
rect 35758 37938 35810 37950
rect 45054 37938 45106 37950
rect 41570 37886 41582 37938
rect 41634 37886 41646 37938
rect 35758 37874 35810 37886
rect 45054 37874 45106 37886
rect 5966 37826 6018 37838
rect 5966 37762 6018 37774
rect 10782 37826 10834 37838
rect 10782 37762 10834 37774
rect 15038 37826 15090 37838
rect 17278 37826 17330 37838
rect 16482 37774 16494 37826
rect 16546 37774 16558 37826
rect 15038 37762 15090 37774
rect 17278 37762 17330 37774
rect 17390 37826 17442 37838
rect 17390 37762 17442 37774
rect 21758 37826 21810 37838
rect 21758 37762 21810 37774
rect 22654 37826 22706 37838
rect 22654 37762 22706 37774
rect 22878 37826 22930 37838
rect 22878 37762 22930 37774
rect 26686 37826 26738 37838
rect 26686 37762 26738 37774
rect 27918 37826 27970 37838
rect 27918 37762 27970 37774
rect 29822 37826 29874 37838
rect 35870 37826 35922 37838
rect 34402 37774 34414 37826
rect 34466 37774 34478 37826
rect 29822 37762 29874 37774
rect 35870 37762 35922 37774
rect 35982 37826 36034 37838
rect 35982 37762 36034 37774
rect 37102 37826 37154 37838
rect 37102 37762 37154 37774
rect 44270 37826 44322 37838
rect 44270 37762 44322 37774
rect 1344 37658 49616 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 49616 37658
rect 1344 37572 49616 37606
rect 1934 37490 1986 37502
rect 1934 37426 1986 37438
rect 3278 37490 3330 37502
rect 18958 37490 19010 37502
rect 17938 37438 17950 37490
rect 18002 37438 18014 37490
rect 3278 37426 3330 37438
rect 18958 37426 19010 37438
rect 19182 37490 19234 37502
rect 19182 37426 19234 37438
rect 24670 37490 24722 37502
rect 24670 37426 24722 37438
rect 25454 37490 25506 37502
rect 25454 37426 25506 37438
rect 26462 37490 26514 37502
rect 26462 37426 26514 37438
rect 26574 37490 26626 37502
rect 26574 37426 26626 37438
rect 27806 37490 27858 37502
rect 27806 37426 27858 37438
rect 28254 37490 28306 37502
rect 28254 37426 28306 37438
rect 28814 37490 28866 37502
rect 28814 37426 28866 37438
rect 29934 37490 29986 37502
rect 32398 37490 32450 37502
rect 31042 37438 31054 37490
rect 31106 37438 31118 37490
rect 32050 37438 32062 37490
rect 32114 37438 32126 37490
rect 29934 37426 29986 37438
rect 32398 37426 32450 37438
rect 39678 37490 39730 37502
rect 39678 37426 39730 37438
rect 41022 37490 41074 37502
rect 41022 37426 41074 37438
rect 45726 37490 45778 37502
rect 45726 37426 45778 37438
rect 3502 37378 3554 37390
rect 16158 37378 16210 37390
rect 4610 37326 4622 37378
rect 4674 37326 4686 37378
rect 6402 37326 6414 37378
rect 6466 37326 6478 37378
rect 11778 37326 11790 37378
rect 11842 37326 11854 37378
rect 3502 37314 3554 37326
rect 16158 37314 16210 37326
rect 16382 37378 16434 37390
rect 16382 37314 16434 37326
rect 17390 37378 17442 37390
rect 17390 37314 17442 37326
rect 25678 37378 25730 37390
rect 25678 37314 25730 37326
rect 29486 37378 29538 37390
rect 29486 37314 29538 37326
rect 30494 37378 30546 37390
rect 30494 37314 30546 37326
rect 32510 37378 32562 37390
rect 40238 37378 40290 37390
rect 45166 37378 45218 37390
rect 33842 37326 33854 37378
rect 33906 37326 33918 37378
rect 37090 37326 37102 37378
rect 37154 37326 37166 37378
rect 42690 37326 42702 37378
rect 42754 37326 42766 37378
rect 32510 37314 32562 37326
rect 40238 37314 40290 37326
rect 45166 37314 45218 37326
rect 45614 37378 45666 37390
rect 47954 37326 47966 37378
rect 48018 37326 48030 37378
rect 48738 37326 48750 37378
rect 48802 37326 48814 37378
rect 45614 37314 45666 37326
rect 2270 37266 2322 37278
rect 4958 37266 5010 37278
rect 3042 37214 3054 37266
rect 3106 37214 3118 37266
rect 2270 37202 2322 37214
rect 4958 37202 5010 37214
rect 6078 37266 6130 37278
rect 8542 37266 8594 37278
rect 17614 37266 17666 37278
rect 8082 37214 8094 37266
rect 8146 37214 8158 37266
rect 12450 37214 12462 37266
rect 12514 37214 12526 37266
rect 12898 37214 12910 37266
rect 12962 37214 12974 37266
rect 6078 37202 6130 37214
rect 8542 37202 8594 37214
rect 17614 37202 17666 37214
rect 18510 37266 18562 37278
rect 26686 37266 26738 37278
rect 19730 37214 19742 37266
rect 19794 37214 19806 37266
rect 21858 37214 21870 37266
rect 21922 37214 21934 37266
rect 22530 37214 22542 37266
rect 22594 37214 22606 37266
rect 23090 37214 23102 37266
rect 23154 37214 23166 37266
rect 25218 37214 25230 37266
rect 25282 37214 25294 37266
rect 25890 37214 25902 37266
rect 25954 37214 25966 37266
rect 26226 37214 26238 37266
rect 26290 37214 26302 37266
rect 18510 37202 18562 37214
rect 26686 37202 26738 37214
rect 26798 37266 26850 37278
rect 26798 37202 26850 37214
rect 27470 37266 27522 37278
rect 27470 37202 27522 37214
rect 29150 37266 29202 37278
rect 31726 37266 31778 37278
rect 39790 37266 39842 37278
rect 31266 37214 31278 37266
rect 31330 37214 31342 37266
rect 33058 37214 33070 37266
rect 33122 37214 33134 37266
rect 36418 37214 36430 37266
rect 36482 37214 36494 37266
rect 29150 37202 29202 37214
rect 31726 37202 31778 37214
rect 39790 37202 39842 37214
rect 40014 37266 40066 37278
rect 46846 37266 46898 37278
rect 41906 37214 41918 37266
rect 41970 37214 41982 37266
rect 45378 37214 45390 37266
rect 45442 37214 45454 37266
rect 46610 37214 46622 37266
rect 46674 37214 46686 37266
rect 40014 37202 40066 37214
rect 46846 37202 46898 37214
rect 47630 37266 47682 37278
rect 47630 37202 47682 37214
rect 49086 37266 49138 37278
rect 49086 37202 49138 37214
rect 16270 37154 16322 37166
rect 9650 37102 9662 37154
rect 9714 37102 9726 37154
rect 13682 37102 13694 37154
rect 13746 37102 13758 37154
rect 15810 37102 15822 37154
rect 15874 37102 15886 37154
rect 16270 37090 16322 37102
rect 19070 37154 19122 37166
rect 24558 37154 24610 37166
rect 20738 37102 20750 37154
rect 20802 37102 20814 37154
rect 19070 37090 19122 37102
rect 24558 37090 24610 37102
rect 25566 37154 25618 37166
rect 39902 37154 39954 37166
rect 35970 37102 35982 37154
rect 36034 37102 36046 37154
rect 39218 37102 39230 37154
rect 39282 37102 39294 37154
rect 25566 37090 25618 37102
rect 39902 37090 39954 37102
rect 40910 37154 40962 37166
rect 40910 37090 40962 37102
rect 41470 37154 41522 37166
rect 44818 37102 44830 37154
rect 44882 37102 44894 37154
rect 41470 37090 41522 37102
rect 3614 37042 3666 37054
rect 3614 36978 3666 36990
rect 8318 37042 8370 37054
rect 8318 36978 8370 36990
rect 8654 37042 8706 37054
rect 30270 37042 30322 37054
rect 20626 36990 20638 37042
rect 20690 36990 20702 37042
rect 8654 36978 8706 36990
rect 30270 36978 30322 36990
rect 30606 37042 30658 37054
rect 46722 36990 46734 37042
rect 46786 36990 46798 37042
rect 30606 36978 30658 36990
rect 1344 36874 49616 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 49616 36874
rect 1344 36788 49616 36822
rect 14926 36706 14978 36718
rect 46062 36706 46114 36718
rect 10882 36654 10894 36706
rect 10946 36654 10958 36706
rect 28578 36654 28590 36706
rect 28642 36654 28654 36706
rect 14926 36642 14978 36654
rect 46062 36642 46114 36654
rect 17614 36594 17666 36606
rect 28030 36594 28082 36606
rect 32734 36594 32786 36606
rect 45054 36594 45106 36606
rect 4610 36542 4622 36594
rect 4674 36542 4686 36594
rect 6290 36542 6302 36594
rect 6354 36542 6366 36594
rect 8418 36542 8430 36594
rect 8482 36542 8494 36594
rect 10210 36542 10222 36594
rect 10274 36542 10286 36594
rect 19730 36542 19742 36594
rect 19794 36542 19806 36594
rect 24658 36542 24670 36594
rect 24722 36542 24734 36594
rect 26786 36542 26798 36594
rect 26850 36542 26862 36594
rect 29138 36542 29150 36594
rect 29202 36542 29214 36594
rect 31266 36542 31278 36594
rect 31330 36542 31342 36594
rect 36418 36542 36430 36594
rect 36482 36542 36494 36594
rect 38770 36542 38782 36594
rect 38834 36542 38846 36594
rect 40002 36542 40014 36594
rect 40066 36542 40078 36594
rect 47058 36542 47070 36594
rect 47122 36542 47134 36594
rect 49186 36542 49198 36594
rect 49250 36542 49262 36594
rect 17614 36530 17666 36542
rect 28030 36530 28082 36542
rect 32734 36530 32786 36542
rect 45054 36530 45106 36542
rect 11230 36482 11282 36494
rect 1810 36430 1822 36482
rect 1874 36430 1886 36482
rect 9202 36430 9214 36482
rect 9266 36430 9278 36482
rect 10546 36430 10558 36482
rect 10610 36430 10622 36482
rect 11230 36418 11282 36430
rect 11566 36482 11618 36494
rect 11566 36418 11618 36430
rect 11790 36482 11842 36494
rect 14142 36482 14194 36494
rect 12674 36430 12686 36482
rect 12738 36430 12750 36482
rect 11790 36418 11842 36430
rect 14142 36418 14194 36430
rect 14366 36482 14418 36494
rect 14366 36418 14418 36430
rect 14702 36482 14754 36494
rect 17838 36482 17890 36494
rect 23326 36482 23378 36494
rect 28254 36482 28306 36494
rect 33294 36482 33346 36494
rect 37550 36482 37602 36494
rect 15250 36430 15262 36482
rect 15314 36430 15326 36482
rect 15810 36430 15822 36482
rect 15874 36430 15886 36482
rect 19282 36430 19294 36482
rect 19346 36430 19358 36482
rect 20066 36430 20078 36482
rect 20130 36430 20142 36482
rect 22306 36430 22318 36482
rect 22370 36430 22382 36482
rect 22866 36430 22878 36482
rect 22930 36430 22942 36482
rect 27570 36430 27582 36482
rect 27634 36430 27646 36482
rect 31938 36430 31950 36482
rect 32002 36430 32014 36482
rect 33618 36430 33630 36482
rect 33682 36430 33694 36482
rect 14702 36418 14754 36430
rect 17838 36418 17890 36430
rect 23326 36418 23378 36430
rect 28254 36418 28306 36430
rect 33294 36418 33346 36430
rect 37550 36418 37602 36430
rect 38334 36482 38386 36494
rect 38334 36418 38386 36430
rect 38446 36482 38498 36494
rect 38446 36418 38498 36430
rect 38670 36482 38722 36494
rect 43486 36482 43538 36494
rect 38882 36430 38894 36482
rect 38946 36430 38958 36482
rect 39890 36430 39902 36482
rect 39954 36430 39966 36482
rect 40898 36430 40910 36482
rect 40962 36430 40974 36482
rect 38670 36418 38722 36430
rect 43486 36418 43538 36430
rect 45278 36482 45330 36494
rect 45278 36418 45330 36430
rect 45390 36482 45442 36494
rect 45390 36418 45442 36430
rect 45838 36482 45890 36494
rect 46274 36430 46286 36482
rect 46338 36430 46350 36482
rect 45838 36418 45890 36430
rect 5070 36370 5122 36382
rect 37326 36370 37378 36382
rect 2482 36318 2494 36370
rect 2546 36318 2558 36370
rect 13794 36318 13806 36370
rect 13858 36318 13870 36370
rect 19170 36318 19182 36370
rect 19234 36318 19246 36370
rect 21858 36318 21870 36370
rect 21922 36318 21934 36370
rect 23874 36318 23886 36370
rect 23938 36318 23950 36370
rect 34290 36318 34302 36370
rect 34354 36318 34366 36370
rect 5070 36306 5122 36318
rect 37326 36306 37378 36318
rect 40350 36370 40402 36382
rect 41694 36370 41746 36382
rect 43598 36370 43650 36382
rect 40674 36318 40686 36370
rect 40738 36318 40750 36370
rect 42802 36318 42814 36370
rect 42866 36318 42878 36370
rect 40350 36306 40402 36318
rect 41694 36306 41746 36318
rect 43598 36306 43650 36318
rect 44046 36370 44098 36382
rect 44046 36306 44098 36318
rect 4958 36258 5010 36270
rect 4958 36194 5010 36206
rect 11454 36258 11506 36270
rect 11454 36194 11506 36206
rect 12910 36258 12962 36270
rect 12910 36194 12962 36206
rect 15598 36258 15650 36270
rect 21646 36258 21698 36270
rect 18162 36206 18174 36258
rect 18226 36206 18238 36258
rect 15598 36194 15650 36206
rect 21646 36194 21698 36206
rect 24110 36258 24162 36270
rect 24110 36194 24162 36206
rect 32622 36258 32674 36270
rect 32622 36194 32674 36206
rect 32846 36258 32898 36270
rect 41358 36258 41410 36270
rect 37874 36206 37886 36258
rect 37938 36206 37950 36258
rect 32846 36194 32898 36206
rect 41358 36194 41410 36206
rect 42142 36258 42194 36270
rect 42142 36194 42194 36206
rect 43150 36258 43202 36270
rect 43150 36194 43202 36206
rect 43822 36258 43874 36270
rect 43822 36194 43874 36206
rect 44158 36258 44210 36270
rect 44158 36194 44210 36206
rect 44382 36258 44434 36270
rect 44382 36194 44434 36206
rect 1344 36090 49616 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 49616 36090
rect 1344 36004 49616 36038
rect 2606 35922 2658 35934
rect 22430 35922 22482 35934
rect 7746 35870 7758 35922
rect 7810 35870 7822 35922
rect 2606 35858 2658 35870
rect 22430 35858 22482 35870
rect 22654 35922 22706 35934
rect 22654 35858 22706 35870
rect 22878 35922 22930 35934
rect 22878 35858 22930 35870
rect 23998 35922 24050 35934
rect 23998 35858 24050 35870
rect 24558 35922 24610 35934
rect 24558 35858 24610 35870
rect 31726 35922 31778 35934
rect 31726 35858 31778 35870
rect 32510 35922 32562 35934
rect 32510 35858 32562 35870
rect 40126 35922 40178 35934
rect 40126 35858 40178 35870
rect 40238 35922 40290 35934
rect 49086 35922 49138 35934
rect 48738 35870 48750 35922
rect 48802 35870 48814 35922
rect 40238 35858 40290 35870
rect 49086 35858 49138 35870
rect 6638 35810 6690 35822
rect 6638 35746 6690 35758
rect 6862 35810 6914 35822
rect 15262 35810 15314 35822
rect 23326 35810 23378 35822
rect 8866 35758 8878 35810
rect 8930 35758 8942 35810
rect 22082 35758 22094 35810
rect 22146 35758 22158 35810
rect 6862 35746 6914 35758
rect 15262 35746 15314 35758
rect 23326 35746 23378 35758
rect 27918 35810 27970 35822
rect 38670 35810 38722 35822
rect 33618 35758 33630 35810
rect 33682 35758 33694 35810
rect 27918 35746 27970 35758
rect 38670 35746 38722 35758
rect 40910 35810 40962 35822
rect 40910 35746 40962 35758
rect 7422 35698 7474 35710
rect 8654 35698 8706 35710
rect 21422 35698 21474 35710
rect 3378 35646 3390 35698
rect 3442 35646 3454 35698
rect 8306 35646 8318 35698
rect 8370 35646 8382 35698
rect 14802 35646 14814 35698
rect 14866 35646 14878 35698
rect 15922 35646 15934 35698
rect 15986 35646 15998 35698
rect 17714 35646 17726 35698
rect 17778 35646 17790 35698
rect 7422 35634 7474 35646
rect 8654 35634 8706 35646
rect 21422 35634 21474 35646
rect 21534 35698 21586 35710
rect 21534 35634 21586 35646
rect 21646 35698 21698 35710
rect 21646 35634 21698 35646
rect 22542 35698 22594 35710
rect 24110 35698 24162 35710
rect 23538 35646 23550 35698
rect 23602 35646 23614 35698
rect 22542 35634 22594 35646
rect 24110 35634 24162 35646
rect 27358 35698 27410 35710
rect 27358 35634 27410 35646
rect 27582 35698 27634 35710
rect 27582 35634 27634 35646
rect 28030 35698 28082 35710
rect 30270 35698 30322 35710
rect 28578 35646 28590 35698
rect 28642 35646 28654 35698
rect 28030 35634 28082 35646
rect 30270 35634 30322 35646
rect 31614 35698 31666 35710
rect 32274 35646 32286 35698
rect 32338 35646 32350 35698
rect 36978 35646 36990 35698
rect 37042 35646 37054 35698
rect 39330 35646 39342 35698
rect 39394 35646 39406 35698
rect 41234 35646 41246 35698
rect 41298 35646 41310 35698
rect 45826 35646 45838 35698
rect 45890 35646 45902 35698
rect 31614 35634 31666 35646
rect 7198 35586 7250 35598
rect 4050 35534 4062 35586
rect 4114 35534 4126 35586
rect 6178 35534 6190 35586
rect 6242 35534 6254 35586
rect 6514 35534 6526 35586
rect 6578 35534 6590 35586
rect 7198 35522 7250 35534
rect 8990 35586 9042 35598
rect 16718 35586 16770 35598
rect 20974 35586 21026 35598
rect 9874 35534 9886 35586
rect 9938 35534 9950 35586
rect 16146 35534 16158 35586
rect 16210 35534 16222 35586
rect 18386 35534 18398 35586
rect 18450 35534 18462 35586
rect 20514 35534 20526 35586
rect 20578 35534 20590 35586
rect 8990 35522 9042 35534
rect 16718 35522 16770 35534
rect 20974 35522 21026 35534
rect 26798 35586 26850 35598
rect 26798 35522 26850 35534
rect 29262 35586 29314 35598
rect 29262 35522 29314 35534
rect 29710 35586 29762 35598
rect 41694 35586 41746 35598
rect 48190 35586 48242 35598
rect 39442 35534 39454 35586
rect 39506 35534 39518 35586
rect 45266 35534 45278 35586
rect 45330 35534 45342 35586
rect 29710 35522 29762 35534
rect 41694 35522 41746 35534
rect 48190 35522 48242 35534
rect 2270 35474 2322 35486
rect 2270 35410 2322 35422
rect 2494 35474 2546 35486
rect 2494 35410 2546 35422
rect 2606 35474 2658 35486
rect 2606 35410 2658 35422
rect 7982 35474 8034 35486
rect 29374 35474 29426 35486
rect 27010 35422 27022 35474
rect 27074 35422 27086 35474
rect 7982 35410 8034 35422
rect 29374 35410 29426 35422
rect 29822 35474 29874 35486
rect 29822 35410 29874 35422
rect 30158 35474 30210 35486
rect 30158 35410 30210 35422
rect 31726 35474 31778 35486
rect 31726 35410 31778 35422
rect 40350 35474 40402 35486
rect 40350 35410 40402 35422
rect 41246 35474 41298 35486
rect 47966 35474 48018 35486
rect 47618 35422 47630 35474
rect 47682 35422 47694 35474
rect 41246 35410 41298 35422
rect 47966 35410 48018 35422
rect 1344 35306 49616 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 49616 35306
rect 1344 35220 49616 35254
rect 3502 35138 3554 35150
rect 2594 35086 2606 35138
rect 2658 35086 2670 35138
rect 3502 35074 3554 35086
rect 9214 35138 9266 35150
rect 9214 35074 9266 35086
rect 9326 35138 9378 35150
rect 9326 35074 9378 35086
rect 27470 35138 27522 35150
rect 27470 35074 27522 35086
rect 30382 35138 30434 35150
rect 30382 35074 30434 35086
rect 44158 35138 44210 35150
rect 44158 35074 44210 35086
rect 3166 35026 3218 35038
rect 3166 34962 3218 34974
rect 3614 35026 3666 35038
rect 3614 34962 3666 34974
rect 5070 35026 5122 35038
rect 18286 35026 18338 35038
rect 36094 35026 36146 35038
rect 49086 35026 49138 35038
rect 8530 34974 8542 35026
rect 8594 34974 8606 35026
rect 12674 34974 12686 35026
rect 12738 34974 12750 35026
rect 14242 34974 14254 35026
rect 14306 34974 14318 35026
rect 16370 34974 16382 35026
rect 16434 34974 16446 35026
rect 20402 34974 20414 35026
rect 20466 34974 20478 35026
rect 32610 34974 32622 35026
rect 32674 34974 32686 35026
rect 34738 34974 34750 35026
rect 34802 34974 34814 35026
rect 35410 34974 35422 35026
rect 35474 34974 35486 35026
rect 37314 34974 37326 35026
rect 37378 34974 37390 35026
rect 39442 34974 39454 35026
rect 39506 34974 39518 35026
rect 41682 34974 41694 35026
rect 41746 34974 41758 35026
rect 43810 34974 43822 35026
rect 43874 34974 43886 35026
rect 44818 34974 44830 35026
rect 44882 34974 44894 35026
rect 48178 34974 48190 35026
rect 48242 34974 48254 35026
rect 5070 34962 5122 34974
rect 18286 34962 18338 34974
rect 36094 34962 36146 34974
rect 49086 34962 49138 34974
rect 2942 34914 2994 34926
rect 2942 34850 2994 34862
rect 4286 34914 4338 34926
rect 8990 34914 9042 34926
rect 28366 34914 28418 34926
rect 5618 34862 5630 34914
rect 5682 34862 5694 34914
rect 9874 34862 9886 34914
rect 9938 34862 9950 34914
rect 13458 34862 13470 34914
rect 13522 34862 13534 34914
rect 17826 34862 17838 34914
rect 17890 34862 17902 34914
rect 18050 34862 18062 34914
rect 18114 34862 18126 34914
rect 18834 34862 18846 34914
rect 18898 34862 18910 34914
rect 20514 34862 20526 34914
rect 20578 34862 20590 34914
rect 22978 34862 22990 34914
rect 23042 34862 23054 34914
rect 4286 34850 4338 34862
rect 8990 34850 9042 34862
rect 28366 34850 28418 34862
rect 29486 34914 29538 34926
rect 29486 34850 29538 34862
rect 30046 34914 30098 34926
rect 31938 34862 31950 34914
rect 32002 34862 32014 34914
rect 35074 34862 35086 34914
rect 35138 34862 35150 34914
rect 40226 34862 40238 34914
rect 40290 34862 40302 34914
rect 41010 34862 41022 34914
rect 41074 34862 41086 34914
rect 47618 34862 47630 34914
rect 47682 34862 47694 34914
rect 48402 34862 48414 34914
rect 48466 34862 48478 34914
rect 30046 34850 30098 34862
rect 4734 34802 4786 34814
rect 1922 34750 1934 34802
rect 1986 34750 1998 34802
rect 4734 34738 4786 34750
rect 4846 34802 4898 34814
rect 18622 34802 18674 34814
rect 27694 34802 27746 34814
rect 6402 34750 6414 34802
rect 6466 34750 6478 34802
rect 10546 34750 10558 34802
rect 10610 34750 10622 34802
rect 23538 34750 23550 34802
rect 23602 34750 23614 34802
rect 4846 34738 4898 34750
rect 18622 34738 18674 34750
rect 27694 34738 27746 34750
rect 28030 34802 28082 34814
rect 28030 34738 28082 34750
rect 29150 34802 29202 34814
rect 29150 34738 29202 34750
rect 29822 34802 29874 34814
rect 29822 34738 29874 34750
rect 44270 34802 44322 34814
rect 46946 34750 46958 34802
rect 47010 34750 47022 34802
rect 44270 34738 44322 34750
rect 2270 34690 2322 34702
rect 2270 34626 2322 34638
rect 3726 34690 3778 34702
rect 3726 34626 3778 34638
rect 4062 34690 4114 34702
rect 4062 34626 4114 34638
rect 9326 34690 9378 34702
rect 29262 34690 29314 34702
rect 27122 34638 27134 34690
rect 27186 34638 27198 34690
rect 9326 34626 9378 34638
rect 29262 34626 29314 34638
rect 35982 34690 36034 34702
rect 35982 34626 36034 34638
rect 1344 34522 49616 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 49616 34522
rect 1344 34436 49616 34470
rect 1934 34354 1986 34366
rect 1934 34290 1986 34302
rect 4174 34354 4226 34366
rect 4174 34290 4226 34302
rect 5630 34354 5682 34366
rect 5630 34290 5682 34302
rect 6414 34354 6466 34366
rect 6414 34290 6466 34302
rect 7758 34354 7810 34366
rect 14254 34354 14306 34366
rect 10098 34302 10110 34354
rect 10162 34302 10174 34354
rect 7758 34290 7810 34302
rect 14254 34290 14306 34302
rect 18062 34354 18114 34366
rect 24334 34354 24386 34366
rect 19842 34302 19854 34354
rect 19906 34302 19918 34354
rect 18062 34290 18114 34302
rect 24334 34290 24386 34302
rect 28590 34354 28642 34366
rect 28590 34290 28642 34302
rect 29486 34354 29538 34366
rect 29486 34290 29538 34302
rect 30382 34354 30434 34366
rect 41134 34354 41186 34366
rect 33394 34302 33406 34354
rect 33458 34302 33470 34354
rect 40226 34302 40238 34354
rect 40290 34302 40302 34354
rect 30382 34290 30434 34302
rect 41134 34290 41186 34302
rect 43934 34354 43986 34366
rect 47182 34354 47234 34366
rect 44370 34302 44382 34354
rect 44434 34302 44446 34354
rect 43934 34290 43986 34302
rect 47182 34290 47234 34302
rect 47406 34354 47458 34366
rect 47406 34290 47458 34302
rect 48190 34354 48242 34366
rect 48190 34290 48242 34302
rect 48862 34354 48914 34366
rect 48862 34290 48914 34302
rect 1710 34242 1762 34254
rect 1710 34178 1762 34190
rect 2270 34242 2322 34254
rect 2270 34178 2322 34190
rect 2718 34242 2770 34254
rect 2718 34178 2770 34190
rect 2830 34242 2882 34254
rect 2830 34178 2882 34190
rect 4062 34242 4114 34254
rect 4062 34178 4114 34190
rect 6302 34242 6354 34254
rect 6302 34178 6354 34190
rect 7310 34242 7362 34254
rect 7310 34178 7362 34190
rect 7870 34242 7922 34254
rect 28702 34242 28754 34254
rect 9650 34190 9662 34242
rect 9714 34190 9726 34242
rect 11218 34190 11230 34242
rect 11282 34190 11294 34242
rect 21634 34190 21646 34242
rect 21698 34190 21710 34242
rect 7870 34178 7922 34190
rect 28702 34178 28754 34190
rect 30606 34242 30658 34254
rect 30606 34178 30658 34190
rect 31502 34242 31554 34254
rect 40910 34242 40962 34254
rect 36194 34190 36206 34242
rect 36258 34190 36270 34242
rect 37426 34190 37438 34242
rect 37490 34190 37502 34242
rect 39554 34190 39566 34242
rect 39618 34190 39630 34242
rect 39890 34190 39902 34242
rect 39954 34190 39966 34242
rect 31502 34178 31554 34190
rect 40910 34178 40962 34190
rect 48750 34242 48802 34254
rect 48750 34178 48802 34190
rect 2046 34130 2098 34142
rect 2046 34066 2098 34078
rect 2942 34130 2994 34142
rect 2942 34066 2994 34078
rect 4398 34130 4450 34142
rect 4398 34066 4450 34078
rect 4510 34130 4562 34142
rect 5966 34130 6018 34142
rect 14590 34130 14642 34142
rect 4610 34078 4622 34130
rect 4674 34078 4686 34130
rect 6626 34078 6638 34130
rect 6690 34078 6702 34130
rect 9538 34078 9550 34130
rect 9602 34078 9614 34130
rect 10546 34078 10558 34130
rect 10610 34078 10622 34130
rect 4510 34066 4562 34078
rect 5966 34066 6018 34078
rect 14590 34066 14642 34078
rect 15934 34130 15986 34142
rect 15934 34066 15986 34078
rect 16158 34130 16210 34142
rect 16158 34066 16210 34078
rect 17390 34130 17442 34142
rect 28366 34130 28418 34142
rect 20850 34078 20862 34130
rect 20914 34078 20926 34130
rect 25218 34078 25230 34130
rect 25282 34078 25294 34130
rect 17390 34066 17442 34078
rect 28366 34066 28418 34078
rect 29262 34130 29314 34142
rect 33070 34130 33122 34142
rect 43038 34130 43090 34142
rect 29698 34078 29710 34130
rect 29762 34078 29774 34130
rect 29922 34078 29934 34130
rect 29986 34078 29998 34130
rect 30930 34078 30942 34130
rect 30994 34078 31006 34130
rect 32162 34078 32174 34130
rect 32226 34078 32238 34130
rect 34738 34078 34750 34130
rect 34802 34078 34814 34130
rect 36978 34078 36990 34130
rect 37042 34078 37054 34130
rect 39218 34078 39230 34130
rect 39282 34078 39294 34130
rect 42466 34078 42478 34130
rect 42530 34078 42542 34130
rect 29262 34066 29314 34078
rect 33070 34066 33122 34078
rect 43038 34066 43090 34078
rect 43710 34130 43762 34142
rect 43710 34066 43762 34078
rect 44718 34130 44770 34142
rect 44718 34066 44770 34078
rect 45390 34130 45442 34142
rect 45390 34066 45442 34078
rect 45502 34130 45554 34142
rect 45502 34066 45554 34078
rect 45726 34130 45778 34142
rect 45726 34066 45778 34078
rect 47070 34130 47122 34142
rect 49074 34078 49086 34130
rect 49138 34078 49150 34130
rect 47070 34066 47122 34078
rect 12126 34018 12178 34030
rect 12126 33954 12178 33966
rect 18622 34018 18674 34030
rect 18622 33954 18674 33966
rect 18846 34018 18898 34030
rect 18846 33954 18898 33966
rect 19294 34018 19346 34030
rect 19294 33954 19346 33966
rect 20414 34018 20466 34030
rect 24446 34018 24498 34030
rect 30494 34018 30546 34030
rect 33966 34018 34018 34030
rect 23762 33966 23774 34018
rect 23826 33966 23838 34018
rect 26002 33966 26014 34018
rect 26066 33966 26078 34018
rect 28130 33966 28142 34018
rect 28194 33966 28206 34018
rect 29586 33966 29598 34018
rect 29650 33966 29662 34018
rect 31938 33966 31950 34018
rect 32002 33966 32014 34018
rect 20414 33954 20466 33966
rect 24446 33954 24498 33966
rect 30494 33954 30546 33966
rect 33966 33954 34018 33966
rect 34526 34018 34578 34030
rect 38446 34018 38498 34030
rect 35634 33966 35646 34018
rect 35698 33966 35710 34018
rect 34526 33954 34578 33966
rect 38446 33954 38498 33966
rect 38894 34018 38946 34030
rect 46734 34018 46786 34030
rect 42802 33966 42814 34018
rect 42866 33966 42878 34018
rect 46162 33966 46174 34018
rect 46226 33966 46238 34018
rect 38894 33954 38946 33966
rect 46734 33954 46786 33966
rect 47630 34018 47682 34030
rect 47630 33954 47682 33966
rect 7198 33906 7250 33918
rect 3378 33854 3390 33906
rect 3442 33854 3454 33906
rect 7198 33842 7250 33854
rect 7758 33906 7810 33918
rect 11902 33906 11954 33918
rect 17502 33906 17554 33918
rect 11554 33854 11566 33906
rect 11618 33854 11630 33906
rect 16482 33854 16494 33906
rect 16546 33854 16558 33906
rect 7758 33842 7810 33854
rect 11902 33842 11954 33854
rect 17502 33842 17554 33854
rect 18958 33906 19010 33918
rect 18958 33842 19010 33854
rect 19518 33906 19570 33918
rect 19518 33842 19570 33854
rect 41246 33906 41298 33918
rect 41246 33842 41298 33854
rect 44046 33906 44098 33918
rect 44046 33842 44098 33854
rect 45838 33906 45890 33918
rect 45838 33842 45890 33854
rect 46510 33906 46562 33918
rect 46510 33842 46562 33854
rect 1344 33738 49616 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 49616 33738
rect 1344 33652 49616 33686
rect 5854 33570 5906 33582
rect 5854 33506 5906 33518
rect 6078 33570 6130 33582
rect 6078 33506 6130 33518
rect 6302 33570 6354 33582
rect 6302 33506 6354 33518
rect 17166 33570 17218 33582
rect 28254 33570 28306 33582
rect 20738 33518 20750 33570
rect 20802 33518 20814 33570
rect 17166 33506 17218 33518
rect 28254 33506 28306 33518
rect 30382 33570 30434 33582
rect 30706 33518 30718 33570
rect 30770 33518 30782 33570
rect 30382 33506 30434 33518
rect 8430 33458 8482 33470
rect 16830 33458 16882 33470
rect 22094 33458 22146 33470
rect 29486 33458 29538 33470
rect 5058 33406 5070 33458
rect 5122 33406 5134 33458
rect 12674 33406 12686 33458
rect 12738 33406 12750 33458
rect 18610 33406 18622 33458
rect 18674 33406 18686 33458
rect 19282 33406 19294 33458
rect 19346 33406 19358 33458
rect 23650 33406 23662 33458
rect 23714 33406 23726 33458
rect 8430 33394 8482 33406
rect 16830 33394 16882 33406
rect 22094 33394 22146 33406
rect 29486 33394 29538 33406
rect 33182 33458 33234 33470
rect 43710 33458 43762 33470
rect 36418 33406 36430 33458
rect 36482 33406 36494 33458
rect 40450 33406 40462 33458
rect 40514 33406 40526 33458
rect 42578 33406 42590 33458
rect 42642 33406 42654 33458
rect 47058 33406 47070 33458
rect 47122 33406 47134 33458
rect 49186 33406 49198 33458
rect 49250 33406 49262 33458
rect 33182 33394 33234 33406
rect 43710 33394 43762 33406
rect 7310 33346 7362 33358
rect 2146 33294 2158 33346
rect 2210 33294 2222 33346
rect 5618 33294 5630 33346
rect 5682 33294 5694 33346
rect 7310 33282 7362 33294
rect 7982 33346 8034 33358
rect 9102 33346 9154 33358
rect 8866 33294 8878 33346
rect 8930 33294 8942 33346
rect 7982 33282 8034 33294
rect 9102 33282 9154 33294
rect 9326 33346 9378 33358
rect 16270 33346 16322 33358
rect 9874 33294 9886 33346
rect 9938 33294 9950 33346
rect 15138 33294 15150 33346
rect 15202 33294 15214 33346
rect 9326 33282 9378 33294
rect 16270 33282 16322 33294
rect 18174 33346 18226 33358
rect 18174 33282 18226 33294
rect 20190 33346 20242 33358
rect 20190 33282 20242 33294
rect 20414 33346 20466 33358
rect 27246 33346 27298 33358
rect 24770 33294 24782 33346
rect 24834 33294 24846 33346
rect 26450 33294 26462 33346
rect 26514 33294 26526 33346
rect 20414 33282 20466 33294
rect 27246 33282 27298 33294
rect 27358 33346 27410 33358
rect 28478 33346 28530 33358
rect 27570 33294 27582 33346
rect 27634 33294 27646 33346
rect 28130 33294 28142 33346
rect 28194 33294 28206 33346
rect 27358 33282 27410 33294
rect 28478 33282 28530 33294
rect 29374 33346 29426 33358
rect 29374 33282 29426 33294
rect 29598 33346 29650 33358
rect 30158 33346 30210 33358
rect 44830 33346 44882 33358
rect 29810 33294 29822 33346
rect 29874 33294 29886 33346
rect 31826 33294 31838 33346
rect 31890 33294 31902 33346
rect 33618 33294 33630 33346
rect 33682 33294 33694 33346
rect 36978 33294 36990 33346
rect 37042 33294 37054 33346
rect 43362 33294 43374 33346
rect 43426 33294 43438 33346
rect 45378 33294 45390 33346
rect 45442 33294 45454 33346
rect 46386 33294 46398 33346
rect 46450 33294 46462 33346
rect 29598 33282 29650 33294
rect 30158 33282 30210 33294
rect 44830 33282 44882 33294
rect 6414 33234 6466 33246
rect 2930 33182 2942 33234
rect 2994 33182 3006 33234
rect 6414 33170 6466 33182
rect 6974 33234 7026 33246
rect 6974 33170 7026 33182
rect 7758 33234 7810 33246
rect 7758 33170 7810 33182
rect 9438 33234 9490 33246
rect 13806 33234 13858 33246
rect 16158 33234 16210 33246
rect 10546 33182 10558 33234
rect 10610 33182 10622 33234
rect 15698 33182 15710 33234
rect 15762 33182 15774 33234
rect 9438 33170 9490 33182
rect 13806 33170 13858 33182
rect 16158 33170 16210 33182
rect 16382 33234 16434 33246
rect 16382 33170 16434 33182
rect 17390 33234 17442 33246
rect 17390 33170 17442 33182
rect 19294 33234 19346 33246
rect 19294 33170 19346 33182
rect 19406 33234 19458 33246
rect 32062 33234 32114 33246
rect 45054 33234 45106 33246
rect 19618 33182 19630 33234
rect 19682 33182 19694 33234
rect 24658 33182 24670 33234
rect 24722 33182 24734 33234
rect 25890 33182 25902 33234
rect 25954 33182 25966 33234
rect 34290 33182 34302 33234
rect 34354 33182 34366 33234
rect 37762 33182 37774 33234
rect 37826 33182 37838 33234
rect 19406 33170 19458 33182
rect 32062 33170 32114 33182
rect 45054 33170 45106 33182
rect 45166 33234 45218 33246
rect 45166 33170 45218 33182
rect 45838 33234 45890 33246
rect 45838 33170 45890 33182
rect 6862 33122 6914 33134
rect 6862 33058 6914 33070
rect 7534 33122 7586 33134
rect 7534 33058 7586 33070
rect 13470 33122 13522 33134
rect 13470 33058 13522 33070
rect 15374 33122 15426 33134
rect 15374 33058 15426 33070
rect 18286 33122 18338 33134
rect 18286 33058 18338 33070
rect 18510 33122 18562 33134
rect 18510 33058 18562 33070
rect 18622 33122 18674 33134
rect 18622 33058 18674 33070
rect 19070 33122 19122 33134
rect 27918 33122 27970 33134
rect 26786 33070 26798 33122
rect 26850 33070 26862 33122
rect 19070 33058 19122 33070
rect 27918 33058 27970 33070
rect 29262 33122 29314 33134
rect 29262 33058 29314 33070
rect 31166 33122 31218 33134
rect 31166 33058 31218 33070
rect 32846 33122 32898 33134
rect 43822 33122 43874 33134
rect 40002 33070 40014 33122
rect 40066 33070 40078 33122
rect 32846 33058 32898 33070
rect 43822 33058 43874 33070
rect 1344 32954 49616 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 49616 32954
rect 1344 32868 49616 32902
rect 3166 32786 3218 32798
rect 3166 32722 3218 32734
rect 11006 32786 11058 32798
rect 11006 32722 11058 32734
rect 15710 32786 15762 32798
rect 15710 32722 15762 32734
rect 19294 32786 19346 32798
rect 19294 32722 19346 32734
rect 19406 32786 19458 32798
rect 19406 32722 19458 32734
rect 19742 32786 19794 32798
rect 19742 32722 19794 32734
rect 20078 32786 20130 32798
rect 20078 32722 20130 32734
rect 20862 32786 20914 32798
rect 20862 32722 20914 32734
rect 25790 32786 25842 32798
rect 25790 32722 25842 32734
rect 27470 32786 27522 32798
rect 27470 32722 27522 32734
rect 28702 32786 28754 32798
rect 28702 32722 28754 32734
rect 33294 32786 33346 32798
rect 33294 32722 33346 32734
rect 34302 32786 34354 32798
rect 34302 32722 34354 32734
rect 40910 32786 40962 32798
rect 40910 32722 40962 32734
rect 44942 32786 44994 32798
rect 44942 32722 44994 32734
rect 45166 32786 45218 32798
rect 45166 32722 45218 32734
rect 45278 32786 45330 32798
rect 45278 32722 45330 32734
rect 46286 32786 46338 32798
rect 46286 32722 46338 32734
rect 47294 32786 47346 32798
rect 47294 32722 47346 32734
rect 10110 32674 10162 32686
rect 17502 32674 17554 32686
rect 5506 32622 5518 32674
rect 5570 32622 5582 32674
rect 13122 32622 13134 32674
rect 13186 32622 13198 32674
rect 10110 32610 10162 32622
rect 17502 32610 17554 32622
rect 17614 32674 17666 32686
rect 17614 32610 17666 32622
rect 18062 32674 18114 32686
rect 18062 32610 18114 32622
rect 20302 32674 20354 32686
rect 20302 32610 20354 32622
rect 20414 32674 20466 32686
rect 20414 32610 20466 32622
rect 26910 32674 26962 32686
rect 26910 32610 26962 32622
rect 27022 32674 27074 32686
rect 27022 32610 27074 32622
rect 27694 32674 27746 32686
rect 27694 32610 27746 32622
rect 27806 32674 27858 32686
rect 27806 32610 27858 32622
rect 28254 32674 28306 32686
rect 28254 32610 28306 32622
rect 29374 32674 29426 32686
rect 29374 32610 29426 32622
rect 29710 32674 29762 32686
rect 29710 32610 29762 32622
rect 34750 32674 34802 32686
rect 45502 32674 45554 32686
rect 42130 32622 42142 32674
rect 42194 32622 42206 32674
rect 34750 32610 34802 32622
rect 45502 32610 45554 32622
rect 48078 32674 48130 32686
rect 48738 32622 48750 32674
rect 48802 32622 48814 32674
rect 48078 32610 48130 32622
rect 2270 32562 2322 32574
rect 10222 32562 10274 32574
rect 11118 32562 11170 32574
rect 16494 32562 16546 32574
rect 1810 32510 1822 32562
rect 1874 32510 1886 32562
rect 3266 32510 3278 32562
rect 3330 32510 3342 32562
rect 8866 32510 8878 32562
rect 8930 32510 8942 32562
rect 9762 32510 9774 32562
rect 9826 32510 9838 32562
rect 10770 32510 10782 32562
rect 10834 32510 10846 32562
rect 12450 32510 12462 32562
rect 12514 32510 12526 32562
rect 2270 32498 2322 32510
rect 10222 32498 10274 32510
rect 11118 32498 11170 32510
rect 16494 32498 16546 32510
rect 16606 32562 16658 32574
rect 17278 32562 17330 32574
rect 16818 32510 16830 32562
rect 16882 32510 16894 32562
rect 16606 32498 16658 32510
rect 17278 32498 17330 32510
rect 18286 32562 18338 32574
rect 18286 32498 18338 32510
rect 18510 32562 18562 32574
rect 19518 32562 19570 32574
rect 18722 32510 18734 32562
rect 18786 32510 18798 32562
rect 18510 32498 18562 32510
rect 19518 32498 19570 32510
rect 21198 32562 21250 32574
rect 28478 32562 28530 32574
rect 31502 32562 31554 32574
rect 21522 32510 21534 32562
rect 21586 32510 21598 32562
rect 25554 32510 25566 32562
rect 25618 32510 25630 32562
rect 27234 32510 27246 32562
rect 27298 32510 27310 32562
rect 28914 32510 28926 32562
rect 28978 32510 28990 32562
rect 21198 32498 21250 32510
rect 28478 32498 28530 32510
rect 31502 32498 31554 32510
rect 32062 32562 32114 32574
rect 32062 32498 32114 32510
rect 34190 32562 34242 32574
rect 34190 32498 34242 32510
rect 34526 32562 34578 32574
rect 46622 32562 46674 32574
rect 38882 32510 38894 32562
rect 38946 32510 38958 32562
rect 41458 32510 41470 32562
rect 41522 32510 41534 32562
rect 44706 32510 44718 32562
rect 44770 32510 44782 32562
rect 34526 32498 34578 32510
rect 46622 32498 46674 32510
rect 47070 32562 47122 32574
rect 47070 32498 47122 32510
rect 47406 32562 47458 32574
rect 47406 32498 47458 32510
rect 47630 32562 47682 32574
rect 47630 32498 47682 32510
rect 47966 32562 48018 32574
rect 47966 32498 48018 32510
rect 49086 32562 49138 32574
rect 49086 32498 49138 32510
rect 3054 32450 3106 32462
rect 3054 32386 3106 32398
rect 10446 32450 10498 32462
rect 15598 32450 15650 32462
rect 29822 32450 29874 32462
rect 15250 32398 15262 32450
rect 15314 32398 15326 32450
rect 18610 32398 18622 32450
rect 18674 32398 18686 32450
rect 22306 32398 22318 32450
rect 22370 32398 22382 32450
rect 24434 32398 24446 32450
rect 24498 32398 24510 32450
rect 28802 32398 28814 32450
rect 28866 32398 28878 32450
rect 10446 32386 10498 32398
rect 15598 32386 15650 32398
rect 29822 32386 29874 32398
rect 30718 32450 30770 32462
rect 30718 32386 30770 32398
rect 31278 32450 31330 32462
rect 31278 32386 31330 32398
rect 32622 32450 32674 32462
rect 32622 32386 32674 32398
rect 33182 32450 33234 32462
rect 33182 32386 33234 32398
rect 33742 32450 33794 32462
rect 33742 32386 33794 32398
rect 34414 32450 34466 32462
rect 41022 32450 41074 32462
rect 36194 32398 36206 32450
rect 36258 32398 36270 32450
rect 44258 32398 44270 32450
rect 44322 32398 44334 32450
rect 45714 32398 45726 32450
rect 45778 32398 45790 32450
rect 34414 32386 34466 32398
rect 41022 32386 41074 32398
rect 2046 32338 2098 32350
rect 2046 32274 2098 32286
rect 2382 32338 2434 32350
rect 2382 32274 2434 32286
rect 2830 32338 2882 32350
rect 2830 32274 2882 32286
rect 9438 32338 9490 32350
rect 29262 32338 29314 32350
rect 16034 32286 16046 32338
rect 16098 32286 16110 32338
rect 26450 32286 26462 32338
rect 26514 32286 26526 32338
rect 9438 32274 9490 32286
rect 29262 32274 29314 32286
rect 33630 32338 33682 32350
rect 33630 32274 33682 32286
rect 46286 32338 46338 32350
rect 46286 32274 46338 32286
rect 46398 32338 46450 32350
rect 46398 32274 46450 32286
rect 48078 32338 48130 32350
rect 48078 32274 48130 32286
rect 1344 32170 49616 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 49616 32170
rect 1344 32084 49616 32118
rect 20190 32002 20242 32014
rect 20190 31938 20242 31950
rect 22542 32002 22594 32014
rect 22542 31938 22594 31950
rect 9214 31890 9266 31902
rect 2482 31838 2494 31890
rect 2546 31838 2558 31890
rect 4610 31838 4622 31890
rect 4674 31838 4686 31890
rect 6626 31838 6638 31890
rect 6690 31838 6702 31890
rect 8754 31838 8766 31890
rect 8818 31838 8830 31890
rect 9214 31826 9266 31838
rect 9774 31890 9826 31902
rect 28030 31890 28082 31902
rect 30382 31890 30434 31902
rect 35870 31890 35922 31902
rect 19618 31838 19630 31890
rect 19682 31838 19694 31890
rect 23874 31838 23886 31890
rect 23938 31838 23950 31890
rect 27458 31838 27470 31890
rect 27522 31838 27534 31890
rect 29922 31838 29934 31890
rect 29986 31838 29998 31890
rect 33058 31838 33070 31890
rect 33122 31838 33134 31890
rect 35186 31838 35198 31890
rect 35250 31838 35262 31890
rect 9774 31826 9826 31838
rect 28030 31826 28082 31838
rect 30382 31826 30434 31838
rect 35870 31826 35922 31838
rect 38446 31890 38498 31902
rect 38446 31826 38498 31838
rect 39118 31890 39170 31902
rect 39118 31826 39170 31838
rect 44830 31890 44882 31902
rect 44830 31826 44882 31838
rect 44942 31890 44994 31902
rect 47058 31838 47070 31890
rect 47122 31838 47134 31890
rect 49186 31838 49198 31890
rect 49250 31838 49262 31890
rect 44942 31826 44994 31838
rect 9998 31778 10050 31790
rect 1810 31726 1822 31778
rect 1874 31726 1886 31778
rect 5954 31726 5966 31778
rect 6018 31726 6030 31778
rect 9538 31726 9550 31778
rect 9602 31726 9614 31778
rect 9998 31714 10050 31726
rect 10446 31778 10498 31790
rect 10446 31714 10498 31726
rect 11006 31778 11058 31790
rect 20526 31778 20578 31790
rect 22430 31778 22482 31790
rect 13570 31726 13582 31778
rect 13634 31726 13646 31778
rect 19170 31726 19182 31778
rect 19234 31726 19246 31778
rect 19842 31726 19854 31778
rect 19906 31726 19918 31778
rect 21858 31726 21870 31778
rect 21922 31726 21934 31778
rect 11006 31714 11058 31726
rect 20526 31714 20578 31726
rect 22430 31714 22482 31726
rect 22990 31778 23042 31790
rect 30718 31778 30770 31790
rect 23426 31726 23438 31778
rect 23490 31726 23502 31778
rect 24546 31726 24558 31778
rect 24610 31726 24622 31778
rect 30034 31726 30046 31778
rect 30098 31726 30110 31778
rect 22990 31714 23042 31726
rect 30718 31714 30770 31726
rect 31390 31778 31442 31790
rect 35982 31778 36034 31790
rect 32386 31726 32398 31778
rect 32450 31726 32462 31778
rect 31390 31714 31442 31726
rect 35982 31714 36034 31726
rect 40014 31778 40066 31790
rect 40014 31714 40066 31726
rect 41134 31778 41186 31790
rect 45166 31778 45218 31790
rect 41682 31726 41694 31778
rect 41746 31726 41758 31778
rect 42242 31726 42254 31778
rect 42306 31726 42318 31778
rect 42914 31726 42926 31778
rect 42978 31726 42990 31778
rect 44258 31726 44270 31778
rect 44322 31726 44334 31778
rect 41134 31714 41186 31726
rect 45166 31714 45218 31726
rect 45726 31778 45778 31790
rect 46274 31726 46286 31778
rect 46338 31726 46350 31778
rect 45726 31714 45778 31726
rect 10110 31666 10162 31678
rect 10110 31602 10162 31614
rect 10670 31666 10722 31678
rect 20750 31666 20802 31678
rect 17490 31614 17502 31666
rect 17554 31614 17566 31666
rect 10670 31602 10722 31614
rect 20750 31602 20802 31614
rect 22094 31666 22146 31678
rect 22094 31602 22146 31614
rect 22542 31666 22594 31678
rect 27918 31666 27970 31678
rect 25330 31614 25342 31666
rect 25394 31614 25406 31666
rect 22542 31602 22594 31614
rect 27918 31602 27970 31614
rect 29374 31666 29426 31678
rect 29374 31602 29426 31614
rect 30942 31666 30994 31678
rect 30942 31602 30994 31614
rect 31278 31666 31330 31678
rect 31278 31602 31330 31614
rect 31614 31666 31666 31678
rect 31614 31602 31666 31614
rect 31838 31666 31890 31678
rect 31838 31602 31890 31614
rect 35534 31666 35586 31678
rect 35534 31602 35586 31614
rect 37326 31666 37378 31678
rect 37326 31602 37378 31614
rect 37774 31666 37826 31678
rect 37774 31602 37826 31614
rect 38782 31666 38834 31678
rect 45614 31666 45666 31678
rect 42466 31614 42478 31666
rect 42530 31614 42542 31666
rect 43026 31614 43038 31666
rect 43090 31614 43102 31666
rect 38782 31602 38834 31614
rect 45614 31602 45666 31614
rect 10782 31554 10834 31566
rect 10782 31490 10834 31502
rect 19406 31554 19458 31566
rect 19406 31490 19458 31502
rect 19630 31554 19682 31566
rect 19630 31490 19682 31502
rect 21534 31554 21586 31566
rect 21534 31490 21586 31502
rect 28478 31554 28530 31566
rect 28478 31490 28530 31502
rect 29598 31554 29650 31566
rect 29598 31490 29650 31502
rect 29822 31554 29874 31566
rect 29822 31490 29874 31502
rect 35758 31554 35810 31566
rect 35758 31490 35810 31502
rect 36094 31554 36146 31566
rect 36094 31490 36146 31502
rect 37214 31554 37266 31566
rect 37214 31490 37266 31502
rect 37438 31554 37490 31566
rect 37438 31490 37490 31502
rect 37550 31554 37602 31566
rect 37550 31490 37602 31502
rect 38222 31554 38274 31566
rect 38222 31490 38274 31502
rect 38334 31554 38386 31566
rect 38334 31490 38386 31502
rect 38558 31554 38610 31566
rect 38558 31490 38610 31502
rect 39678 31554 39730 31566
rect 39678 31490 39730 31502
rect 40574 31554 40626 31566
rect 40574 31490 40626 31502
rect 41246 31554 41298 31566
rect 41246 31490 41298 31502
rect 41358 31554 41410 31566
rect 41358 31490 41410 31502
rect 41470 31554 41522 31566
rect 45502 31554 45554 31566
rect 43138 31502 43150 31554
rect 43202 31502 43214 31554
rect 41470 31490 41522 31502
rect 45502 31490 45554 31502
rect 1344 31386 49616 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 49616 31386
rect 1344 31300 49616 31334
rect 2382 31218 2434 31230
rect 9886 31218 9938 31230
rect 9538 31166 9550 31218
rect 9602 31166 9614 31218
rect 2382 31154 2434 31166
rect 9886 31154 9938 31166
rect 16830 31218 16882 31230
rect 16830 31154 16882 31166
rect 17390 31218 17442 31230
rect 17390 31154 17442 31166
rect 17614 31218 17666 31230
rect 17614 31154 17666 31166
rect 18062 31218 18114 31230
rect 18062 31154 18114 31166
rect 18734 31218 18786 31230
rect 18734 31154 18786 31166
rect 19182 31218 19234 31230
rect 19182 31154 19234 31166
rect 20750 31218 20802 31230
rect 20750 31154 20802 31166
rect 25566 31218 25618 31230
rect 25566 31154 25618 31166
rect 26686 31218 26738 31230
rect 26686 31154 26738 31166
rect 27134 31218 27186 31230
rect 27134 31154 27186 31166
rect 30942 31218 30994 31230
rect 30942 31154 30994 31166
rect 31726 31218 31778 31230
rect 45614 31218 45666 31230
rect 34066 31166 34078 31218
rect 34130 31166 34142 31218
rect 34738 31166 34750 31218
rect 34802 31166 34814 31218
rect 43474 31166 43486 31218
rect 43538 31166 43550 31218
rect 31726 31154 31778 31166
rect 45614 31154 45666 31166
rect 45838 31218 45890 31230
rect 49086 31218 49138 31230
rect 48738 31166 48750 31218
rect 48802 31166 48814 31218
rect 45838 31154 45890 31166
rect 49086 31154 49138 31166
rect 4622 31106 4674 31118
rect 4622 31042 4674 31054
rect 6302 31106 6354 31118
rect 6302 31042 6354 31054
rect 6414 31106 6466 31118
rect 8206 31106 8258 31118
rect 6626 31054 6638 31106
rect 6690 31054 6702 31106
rect 6414 31042 6466 31054
rect 8206 31042 8258 31054
rect 8654 31106 8706 31118
rect 8654 31042 8706 31054
rect 16718 31106 16770 31118
rect 16718 31042 16770 31054
rect 17838 31106 17890 31118
rect 17838 31042 17890 31054
rect 18286 31106 18338 31118
rect 18286 31042 18338 31054
rect 18398 31106 18450 31118
rect 18398 31042 18450 31054
rect 20302 31106 20354 31118
rect 20302 31042 20354 31054
rect 25902 31106 25954 31118
rect 25902 31042 25954 31054
rect 30494 31106 30546 31118
rect 30494 31042 30546 31054
rect 31950 31106 32002 31118
rect 31950 31042 32002 31054
rect 34414 31106 34466 31118
rect 42590 31106 42642 31118
rect 37986 31054 37998 31106
rect 38050 31054 38062 31106
rect 34414 31042 34466 31054
rect 42590 31042 42642 31054
rect 44046 31106 44098 31118
rect 44046 31042 44098 31054
rect 46958 31106 47010 31118
rect 46958 31042 47010 31054
rect 2606 30994 2658 31006
rect 4510 30994 4562 31006
rect 6078 30994 6130 31006
rect 3490 30942 3502 30994
rect 3554 30942 3566 30994
rect 4050 30942 4062 30994
rect 4114 30942 4126 30994
rect 4834 30942 4846 30994
rect 4898 30942 4910 30994
rect 2606 30930 2658 30942
rect 4510 30930 4562 30942
rect 6078 30930 6130 30942
rect 7758 30994 7810 31006
rect 7758 30930 7810 30942
rect 7982 30994 8034 31006
rect 7982 30930 8034 30942
rect 8318 30994 8370 31006
rect 31502 30994 31554 31006
rect 13010 30942 13022 30994
rect 13074 30942 13086 30994
rect 13458 30942 13470 30994
rect 13522 30942 13534 30994
rect 20066 30942 20078 30994
rect 20130 30942 20142 30994
rect 21410 30942 21422 30994
rect 21474 30942 21486 30994
rect 8318 30930 8370 30942
rect 31502 30930 31554 30942
rect 31726 30994 31778 31006
rect 40910 30994 40962 31006
rect 33842 30942 33854 30994
rect 33906 30942 33918 30994
rect 35298 30942 35310 30994
rect 35362 30942 35374 30994
rect 31726 30930 31778 30942
rect 40910 30930 40962 30942
rect 41022 30994 41074 31006
rect 46062 30994 46114 31006
rect 41346 30942 41358 30994
rect 41410 30942 41422 30994
rect 43586 30942 43598 30994
rect 43650 30942 43662 30994
rect 41022 30930 41074 30942
rect 46062 30930 46114 30942
rect 46510 30994 46562 31006
rect 46510 30930 46562 30942
rect 47630 30994 47682 31006
rect 47630 30930 47682 30942
rect 47742 30994 47794 31006
rect 47742 30930 47794 30942
rect 47966 30994 48018 31006
rect 47966 30930 48018 30942
rect 48078 30994 48130 31006
rect 48078 30930 48130 30942
rect 7534 30882 7586 30894
rect 18846 30882 18898 30894
rect 2258 30830 2270 30882
rect 2322 30830 2334 30882
rect 6850 30830 6862 30882
rect 6914 30830 6926 30882
rect 10210 30830 10222 30882
rect 10274 30830 10286 30882
rect 12338 30830 12350 30882
rect 12402 30830 12414 30882
rect 14242 30830 14254 30882
rect 14306 30830 14318 30882
rect 16370 30830 16382 30882
rect 16434 30830 16446 30882
rect 7534 30818 7586 30830
rect 18846 30818 18898 30830
rect 19294 30882 19346 30894
rect 19294 30818 19346 30830
rect 20638 30882 20690 30894
rect 24670 30882 24722 30894
rect 22082 30830 22094 30882
rect 22146 30830 22158 30882
rect 24210 30830 24222 30882
rect 24274 30830 24286 30882
rect 20638 30818 20690 30830
rect 24670 30818 24722 30830
rect 27694 30882 27746 30894
rect 27694 30818 27746 30830
rect 28142 30882 28194 30894
rect 28142 30818 28194 30830
rect 28590 30882 28642 30894
rect 28590 30818 28642 30830
rect 29150 30882 29202 30894
rect 29150 30818 29202 30830
rect 29710 30882 29762 30894
rect 29710 30818 29762 30830
rect 30046 30882 30098 30894
rect 30046 30818 30098 30830
rect 32622 30882 32674 30894
rect 32622 30818 32674 30830
rect 33294 30882 33346 30894
rect 46286 30882 46338 30894
rect 45826 30830 45838 30882
rect 45890 30830 45902 30882
rect 33294 30818 33346 30830
rect 46286 30818 46338 30830
rect 47854 30882 47906 30894
rect 47854 30818 47906 30830
rect 2942 30770 2994 30782
rect 2942 30706 2994 30718
rect 3054 30770 3106 30782
rect 3054 30706 3106 30718
rect 3278 30770 3330 30782
rect 17726 30770 17778 30782
rect 7186 30718 7198 30770
rect 7250 30718 7262 30770
rect 3278 30706 3330 30718
rect 17726 30706 17778 30718
rect 29934 30770 29986 30782
rect 29934 30706 29986 30718
rect 33406 30770 33458 30782
rect 33406 30706 33458 30718
rect 46846 30770 46898 30782
rect 46846 30706 46898 30718
rect 1344 30602 49616 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 49616 30602
rect 1344 30516 49616 30550
rect 28142 30434 28194 30446
rect 28142 30370 28194 30382
rect 43486 30434 43538 30446
rect 43486 30370 43538 30382
rect 47406 30434 47458 30446
rect 47406 30370 47458 30382
rect 48862 30434 48914 30446
rect 48862 30370 48914 30382
rect 7086 30322 7138 30334
rect 43262 30322 43314 30334
rect 2482 30270 2494 30322
rect 2546 30270 2558 30322
rect 4610 30270 4622 30322
rect 4674 30270 4686 30322
rect 9202 30270 9214 30322
rect 9266 30270 9278 30322
rect 11330 30270 11342 30322
rect 11394 30270 11406 30322
rect 24098 30270 24110 30322
rect 24162 30270 24174 30322
rect 32050 30270 32062 30322
rect 32114 30270 32126 30322
rect 33058 30270 33070 30322
rect 33122 30270 33134 30322
rect 36978 30270 36990 30322
rect 37042 30270 37054 30322
rect 41570 30270 41582 30322
rect 41634 30270 41646 30322
rect 7086 30258 7138 30270
rect 43262 30258 43314 30270
rect 43934 30322 43986 30334
rect 48302 30322 48354 30334
rect 45042 30270 45054 30322
rect 45106 30270 45118 30322
rect 43934 30258 43986 30270
rect 48302 30258 48354 30270
rect 5966 30210 6018 30222
rect 6974 30210 7026 30222
rect 1810 30158 1822 30210
rect 1874 30158 1886 30210
rect 6402 30158 6414 30210
rect 6466 30158 6478 30210
rect 5966 30146 6018 30158
rect 6974 30146 7026 30158
rect 7198 30210 7250 30222
rect 13806 30210 13858 30222
rect 8082 30158 8094 30210
rect 8146 30158 8158 30210
rect 12114 30158 12126 30210
rect 12178 30158 12190 30210
rect 12674 30158 12686 30210
rect 12738 30158 12750 30210
rect 7198 30146 7250 30158
rect 13806 30146 13858 30158
rect 14478 30210 14530 30222
rect 14478 30146 14530 30158
rect 14702 30210 14754 30222
rect 21870 30210 21922 30222
rect 25566 30210 25618 30222
rect 27358 30210 27410 30222
rect 20626 30158 20638 30210
rect 20690 30158 20702 30210
rect 23762 30158 23774 30210
rect 23826 30158 23838 30210
rect 26226 30158 26238 30210
rect 26290 30158 26302 30210
rect 14702 30146 14754 30158
rect 21870 30146 21922 30158
rect 25566 30146 25618 30158
rect 27358 30146 27410 30158
rect 27694 30210 27746 30222
rect 27694 30146 27746 30158
rect 27918 30210 27970 30222
rect 28702 30210 28754 30222
rect 28354 30158 28366 30210
rect 28418 30158 28430 30210
rect 27918 30146 27970 30158
rect 28702 30146 28754 30158
rect 31054 30210 31106 30222
rect 36318 30210 36370 30222
rect 40686 30210 40738 30222
rect 42030 30210 42082 30222
rect 35186 30158 35198 30210
rect 35250 30158 35262 30210
rect 35970 30158 35982 30210
rect 36034 30158 36046 30210
rect 39778 30158 39790 30210
rect 39842 30158 39854 30210
rect 41122 30158 41134 30210
rect 41186 30158 41198 30210
rect 31054 30146 31106 30158
rect 36318 30146 36370 30158
rect 40686 30146 40738 30158
rect 42030 30146 42082 30158
rect 42254 30210 42306 30222
rect 42254 30146 42306 30158
rect 42814 30210 42866 30222
rect 42814 30146 42866 30158
rect 42926 30210 42978 30222
rect 42926 30146 42978 30158
rect 43710 30210 43762 30222
rect 45278 30210 45330 30222
rect 44818 30158 44830 30210
rect 44882 30158 44894 30210
rect 43710 30146 43762 30158
rect 45278 30146 45330 30158
rect 46062 30210 46114 30222
rect 46846 30210 46898 30222
rect 48190 30210 48242 30222
rect 46386 30158 46398 30210
rect 46450 30158 46462 30210
rect 47058 30158 47070 30210
rect 47122 30158 47134 30210
rect 47394 30158 47406 30210
rect 47458 30158 47470 30210
rect 46062 30146 46114 30158
rect 46846 30146 46898 30158
rect 48190 30146 48242 30158
rect 48414 30210 48466 30222
rect 48514 30158 48526 30210
rect 48578 30158 48590 30210
rect 48414 30146 48466 30158
rect 7422 30098 7474 30110
rect 12462 30098 12514 30110
rect 7858 30046 7870 30098
rect 7922 30046 7934 30098
rect 7422 30034 7474 30046
rect 12462 30034 12514 30046
rect 14142 30098 14194 30110
rect 22990 30098 23042 30110
rect 18386 30046 18398 30098
rect 18450 30046 18462 30098
rect 22642 30046 22654 30098
rect 22706 30046 22718 30098
rect 14142 30034 14194 30046
rect 22990 30034 23042 30046
rect 23326 30098 23378 30110
rect 23326 30034 23378 30046
rect 26798 30098 26850 30110
rect 26798 30034 26850 30046
rect 31614 30098 31666 30110
rect 31614 30034 31666 30046
rect 36430 30098 36482 30110
rect 40350 30098 40402 30110
rect 39106 30046 39118 30098
rect 39170 30046 39182 30098
rect 36430 30034 36482 30046
rect 40350 30034 40402 30046
rect 40462 30098 40514 30110
rect 40462 30034 40514 30046
rect 45054 30098 45106 30110
rect 45054 30034 45106 30046
rect 45502 30098 45554 30110
rect 45502 30034 45554 30046
rect 47742 30098 47794 30110
rect 47742 30034 47794 30046
rect 5630 29986 5682 29998
rect 5630 29922 5682 29934
rect 6638 29986 6690 29998
rect 21422 29986 21474 29998
rect 15026 29934 15038 29986
rect 15090 29934 15102 29986
rect 6638 29922 6690 29934
rect 21422 29922 21474 29934
rect 21646 29986 21698 29998
rect 21646 29922 21698 29934
rect 21758 29986 21810 29998
rect 21758 29922 21810 29934
rect 22430 29986 22482 29998
rect 22430 29922 22482 29934
rect 25006 29986 25058 29998
rect 28142 29986 28194 29998
rect 26450 29934 26462 29986
rect 26514 29934 26526 29986
rect 25006 29922 25058 29934
rect 28142 29922 28194 29934
rect 29374 29986 29426 29998
rect 29374 29922 29426 29934
rect 29710 29986 29762 29998
rect 29710 29922 29762 29934
rect 30270 29986 30322 29998
rect 30270 29922 30322 29934
rect 30718 29986 30770 29998
rect 30718 29922 30770 29934
rect 32510 29986 32562 29998
rect 32510 29922 32562 29934
rect 42702 29986 42754 29998
rect 42702 29922 42754 29934
rect 44382 29986 44434 29998
rect 44382 29922 44434 29934
rect 45726 29986 45778 29998
rect 45726 29922 45778 29934
rect 45950 29986 46002 29998
rect 45950 29922 46002 29934
rect 46622 29986 46674 29998
rect 46622 29922 46674 29934
rect 46734 29986 46786 29998
rect 46734 29922 46786 29934
rect 1344 29818 49616 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 49616 29818
rect 1344 29732 49616 29766
rect 3278 29650 3330 29662
rect 3278 29586 3330 29598
rect 5294 29650 5346 29662
rect 23886 29650 23938 29662
rect 7634 29598 7646 29650
rect 7698 29598 7710 29650
rect 12674 29598 12686 29650
rect 12738 29598 12750 29650
rect 5294 29586 5346 29598
rect 23886 29586 23938 29598
rect 24782 29650 24834 29662
rect 24782 29586 24834 29598
rect 34750 29650 34802 29662
rect 34750 29586 34802 29598
rect 34974 29650 35026 29662
rect 34974 29586 35026 29598
rect 35086 29650 35138 29662
rect 35086 29586 35138 29598
rect 36430 29650 36482 29662
rect 36430 29586 36482 29598
rect 36542 29650 36594 29662
rect 36542 29586 36594 29598
rect 40350 29650 40402 29662
rect 40350 29586 40402 29598
rect 41022 29650 41074 29662
rect 41022 29586 41074 29598
rect 41134 29650 41186 29662
rect 41134 29586 41186 29598
rect 41358 29650 41410 29662
rect 41358 29586 41410 29598
rect 42478 29650 42530 29662
rect 42478 29586 42530 29598
rect 42702 29650 42754 29662
rect 42702 29586 42754 29598
rect 48750 29650 48802 29662
rect 48750 29586 48802 29598
rect 8766 29538 8818 29550
rect 4834 29486 4846 29538
rect 4898 29486 4910 29538
rect 8306 29486 8318 29538
rect 8370 29486 8382 29538
rect 8766 29474 8818 29486
rect 10670 29538 10722 29550
rect 31726 29538 31778 29550
rect 34862 29538 34914 29550
rect 21410 29486 21422 29538
rect 21474 29486 21486 29538
rect 33394 29486 33406 29538
rect 33458 29486 33470 29538
rect 10670 29474 10722 29486
rect 31726 29474 31778 29486
rect 34862 29474 34914 29486
rect 36654 29538 36706 29550
rect 36654 29474 36706 29486
rect 42366 29538 42418 29550
rect 48862 29538 48914 29550
rect 46162 29486 46174 29538
rect 46226 29486 46238 29538
rect 42366 29474 42418 29486
rect 48862 29474 48914 29486
rect 3166 29426 3218 29438
rect 3166 29362 3218 29374
rect 3502 29426 3554 29438
rect 3502 29362 3554 29374
rect 3726 29426 3778 29438
rect 3726 29362 3778 29374
rect 3950 29426 4002 29438
rect 4622 29426 4674 29438
rect 4274 29374 4286 29426
rect 4338 29374 4350 29426
rect 3950 29362 4002 29374
rect 4622 29362 4674 29374
rect 4958 29426 5010 29438
rect 7310 29426 7362 29438
rect 5506 29374 5518 29426
rect 5570 29374 5582 29426
rect 4958 29362 5010 29374
rect 7310 29362 7362 29374
rect 7982 29426 8034 29438
rect 7982 29362 8034 29374
rect 11006 29426 11058 29438
rect 23998 29426 24050 29438
rect 33070 29426 33122 29438
rect 13906 29374 13918 29426
rect 13970 29374 13982 29426
rect 17490 29374 17502 29426
rect 17554 29374 17566 29426
rect 20738 29374 20750 29426
rect 20802 29374 20814 29426
rect 25218 29374 25230 29426
rect 25282 29374 25294 29426
rect 31378 29374 31390 29426
rect 31442 29374 31454 29426
rect 32162 29374 32174 29426
rect 32226 29374 32238 29426
rect 11006 29362 11058 29374
rect 23998 29362 24050 29374
rect 33070 29362 33122 29374
rect 33742 29426 33794 29438
rect 33742 29362 33794 29374
rect 33966 29426 34018 29438
rect 33966 29362 34018 29374
rect 34414 29426 34466 29438
rect 34414 29362 34466 29374
rect 35198 29426 35250 29438
rect 39342 29426 39394 29438
rect 35970 29374 35982 29426
rect 36034 29374 36046 29426
rect 36754 29374 36766 29426
rect 36818 29423 36830 29426
rect 36818 29377 37039 29423
rect 36818 29374 36830 29377
rect 35198 29362 35250 29374
rect 12126 29314 12178 29326
rect 30830 29314 30882 29326
rect 14690 29262 14702 29314
rect 14754 29262 14766 29314
rect 16818 29262 16830 29314
rect 16882 29262 16894 29314
rect 18162 29262 18174 29314
rect 18226 29262 18238 29314
rect 20290 29262 20302 29314
rect 20354 29262 20366 29314
rect 23538 29262 23550 29314
rect 23602 29262 23614 29314
rect 27458 29262 27470 29314
rect 27522 29262 27534 29314
rect 12126 29250 12178 29262
rect 30830 29250 30882 29262
rect 33854 29314 33906 29326
rect 36993 29314 37039 29377
rect 37650 29374 37662 29426
rect 37714 29374 37726 29426
rect 37874 29374 37886 29426
rect 37938 29374 37950 29426
rect 38322 29374 38334 29426
rect 38386 29374 38398 29426
rect 39342 29362 39394 29374
rect 39902 29426 39954 29438
rect 39902 29362 39954 29374
rect 40910 29426 40962 29438
rect 42914 29374 42926 29426
rect 42978 29374 42990 29426
rect 40910 29362 40962 29374
rect 41918 29314 41970 29326
rect 36978 29262 36990 29314
rect 37042 29262 37054 29314
rect 38434 29262 38446 29314
rect 38498 29262 38510 29314
rect 33854 29250 33906 29262
rect 41918 29250 41970 29262
rect 8654 29202 8706 29214
rect 8654 29138 8706 29150
rect 8990 29202 9042 29214
rect 8990 29138 9042 29150
rect 12350 29202 12402 29214
rect 12350 29138 12402 29150
rect 31054 29202 31106 29214
rect 31054 29138 31106 29150
rect 35646 29202 35698 29214
rect 35646 29138 35698 29150
rect 35982 29202 36034 29214
rect 41806 29202 41858 29214
rect 38546 29150 38558 29202
rect 38610 29150 38622 29202
rect 35982 29138 36034 29150
rect 41806 29138 41858 29150
rect 1344 29034 49616 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 49616 29034
rect 1344 28948 49616 28982
rect 5966 28866 6018 28878
rect 22542 28866 22594 28878
rect 21298 28814 21310 28866
rect 21362 28814 21374 28866
rect 5966 28802 6018 28814
rect 22542 28802 22594 28814
rect 35758 28866 35810 28878
rect 35758 28802 35810 28814
rect 43150 28866 43202 28878
rect 43150 28802 43202 28814
rect 44830 28866 44882 28878
rect 44830 28802 44882 28814
rect 45166 28866 45218 28878
rect 45166 28802 45218 28814
rect 47742 28866 47794 28878
rect 47742 28802 47794 28814
rect 4286 28754 4338 28766
rect 15150 28754 15202 28766
rect 47070 28754 47122 28766
rect 6402 28702 6414 28754
rect 6466 28702 6478 28754
rect 10434 28702 10446 28754
rect 10498 28702 10510 28754
rect 12562 28702 12574 28754
rect 12626 28702 12638 28754
rect 23090 28702 23102 28754
rect 23154 28702 23166 28754
rect 29138 28702 29150 28754
rect 29202 28702 29214 28754
rect 35298 28702 35310 28754
rect 35362 28702 35374 28754
rect 41570 28702 41582 28754
rect 41634 28702 41646 28754
rect 46498 28702 46510 28754
rect 46562 28702 46574 28754
rect 48738 28702 48750 28754
rect 48802 28702 48814 28754
rect 4286 28690 4338 28702
rect 15150 28690 15202 28702
rect 47070 28690 47122 28702
rect 3278 28642 3330 28654
rect 3278 28578 3330 28590
rect 3390 28642 3442 28654
rect 3390 28578 3442 28590
rect 3950 28642 4002 28654
rect 3950 28578 4002 28590
rect 4510 28642 4562 28654
rect 4510 28578 4562 28590
rect 4734 28642 4786 28654
rect 17054 28642 17106 28654
rect 19854 28642 19906 28654
rect 8530 28590 8542 28642
rect 8594 28590 8606 28642
rect 9202 28590 9214 28642
rect 9266 28590 9278 28642
rect 9650 28590 9662 28642
rect 9714 28590 9726 28642
rect 14690 28590 14702 28642
rect 14754 28590 14766 28642
rect 14914 28590 14926 28642
rect 14978 28590 14990 28642
rect 15698 28590 15710 28642
rect 15762 28590 15774 28642
rect 18722 28590 18734 28642
rect 18786 28590 18798 28642
rect 19394 28590 19406 28642
rect 19458 28590 19470 28642
rect 4734 28578 4786 28590
rect 17054 28578 17106 28590
rect 19854 28578 19906 28590
rect 20638 28642 20690 28654
rect 20638 28578 20690 28590
rect 21758 28642 21810 28654
rect 21758 28578 21810 28590
rect 21870 28642 21922 28654
rect 21870 28578 21922 28590
rect 21982 28642 22034 28654
rect 27694 28642 27746 28654
rect 23202 28590 23214 28642
rect 23266 28590 23278 28642
rect 26338 28590 26350 28642
rect 26402 28590 26414 28642
rect 21982 28578 22034 28590
rect 27694 28578 27746 28590
rect 28590 28642 28642 28654
rect 35870 28642 35922 28654
rect 48414 28642 48466 28654
rect 31266 28590 31278 28642
rect 31330 28590 31342 28642
rect 32050 28590 32062 28642
rect 32114 28590 32126 28642
rect 32386 28590 32398 28642
rect 32450 28590 32462 28642
rect 36082 28590 36094 28642
rect 36146 28590 36158 28642
rect 37314 28590 37326 28642
rect 37378 28590 37390 28642
rect 38658 28590 38670 28642
rect 38722 28590 38734 28642
rect 40450 28590 40462 28642
rect 40514 28590 40526 28642
rect 42578 28590 42590 28642
rect 42642 28590 42654 28642
rect 43026 28590 43038 28642
rect 43090 28590 43102 28642
rect 45154 28590 45166 28642
rect 45218 28590 45230 28642
rect 45490 28590 45502 28642
rect 45554 28590 45566 28642
rect 46050 28590 46062 28642
rect 46114 28590 46126 28642
rect 48066 28590 48078 28642
rect 48130 28590 48142 28642
rect 28590 28578 28642 28590
rect 35870 28578 35922 28590
rect 48414 28578 48466 28590
rect 49198 28642 49250 28654
rect 49198 28578 49250 28590
rect 3502 28530 3554 28542
rect 3502 28466 3554 28478
rect 4174 28530 4226 28542
rect 4174 28466 4226 28478
rect 5854 28530 5906 28542
rect 5854 28466 5906 28478
rect 5966 28530 6018 28542
rect 5966 28466 6018 28478
rect 15486 28530 15538 28542
rect 15486 28466 15538 28478
rect 16718 28530 16770 28542
rect 16718 28466 16770 28478
rect 17726 28530 17778 28542
rect 17726 28466 17778 28478
rect 17838 28530 17890 28542
rect 22430 28530 22482 28542
rect 18274 28478 18286 28530
rect 18338 28478 18350 28530
rect 20178 28478 20190 28530
rect 20242 28478 20254 28530
rect 17838 28466 17890 28478
rect 22430 28466 22482 28478
rect 22542 28530 22594 28542
rect 26798 28530 26850 28542
rect 24658 28478 24670 28530
rect 24722 28478 24734 28530
rect 25778 28478 25790 28530
rect 25842 28478 25854 28530
rect 22542 28466 22594 28478
rect 26798 28466 26850 28478
rect 27358 28530 27410 28542
rect 27358 28466 27410 28478
rect 28478 28530 28530 28542
rect 44046 28530 44098 28542
rect 46958 28530 47010 28542
rect 33170 28478 33182 28530
rect 33234 28478 33246 28530
rect 36978 28478 36990 28530
rect 37042 28478 37054 28530
rect 39106 28478 39118 28530
rect 39170 28478 39182 28530
rect 40338 28478 40350 28530
rect 40402 28478 40414 28530
rect 43138 28478 43150 28530
rect 43202 28478 43214 28530
rect 46162 28478 46174 28530
rect 46226 28478 46238 28530
rect 28478 28466 28530 28478
rect 44046 28466 44098 28478
rect 46958 28466 47010 28478
rect 47182 28530 47234 28542
rect 47182 28466 47234 28478
rect 47406 28530 47458 28542
rect 47406 28466 47458 28478
rect 47854 28530 47906 28542
rect 47854 28466 47906 28478
rect 16606 28418 16658 28430
rect 16606 28354 16658 28366
rect 17166 28418 17218 28430
rect 17166 28354 17218 28366
rect 18062 28418 18114 28430
rect 26910 28418 26962 28430
rect 18498 28366 18510 28418
rect 18562 28366 18574 28418
rect 18062 28354 18114 28366
rect 26910 28354 26962 28366
rect 27582 28418 27634 28430
rect 27582 28354 27634 28366
rect 27806 28418 27858 28430
rect 27806 28354 27858 28366
rect 27918 28418 27970 28430
rect 27918 28354 27970 28366
rect 44158 28418 44210 28430
rect 44158 28354 44210 28366
rect 1344 28250 49616 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 49616 28250
rect 1344 28164 49616 28198
rect 16270 28082 16322 28094
rect 6402 28030 6414 28082
rect 6466 28030 6478 28082
rect 11106 28030 11118 28082
rect 11170 28030 11182 28082
rect 16270 28018 16322 28030
rect 16382 28082 16434 28094
rect 16382 28018 16434 28030
rect 18398 28082 18450 28094
rect 18398 28018 18450 28030
rect 19630 28082 19682 28094
rect 19630 28018 19682 28030
rect 20750 28082 20802 28094
rect 20750 28018 20802 28030
rect 21086 28082 21138 28094
rect 21086 28018 21138 28030
rect 26014 28082 26066 28094
rect 26014 28018 26066 28030
rect 26574 28082 26626 28094
rect 26574 28018 26626 28030
rect 26686 28082 26738 28094
rect 26686 28018 26738 28030
rect 26910 28082 26962 28094
rect 26910 28018 26962 28030
rect 31726 28082 31778 28094
rect 31726 28018 31778 28030
rect 35758 28082 35810 28094
rect 35758 28018 35810 28030
rect 48078 28082 48130 28094
rect 48078 28018 48130 28030
rect 8206 27970 8258 27982
rect 4946 27918 4958 27970
rect 5010 27918 5022 27970
rect 6514 27918 6526 27970
rect 6578 27918 6590 27970
rect 7410 27918 7422 27970
rect 7474 27918 7486 27970
rect 7746 27918 7758 27970
rect 7810 27918 7822 27970
rect 8206 27906 8258 27918
rect 13806 27970 13858 27982
rect 13806 27906 13858 27918
rect 14030 27970 14082 27982
rect 14030 27906 14082 27918
rect 16606 27970 16658 27982
rect 16606 27906 16658 27918
rect 17502 27970 17554 27982
rect 25342 27970 25394 27982
rect 32062 27970 32114 27982
rect 18610 27918 18622 27970
rect 18674 27918 18686 27970
rect 28130 27918 28142 27970
rect 28194 27918 28206 27970
rect 17502 27906 17554 27918
rect 25342 27906 25394 27918
rect 32062 27906 32114 27918
rect 33518 27970 33570 27982
rect 33518 27906 33570 27918
rect 33630 27970 33682 27982
rect 33630 27906 33682 27918
rect 33854 27970 33906 27982
rect 33854 27906 33906 27918
rect 34078 27970 34130 27982
rect 34078 27906 34130 27918
rect 5518 27858 5570 27870
rect 7086 27858 7138 27870
rect 1810 27806 1822 27858
rect 1874 27806 1886 27858
rect 5954 27806 5966 27858
rect 6018 27806 6030 27858
rect 5518 27794 5570 27806
rect 7086 27794 7138 27806
rect 8654 27858 8706 27870
rect 8654 27794 8706 27806
rect 11678 27858 11730 27870
rect 16046 27858 16098 27870
rect 12562 27806 12574 27858
rect 12626 27806 12638 27858
rect 15026 27806 15038 27858
rect 15090 27806 15102 27858
rect 15250 27806 15262 27858
rect 15314 27806 15326 27858
rect 11678 27794 11730 27806
rect 16046 27794 16098 27806
rect 16158 27858 16210 27870
rect 16158 27794 16210 27806
rect 17390 27858 17442 27870
rect 17390 27794 17442 27806
rect 17950 27858 18002 27870
rect 17950 27794 18002 27806
rect 18174 27858 18226 27870
rect 18174 27794 18226 27806
rect 18958 27858 19010 27870
rect 18958 27794 19010 27806
rect 19182 27858 19234 27870
rect 19182 27794 19234 27806
rect 19406 27858 19458 27870
rect 19406 27794 19458 27806
rect 19854 27858 19906 27870
rect 19854 27794 19906 27806
rect 21422 27858 21474 27870
rect 26798 27858 26850 27870
rect 31166 27858 31218 27870
rect 34414 27858 34466 27870
rect 38446 27858 38498 27870
rect 24658 27806 24670 27858
rect 24722 27806 24734 27858
rect 26338 27806 26350 27858
rect 26402 27806 26414 27858
rect 27458 27806 27470 27858
rect 27522 27806 27534 27858
rect 32274 27806 32286 27858
rect 32338 27806 32350 27858
rect 32498 27806 32510 27858
rect 32562 27806 32574 27858
rect 34626 27806 34638 27858
rect 34690 27806 34702 27858
rect 35074 27806 35086 27858
rect 35138 27806 35150 27858
rect 36530 27806 36542 27858
rect 36594 27855 36606 27858
rect 36866 27855 36878 27858
rect 36594 27809 36878 27855
rect 36594 27806 36606 27809
rect 36866 27806 36878 27809
rect 36930 27806 36942 27858
rect 38210 27806 38222 27858
rect 38274 27806 38286 27858
rect 21422 27794 21474 27806
rect 26798 27794 26850 27806
rect 31166 27794 31218 27806
rect 34414 27794 34466 27806
rect 38446 27794 38498 27806
rect 38782 27858 38834 27870
rect 46846 27858 46898 27870
rect 39106 27806 39118 27858
rect 39170 27806 39182 27858
rect 44706 27806 44718 27858
rect 44770 27806 44782 27858
rect 38782 27794 38834 27806
rect 46846 27794 46898 27806
rect 7870 27746 7922 27758
rect 2482 27694 2494 27746
rect 2546 27694 2558 27746
rect 4610 27694 4622 27746
rect 4674 27694 4686 27746
rect 7870 27682 7922 27694
rect 8318 27746 8370 27758
rect 8318 27682 8370 27694
rect 11454 27746 11506 27758
rect 11454 27682 11506 27694
rect 12014 27746 12066 27758
rect 19742 27746 19794 27758
rect 25230 27746 25282 27758
rect 30718 27746 30770 27758
rect 33070 27746 33122 27758
rect 12786 27694 12798 27746
rect 12850 27694 12862 27746
rect 13682 27694 13694 27746
rect 13746 27694 13758 27746
rect 14914 27694 14926 27746
rect 14978 27694 14990 27746
rect 21746 27694 21758 27746
rect 21810 27694 21822 27746
rect 23874 27694 23886 27746
rect 23938 27694 23950 27746
rect 30258 27694 30270 27746
rect 30322 27694 30334 27746
rect 32162 27694 32174 27746
rect 32226 27694 32238 27746
rect 12014 27682 12066 27694
rect 19742 27682 19794 27694
rect 25230 27682 25282 27694
rect 30718 27682 30770 27694
rect 33070 27682 33122 27694
rect 36318 27746 36370 27758
rect 47070 27746 47122 27758
rect 44146 27694 44158 27746
rect 44210 27694 44222 27746
rect 36318 27682 36370 27694
rect 47070 27682 47122 27694
rect 47630 27746 47682 27758
rect 47630 27682 47682 27694
rect 48190 27746 48242 27758
rect 48190 27682 48242 27694
rect 48862 27746 48914 27758
rect 48862 27682 48914 27694
rect 6862 27634 6914 27646
rect 6862 27570 6914 27582
rect 8542 27634 8594 27646
rect 17502 27634 17554 27646
rect 14466 27582 14478 27634
rect 14530 27582 14542 27634
rect 8542 27570 8594 27582
rect 17502 27570 17554 27582
rect 18398 27634 18450 27646
rect 18398 27570 18450 27582
rect 33182 27634 33234 27646
rect 46510 27634 46562 27646
rect 37538 27582 37550 27634
rect 37602 27582 37614 27634
rect 33182 27570 33234 27582
rect 46510 27570 46562 27582
rect 47518 27634 47570 27646
rect 47518 27570 47570 27582
rect 48750 27634 48802 27646
rect 48750 27570 48802 27582
rect 1344 27466 49616 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 49616 27466
rect 1344 27380 49616 27414
rect 2494 27298 2546 27310
rect 6414 27298 6466 27310
rect 4498 27246 4510 27298
rect 4562 27246 4574 27298
rect 6066 27246 6078 27298
rect 6130 27246 6142 27298
rect 2494 27234 2546 27246
rect 6414 27234 6466 27246
rect 15934 27298 15986 27310
rect 15934 27234 15986 27246
rect 17390 27298 17442 27310
rect 17390 27234 17442 27246
rect 17614 27298 17666 27310
rect 17614 27234 17666 27246
rect 44942 27298 44994 27310
rect 44942 27234 44994 27246
rect 2606 27186 2658 27198
rect 2606 27122 2658 27134
rect 5070 27186 5122 27198
rect 5070 27122 5122 27134
rect 6638 27186 6690 27198
rect 6638 27122 6690 27134
rect 12798 27186 12850 27198
rect 12798 27122 12850 27134
rect 13470 27186 13522 27198
rect 15822 27186 15874 27198
rect 14354 27134 14366 27186
rect 14418 27134 14430 27186
rect 15362 27134 15374 27186
rect 15426 27134 15438 27186
rect 13470 27122 13522 27134
rect 15822 27122 15874 27134
rect 17166 27186 17218 27198
rect 17166 27122 17218 27134
rect 18622 27186 18674 27198
rect 18622 27122 18674 27134
rect 19406 27186 19458 27198
rect 19406 27122 19458 27134
rect 19854 27186 19906 27198
rect 29486 27186 29538 27198
rect 21298 27134 21310 27186
rect 21362 27134 21374 27186
rect 24882 27134 24894 27186
rect 24946 27134 24958 27186
rect 27010 27134 27022 27186
rect 27074 27134 27086 27186
rect 19854 27122 19906 27134
rect 29486 27122 29538 27134
rect 38334 27186 38386 27198
rect 42814 27186 42866 27198
rect 45390 27186 45442 27198
rect 40002 27134 40014 27186
rect 40066 27134 40078 27186
rect 42130 27134 42142 27186
rect 42194 27134 42206 27186
rect 44034 27134 44046 27186
rect 44098 27134 44110 27186
rect 38334 27122 38386 27134
rect 42814 27122 42866 27134
rect 45390 27122 45442 27134
rect 45838 27186 45890 27198
rect 49186 27134 49198 27186
rect 49250 27134 49262 27186
rect 45838 27122 45890 27134
rect 3278 27074 3330 27086
rect 3278 27010 3330 27022
rect 3726 27074 3778 27086
rect 3726 27010 3778 27022
rect 3950 27074 4002 27086
rect 4846 27074 4898 27086
rect 15262 27074 15314 27086
rect 4162 27022 4174 27074
rect 4226 27022 4238 27074
rect 12226 27022 12238 27074
rect 12290 27022 12302 27074
rect 13906 27022 13918 27074
rect 13970 27022 13982 27074
rect 14802 27022 14814 27074
rect 14866 27022 14878 27074
rect 3950 27010 4002 27022
rect 4846 27010 4898 27022
rect 15262 27010 15314 27022
rect 16606 27074 16658 27086
rect 18734 27074 18786 27086
rect 19294 27074 19346 27086
rect 18274 27022 18286 27074
rect 18338 27022 18350 27074
rect 18946 27022 18958 27074
rect 19010 27022 19022 27074
rect 16606 27010 16658 27022
rect 18734 27010 18786 27022
rect 19294 27010 19346 27022
rect 20750 27074 20802 27086
rect 36990 27074 37042 27086
rect 24210 27022 24222 27074
rect 24274 27022 24286 27074
rect 27794 27022 27806 27074
rect 27858 27022 27870 27074
rect 29138 27022 29150 27074
rect 29202 27022 29214 27074
rect 36194 27022 36206 27074
rect 36258 27022 36270 27074
rect 20750 27010 20802 27022
rect 36990 27010 37042 27022
rect 37326 27074 37378 27086
rect 39330 27022 39342 27074
rect 39394 27022 39406 27074
rect 42466 27022 42478 27074
rect 42530 27022 42542 27074
rect 43474 27022 43486 27074
rect 43538 27022 43550 27074
rect 46274 27022 46286 27074
rect 46338 27022 46350 27074
rect 37326 27010 37378 27022
rect 3614 26962 3666 26974
rect 16382 26962 16434 26974
rect 2930 26910 2942 26962
rect 2994 26910 3006 26962
rect 8418 26910 8430 26962
rect 8482 26910 8494 26962
rect 3614 26898 3666 26910
rect 16382 26898 16434 26910
rect 16830 26962 16882 26974
rect 16830 26898 16882 26910
rect 18510 26962 18562 26974
rect 29374 26962 29426 26974
rect 20402 26910 20414 26962
rect 20466 26910 20478 26962
rect 23426 26910 23438 26962
rect 23490 26910 23502 26962
rect 18510 26898 18562 26910
rect 29374 26898 29426 26910
rect 29598 26962 29650 26974
rect 29598 26898 29650 26910
rect 30382 26962 30434 26974
rect 37102 26962 37154 26974
rect 32386 26910 32398 26962
rect 32450 26910 32462 26962
rect 30382 26898 30434 26910
rect 37102 26898 37154 26910
rect 37662 26962 37714 26974
rect 43710 26962 43762 26974
rect 37986 26910 37998 26962
rect 38050 26910 38062 26962
rect 37662 26898 37714 26910
rect 43710 26898 43762 26910
rect 43934 26962 43986 26974
rect 43934 26898 43986 26910
rect 44830 26962 44882 26974
rect 47058 26910 47070 26962
rect 47122 26910 47134 26962
rect 44830 26898 44882 26910
rect 15038 26850 15090 26862
rect 15038 26786 15090 26798
rect 15374 26850 15426 26862
rect 15374 26786 15426 26798
rect 16718 26850 16770 26862
rect 16718 26786 16770 26798
rect 18062 26850 18114 26862
rect 18062 26786 18114 26798
rect 28254 26850 28306 26862
rect 28254 26786 28306 26798
rect 29710 26850 29762 26862
rect 29710 26786 29762 26798
rect 30718 26850 30770 26862
rect 30718 26786 30770 26798
rect 38894 26850 38946 26862
rect 38894 26786 38946 26798
rect 42702 26850 42754 26862
rect 42702 26786 42754 26798
rect 42926 26850 42978 26862
rect 42926 26786 42978 26798
rect 43038 26850 43090 26862
rect 43038 26786 43090 26798
rect 44046 26850 44098 26862
rect 44046 26786 44098 26798
rect 1344 26682 49616 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 49616 26682
rect 1344 26596 49616 26630
rect 5182 26514 5234 26526
rect 16494 26514 16546 26526
rect 14914 26462 14926 26514
rect 14978 26462 14990 26514
rect 5182 26450 5234 26462
rect 16494 26450 16546 26462
rect 17614 26514 17666 26526
rect 17614 26450 17666 26462
rect 19742 26514 19794 26526
rect 19742 26450 19794 26462
rect 20974 26514 21026 26526
rect 20974 26450 21026 26462
rect 21422 26514 21474 26526
rect 30270 26514 30322 26526
rect 28466 26462 28478 26514
rect 28530 26462 28542 26514
rect 21422 26450 21474 26462
rect 30270 26450 30322 26462
rect 31614 26514 31666 26526
rect 31614 26450 31666 26462
rect 32062 26514 32114 26526
rect 32062 26450 32114 26462
rect 32510 26514 32562 26526
rect 46510 26514 46562 26526
rect 46050 26462 46062 26514
rect 46114 26462 46126 26514
rect 32510 26450 32562 26462
rect 46510 26450 46562 26462
rect 47630 26514 47682 26526
rect 47630 26450 47682 26462
rect 47742 26514 47794 26526
rect 47742 26450 47794 26462
rect 14030 26402 14082 26414
rect 2482 26350 2494 26402
rect 2546 26350 2558 26402
rect 13234 26350 13246 26402
rect 13298 26350 13310 26402
rect 13570 26350 13582 26402
rect 13634 26350 13646 26402
rect 14030 26338 14082 26350
rect 15710 26402 15762 26414
rect 15710 26338 15762 26350
rect 17390 26402 17442 26414
rect 17390 26338 17442 26350
rect 17838 26402 17890 26414
rect 30158 26402 30210 26414
rect 29138 26350 29150 26402
rect 29202 26350 29214 26402
rect 17838 26338 17890 26350
rect 30158 26338 30210 26350
rect 30494 26402 30546 26414
rect 30494 26338 30546 26350
rect 39790 26402 39842 26414
rect 46622 26402 46674 26414
rect 44594 26350 44606 26402
rect 44658 26350 44670 26402
rect 39790 26338 39842 26350
rect 46622 26338 46674 26350
rect 46846 26402 46898 26414
rect 46846 26338 46898 26350
rect 48078 26402 48130 26414
rect 48078 26338 48130 26350
rect 13694 26290 13746 26302
rect 1810 26238 1822 26290
rect 1874 26238 1886 26290
rect 4946 26238 4958 26290
rect 5010 26238 5022 26290
rect 6178 26238 6190 26290
rect 6242 26238 6254 26290
rect 9538 26238 9550 26290
rect 9602 26238 9614 26290
rect 13122 26238 13134 26290
rect 13186 26238 13198 26290
rect 13694 26226 13746 26238
rect 14254 26290 14306 26302
rect 14254 26226 14306 26238
rect 14590 26290 14642 26302
rect 15822 26290 15874 26302
rect 16382 26290 16434 26302
rect 15138 26238 15150 26290
rect 15202 26238 15214 26290
rect 16146 26238 16158 26290
rect 16210 26238 16222 26290
rect 14590 26226 14642 26238
rect 15822 26226 15874 26238
rect 16382 26226 16434 26238
rect 16606 26290 16658 26302
rect 18398 26290 18450 26302
rect 28814 26290 28866 26302
rect 16818 26238 16830 26290
rect 16882 26238 16894 26290
rect 18050 26238 18062 26290
rect 18114 26238 18126 26290
rect 24658 26238 24670 26290
rect 24722 26238 24734 26290
rect 28130 26238 28142 26290
rect 28194 26238 28206 26290
rect 16606 26226 16658 26238
rect 18398 26226 18450 26238
rect 28814 26226 28866 26238
rect 29486 26290 29538 26302
rect 29486 26226 29538 26238
rect 30606 26290 30658 26302
rect 45726 26290 45778 26302
rect 47518 26290 47570 26302
rect 35970 26238 35982 26290
rect 36034 26238 36046 26290
rect 39218 26238 39230 26290
rect 39282 26238 39294 26290
rect 42130 26238 42142 26290
rect 42194 26238 42206 26290
rect 45378 26238 45390 26290
rect 45442 26238 45454 26290
rect 47058 26238 47070 26290
rect 47122 26238 47134 26290
rect 30606 26226 30658 26238
rect 45726 26226 45778 26238
rect 47518 26226 47570 26238
rect 47854 26290 47906 26302
rect 47854 26226 47906 26238
rect 14142 26178 14194 26190
rect 4610 26126 4622 26178
rect 4674 26126 4686 26178
rect 6850 26126 6862 26178
rect 6914 26126 6926 26178
rect 8978 26126 8990 26178
rect 9042 26126 9054 26178
rect 10322 26126 10334 26178
rect 10386 26126 10398 26178
rect 12450 26126 12462 26178
rect 12514 26126 12526 26178
rect 14142 26114 14194 26126
rect 17726 26178 17778 26190
rect 17726 26114 17778 26126
rect 18510 26178 18562 26190
rect 18510 26114 18562 26126
rect 19294 26178 19346 26190
rect 19294 26114 19346 26126
rect 21310 26178 21362 26190
rect 31054 26178 31106 26190
rect 39678 26178 39730 26190
rect 21746 26126 21758 26178
rect 21810 26126 21822 26178
rect 23874 26126 23886 26178
rect 23938 26126 23950 26178
rect 25218 26126 25230 26178
rect 25282 26126 25294 26178
rect 27346 26126 27358 26178
rect 27410 26126 27422 26178
rect 33058 26126 33070 26178
rect 33122 26126 33134 26178
rect 35186 26126 35198 26178
rect 35250 26126 35262 26178
rect 36306 26126 36318 26178
rect 36370 26126 36382 26178
rect 38434 26126 38446 26178
rect 38498 26126 38510 26178
rect 21310 26114 21362 26126
rect 31054 26114 31106 26126
rect 39678 26114 39730 26126
rect 40350 26178 40402 26190
rect 46734 26178 46786 26190
rect 41458 26126 41470 26178
rect 41522 26126 41534 26178
rect 42466 26126 42478 26178
rect 42530 26126 42542 26178
rect 40350 26114 40402 26126
rect 46734 26114 46786 26126
rect 48862 26178 48914 26190
rect 48862 26114 48914 26126
rect 5294 26066 5346 26078
rect 5294 26002 5346 26014
rect 12686 26066 12738 26078
rect 12686 26002 12738 26014
rect 39566 26066 39618 26078
rect 39566 26002 39618 26014
rect 48750 26066 48802 26078
rect 48750 26002 48802 26014
rect 1344 25898 49616 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 49616 25898
rect 1344 25812 49616 25846
rect 4174 25730 4226 25742
rect 4174 25666 4226 25678
rect 4846 25730 4898 25742
rect 4846 25666 4898 25678
rect 6078 25730 6130 25742
rect 6078 25666 6130 25678
rect 6750 25730 6802 25742
rect 6750 25666 6802 25678
rect 7198 25730 7250 25742
rect 7198 25666 7250 25678
rect 14478 25730 14530 25742
rect 14478 25666 14530 25678
rect 14926 25730 14978 25742
rect 14926 25666 14978 25678
rect 15374 25730 15426 25742
rect 15374 25666 15426 25678
rect 23102 25730 23154 25742
rect 23102 25666 23154 25678
rect 26798 25730 26850 25742
rect 26798 25666 26850 25678
rect 32734 25730 32786 25742
rect 32734 25666 32786 25678
rect 33070 25730 33122 25742
rect 33070 25666 33122 25678
rect 5854 25618 5906 25630
rect 5854 25554 5906 25566
rect 6862 25618 6914 25630
rect 6862 25554 6914 25566
rect 14366 25618 14418 25630
rect 14366 25554 14418 25566
rect 15262 25618 15314 25630
rect 25902 25618 25954 25630
rect 33518 25618 33570 25630
rect 17938 25566 17950 25618
rect 18002 25566 18014 25618
rect 22082 25566 22094 25618
rect 22146 25566 22158 25618
rect 32050 25566 32062 25618
rect 32114 25566 32126 25618
rect 15262 25554 15314 25566
rect 25902 25554 25954 25566
rect 33518 25554 33570 25566
rect 35534 25618 35586 25630
rect 35534 25554 35586 25566
rect 36990 25618 37042 25630
rect 36990 25554 37042 25566
rect 37998 25618 38050 25630
rect 46946 25566 46958 25618
rect 47010 25566 47022 25618
rect 49074 25566 49086 25618
rect 49138 25566 49150 25618
rect 37998 25554 38050 25566
rect 5070 25506 5122 25518
rect 5070 25442 5122 25454
rect 7086 25506 7138 25518
rect 7086 25442 7138 25454
rect 7982 25506 8034 25518
rect 7982 25442 8034 25454
rect 8430 25506 8482 25518
rect 9774 25506 9826 25518
rect 10782 25506 10834 25518
rect 8642 25454 8654 25506
rect 8706 25454 8718 25506
rect 10434 25454 10446 25506
rect 10498 25454 10510 25506
rect 8430 25442 8482 25454
rect 9774 25442 9826 25454
rect 10782 25442 10834 25454
rect 11006 25506 11058 25518
rect 11006 25442 11058 25454
rect 12238 25506 12290 25518
rect 16270 25506 16322 25518
rect 12450 25454 12462 25506
rect 12514 25454 12526 25506
rect 12238 25442 12290 25454
rect 16270 25442 16322 25454
rect 16718 25506 16770 25518
rect 16718 25442 16770 25454
rect 16942 25506 16994 25518
rect 19630 25506 19682 25518
rect 17490 25454 17502 25506
rect 17554 25454 17566 25506
rect 18722 25454 18734 25506
rect 18786 25454 18798 25506
rect 16942 25442 16994 25454
rect 19630 25442 19682 25454
rect 20414 25506 20466 25518
rect 20414 25442 20466 25454
rect 20526 25506 20578 25518
rect 22206 25506 22258 25518
rect 20738 25454 20750 25506
rect 20802 25454 20814 25506
rect 21970 25454 21982 25506
rect 22034 25454 22046 25506
rect 20526 25442 20578 25454
rect 22206 25442 22258 25454
rect 22542 25506 22594 25518
rect 23886 25506 23938 25518
rect 23426 25454 23438 25506
rect 23490 25454 23502 25506
rect 22542 25442 22594 25454
rect 23886 25442 23938 25454
rect 23998 25506 24050 25518
rect 23998 25442 24050 25454
rect 24782 25506 24834 25518
rect 24782 25442 24834 25454
rect 25454 25506 25506 25518
rect 27582 25506 27634 25518
rect 27346 25454 27358 25506
rect 27410 25454 27422 25506
rect 25454 25442 25506 25454
rect 27582 25442 27634 25454
rect 27806 25506 27858 25518
rect 33742 25506 33794 25518
rect 28018 25454 28030 25506
rect 28082 25454 28094 25506
rect 29250 25454 29262 25506
rect 29314 25454 29326 25506
rect 27806 25442 27858 25454
rect 33742 25442 33794 25454
rect 33966 25506 34018 25518
rect 34526 25506 34578 25518
rect 34290 25454 34302 25506
rect 34354 25454 34366 25506
rect 33966 25442 34018 25454
rect 34526 25442 34578 25454
rect 34638 25506 34690 25518
rect 34638 25442 34690 25454
rect 35646 25506 35698 25518
rect 35646 25442 35698 25454
rect 35870 25506 35922 25518
rect 35870 25442 35922 25454
rect 36318 25506 36370 25518
rect 36318 25442 36370 25454
rect 37214 25506 37266 25518
rect 37214 25442 37266 25454
rect 37774 25506 37826 25518
rect 37774 25442 37826 25454
rect 38334 25506 38386 25518
rect 44270 25506 44322 25518
rect 40338 25454 40350 25506
rect 40402 25454 40414 25506
rect 40786 25454 40798 25506
rect 40850 25454 40862 25506
rect 42914 25454 42926 25506
rect 42978 25454 42990 25506
rect 38334 25442 38386 25454
rect 44270 25442 44322 25454
rect 45278 25506 45330 25518
rect 45278 25442 45330 25454
rect 45502 25506 45554 25518
rect 46274 25454 46286 25506
rect 46338 25454 46350 25506
rect 45502 25442 45554 25454
rect 8318 25394 8370 25406
rect 6402 25342 6414 25394
rect 6466 25342 6478 25394
rect 7634 25342 7646 25394
rect 7698 25342 7710 25394
rect 8318 25330 8370 25342
rect 10110 25394 10162 25406
rect 10110 25330 10162 25342
rect 12126 25394 12178 25406
rect 12126 25330 12178 25342
rect 14814 25394 14866 25406
rect 14814 25330 14866 25342
rect 16046 25394 16098 25406
rect 16046 25330 16098 25342
rect 18174 25394 18226 25406
rect 18174 25330 18226 25342
rect 18286 25394 18338 25406
rect 18286 25330 18338 25342
rect 20078 25394 20130 25406
rect 20078 25330 20130 25342
rect 21310 25394 21362 25406
rect 21310 25330 21362 25342
rect 22990 25394 23042 25406
rect 22990 25330 23042 25342
rect 23774 25394 23826 25406
rect 26686 25394 26738 25406
rect 25106 25342 25118 25394
rect 25170 25342 25182 25394
rect 23774 25330 23826 25342
rect 26686 25330 26738 25342
rect 27694 25394 27746 25406
rect 32846 25394 32898 25406
rect 29922 25342 29934 25394
rect 29986 25342 29998 25394
rect 27694 25330 27746 25342
rect 32846 25330 32898 25342
rect 33406 25394 33458 25406
rect 36430 25394 36482 25406
rect 35074 25342 35086 25394
rect 35138 25342 35150 25394
rect 33406 25330 33458 25342
rect 36430 25330 36482 25342
rect 38222 25394 38274 25406
rect 41918 25394 41970 25406
rect 38882 25342 38894 25394
rect 38946 25342 38958 25394
rect 38222 25330 38274 25342
rect 41918 25330 41970 25342
rect 43598 25394 43650 25406
rect 43598 25330 43650 25342
rect 45838 25394 45890 25406
rect 45838 25330 45890 25342
rect 3950 25282 4002 25294
rect 3950 25218 4002 25230
rect 4062 25282 4114 25294
rect 15934 25282 15986 25294
rect 4498 25230 4510 25282
rect 4562 25230 4574 25282
rect 4062 25218 4114 25230
rect 15934 25218 15986 25230
rect 16830 25282 16882 25294
rect 16830 25218 16882 25230
rect 19742 25282 19794 25294
rect 19742 25218 19794 25230
rect 20302 25282 20354 25294
rect 20302 25218 20354 25230
rect 21422 25282 21474 25294
rect 21422 25218 21474 25230
rect 22430 25282 22482 25294
rect 22430 25218 22482 25230
rect 23662 25282 23714 25294
rect 26462 25282 26514 25294
rect 24434 25230 24446 25282
rect 24498 25230 24510 25282
rect 23662 25218 23714 25230
rect 26462 25218 26514 25230
rect 28590 25282 28642 25294
rect 28590 25218 28642 25230
rect 35534 25282 35586 25294
rect 43150 25282 43202 25294
rect 37538 25230 37550 25282
rect 37602 25230 37614 25282
rect 40450 25230 40462 25282
rect 40514 25230 40526 25282
rect 35534 25218 35586 25230
rect 43150 25218 43202 25230
rect 43262 25282 43314 25294
rect 43262 25218 43314 25230
rect 43374 25282 43426 25294
rect 45390 25282 45442 25294
rect 43922 25230 43934 25282
rect 43986 25230 43998 25282
rect 43374 25218 43426 25230
rect 45390 25218 45442 25230
rect 45614 25282 45666 25294
rect 45614 25218 45666 25230
rect 1344 25114 49616 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 49616 25114
rect 1344 25028 49616 25062
rect 8430 24946 8482 24958
rect 5842 24894 5854 24946
rect 5906 24894 5918 24946
rect 8430 24882 8482 24894
rect 15598 24946 15650 24958
rect 15598 24882 15650 24894
rect 22654 24946 22706 24958
rect 22654 24882 22706 24894
rect 22766 24946 22818 24958
rect 22766 24882 22818 24894
rect 22990 24946 23042 24958
rect 22990 24882 23042 24894
rect 24446 24946 24498 24958
rect 24446 24882 24498 24894
rect 31054 24946 31106 24958
rect 31054 24882 31106 24894
rect 31614 24946 31666 24958
rect 31614 24882 31666 24894
rect 31838 24946 31890 24958
rect 31838 24882 31890 24894
rect 32622 24946 32674 24958
rect 32622 24882 32674 24894
rect 41358 24946 41410 24958
rect 41358 24882 41410 24894
rect 47182 24946 47234 24958
rect 47182 24882 47234 24894
rect 5406 24834 5458 24846
rect 5406 24770 5458 24782
rect 7646 24834 7698 24846
rect 7646 24770 7698 24782
rect 9998 24834 10050 24846
rect 9998 24770 10050 24782
rect 13806 24834 13858 24846
rect 13806 24770 13858 24782
rect 14590 24834 14642 24846
rect 14590 24770 14642 24782
rect 16158 24834 16210 24846
rect 16158 24770 16210 24782
rect 16270 24834 16322 24846
rect 22430 24834 22482 24846
rect 16818 24782 16830 24834
rect 16882 24782 16894 24834
rect 16270 24770 16322 24782
rect 22430 24770 22482 24782
rect 30830 24834 30882 24846
rect 30830 24770 30882 24782
rect 36654 24834 36706 24846
rect 41582 24834 41634 24846
rect 39218 24782 39230 24834
rect 39282 24782 39294 24834
rect 36654 24770 36706 24782
rect 41582 24770 41634 24782
rect 41694 24834 41746 24846
rect 41694 24770 41746 24782
rect 41918 24834 41970 24846
rect 46286 24834 46338 24846
rect 45826 24782 45838 24834
rect 45890 24782 45902 24834
rect 41918 24770 41970 24782
rect 46286 24770 46338 24782
rect 46734 24834 46786 24846
rect 46734 24770 46786 24782
rect 5182 24722 5234 24734
rect 1810 24670 1822 24722
rect 1874 24670 1886 24722
rect 5182 24658 5234 24670
rect 5294 24722 5346 24734
rect 5294 24658 5346 24670
rect 6302 24722 6354 24734
rect 6302 24658 6354 24670
rect 6638 24722 6690 24734
rect 6638 24658 6690 24670
rect 7982 24722 8034 24734
rect 7982 24658 8034 24670
rect 10334 24722 10386 24734
rect 12574 24722 12626 24734
rect 15262 24722 15314 24734
rect 12114 24670 12126 24722
rect 12178 24670 12190 24722
rect 13122 24670 13134 24722
rect 13186 24670 13198 24722
rect 14018 24670 14030 24722
rect 14082 24670 14094 24722
rect 15026 24670 15038 24722
rect 15090 24670 15102 24722
rect 10334 24658 10386 24670
rect 12574 24658 12626 24670
rect 15262 24658 15314 24670
rect 15486 24722 15538 24734
rect 15486 24658 15538 24670
rect 16382 24722 16434 24734
rect 22878 24722 22930 24734
rect 18162 24670 18174 24722
rect 18226 24670 18238 24722
rect 19394 24670 19406 24722
rect 19458 24670 19470 24722
rect 20738 24670 20750 24722
rect 20802 24670 20814 24722
rect 16382 24658 16434 24670
rect 22878 24658 22930 24670
rect 23886 24722 23938 24734
rect 31390 24722 31442 24734
rect 41470 24722 41522 24734
rect 45502 24722 45554 24734
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 32050 24670 32062 24722
rect 32114 24670 32126 24722
rect 33170 24670 33182 24722
rect 33234 24670 33246 24722
rect 36306 24670 36318 24722
rect 36370 24670 36382 24722
rect 40002 24670 40014 24722
rect 40066 24670 40078 24722
rect 45042 24670 45054 24722
rect 45106 24670 45118 24722
rect 48066 24670 48078 24722
rect 48130 24670 48142 24722
rect 23886 24658 23938 24670
rect 31390 24658 31442 24670
rect 41470 24658 41522 24670
rect 45502 24658 45554 24670
rect 6190 24610 6242 24622
rect 2482 24558 2494 24610
rect 2546 24558 2558 24610
rect 4610 24558 4622 24610
rect 4674 24558 4686 24610
rect 6190 24546 6242 24558
rect 11902 24610 11954 24622
rect 11902 24546 11954 24558
rect 12462 24610 12514 24622
rect 12462 24546 12514 24558
rect 14702 24610 14754 24622
rect 46174 24610 46226 24622
rect 15586 24558 15598 24610
rect 15650 24558 15662 24610
rect 18610 24558 18622 24610
rect 18674 24558 18686 24610
rect 20962 24558 20974 24610
rect 21026 24558 21038 24610
rect 30034 24558 30046 24610
rect 30098 24558 30110 24610
rect 33842 24558 33854 24610
rect 33906 24558 33918 24610
rect 35970 24558 35982 24610
rect 36034 24558 36046 24610
rect 37090 24558 37102 24610
rect 37154 24558 37166 24610
rect 42242 24558 42254 24610
rect 42306 24558 42318 24610
rect 44370 24558 44382 24610
rect 44434 24558 44446 24610
rect 14702 24546 14754 24558
rect 46174 24546 46226 24558
rect 47630 24610 47682 24622
rect 47630 24546 47682 24558
rect 48862 24610 48914 24622
rect 48862 24546 48914 24558
rect 6526 24498 6578 24510
rect 6526 24434 6578 24446
rect 11790 24498 11842 24510
rect 30718 24498 30770 24510
rect 21634 24446 21646 24498
rect 21698 24446 21710 24498
rect 11790 24434 11842 24446
rect 30718 24434 30770 24446
rect 31502 24498 31554 24510
rect 31502 24434 31554 24446
rect 36318 24498 36370 24510
rect 36318 24434 36370 24446
rect 46622 24498 46674 24510
rect 46622 24434 46674 24446
rect 48750 24498 48802 24510
rect 48750 24434 48802 24446
rect 1344 24330 49616 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 49616 24330
rect 1344 24244 49616 24278
rect 12574 24162 12626 24174
rect 14814 24162 14866 24174
rect 12898 24110 12910 24162
rect 12962 24110 12974 24162
rect 13458 24110 13470 24162
rect 13522 24110 13534 24162
rect 12574 24098 12626 24110
rect 14814 24098 14866 24110
rect 15710 24162 15762 24174
rect 15710 24098 15762 24110
rect 34862 24162 34914 24174
rect 34862 24098 34914 24110
rect 38446 24162 38498 24174
rect 38446 24098 38498 24110
rect 6078 24050 6130 24062
rect 4610 23998 4622 24050
rect 4674 23998 4686 24050
rect 6078 23986 6130 23998
rect 6638 24050 6690 24062
rect 8206 24050 8258 24062
rect 12350 24050 12402 24062
rect 7858 23998 7870 24050
rect 7922 23998 7934 24050
rect 9874 23998 9886 24050
rect 9938 23998 9950 24050
rect 12002 23998 12014 24050
rect 12066 23998 12078 24050
rect 6638 23986 6690 23998
rect 8206 23986 8258 23998
rect 12350 23986 12402 23998
rect 15486 24050 15538 24062
rect 15486 23986 15538 23998
rect 16046 24050 16098 24062
rect 29262 24050 29314 24062
rect 36430 24050 36482 24062
rect 37998 24050 38050 24062
rect 48414 24050 48466 24062
rect 17042 23998 17054 24050
rect 17106 23998 17118 24050
rect 17826 23998 17838 24050
rect 17890 23998 17902 24050
rect 19954 23998 19966 24050
rect 20018 23998 20030 24050
rect 21522 23998 21534 24050
rect 21586 23998 21598 24050
rect 32946 23998 32958 24050
rect 33010 23998 33022 24050
rect 36082 23998 36094 24050
rect 36146 23998 36158 24050
rect 37538 23998 37550 24050
rect 37602 23998 37614 24050
rect 38994 23998 39006 24050
rect 39058 23998 39070 24050
rect 39890 23998 39902 24050
rect 39954 23998 39966 24050
rect 40674 23998 40686 24050
rect 40738 23998 40750 24050
rect 45602 23998 45614 24050
rect 45666 23998 45678 24050
rect 47730 23998 47742 24050
rect 47794 23998 47806 24050
rect 16046 23986 16098 23998
rect 29262 23986 29314 23998
rect 36430 23986 36482 23998
rect 37998 23986 38050 23998
rect 48414 23986 48466 23998
rect 49198 24050 49250 24062
rect 49198 23986 49250 23998
rect 5630 23938 5682 23950
rect 13918 23938 13970 23950
rect 27694 23938 27746 23950
rect 28366 23938 28418 23950
rect 1810 23886 1822 23938
rect 1874 23886 1886 23938
rect 7746 23886 7758 23938
rect 7810 23886 7822 23938
rect 9090 23886 9102 23938
rect 9154 23886 9166 23938
rect 14242 23886 14254 23938
rect 14306 23886 14318 23938
rect 16370 23886 16382 23938
rect 16434 23886 16446 23938
rect 17490 23886 17502 23938
rect 17554 23886 17566 23938
rect 20738 23886 20750 23938
rect 20802 23886 20814 23938
rect 25442 23886 25454 23938
rect 25506 23886 25518 23938
rect 27458 23886 27470 23938
rect 27522 23886 27534 23938
rect 28018 23886 28030 23938
rect 28082 23886 28094 23938
rect 5630 23874 5682 23886
rect 13918 23874 13970 23886
rect 27694 23874 27746 23886
rect 28366 23874 28418 23886
rect 29822 23938 29874 23950
rect 34414 23938 34466 23950
rect 30146 23886 30158 23938
rect 30210 23886 30222 23938
rect 29822 23874 29874 23886
rect 34414 23874 34466 23886
rect 34974 23938 35026 23950
rect 34974 23874 35026 23886
rect 35198 23938 35250 23950
rect 38558 23938 38610 23950
rect 48190 23938 48242 23950
rect 35410 23886 35422 23938
rect 35474 23886 35486 23938
rect 37314 23886 37326 23938
rect 37378 23886 37390 23938
rect 43474 23886 43486 23938
rect 43538 23886 43550 23938
rect 44146 23886 44158 23938
rect 44210 23886 44222 23938
rect 44818 23886 44830 23938
rect 44882 23886 44894 23938
rect 35198 23874 35250 23886
rect 38558 23874 38610 23886
rect 48190 23874 48242 23886
rect 48302 23938 48354 23950
rect 48302 23874 48354 23886
rect 5854 23826 5906 23838
rect 2482 23774 2494 23826
rect 2546 23774 2558 23826
rect 5854 23762 5906 23774
rect 6190 23826 6242 23838
rect 6190 23762 6242 23774
rect 14030 23826 14082 23838
rect 14030 23762 14082 23774
rect 14590 23826 14642 23838
rect 33854 23826 33906 23838
rect 48526 23826 48578 23838
rect 16706 23774 16718 23826
rect 16770 23774 16782 23826
rect 30818 23774 30830 23826
rect 30882 23774 30894 23826
rect 42802 23774 42814 23826
rect 42866 23774 42878 23826
rect 43922 23774 43934 23826
rect 43986 23774 43998 23826
rect 14590 23762 14642 23774
rect 33854 23762 33906 23774
rect 48526 23762 48578 23774
rect 48750 23826 48802 23838
rect 48750 23762 48802 23774
rect 8766 23714 8818 23726
rect 26910 23714 26962 23726
rect 15138 23662 15150 23714
rect 15202 23662 15214 23714
rect 8766 23650 8818 23662
rect 26910 23650 26962 23662
rect 27022 23714 27074 23726
rect 27022 23650 27074 23662
rect 27134 23714 27186 23726
rect 27134 23650 27186 23662
rect 27806 23714 27858 23726
rect 27806 23650 27858 23662
rect 29150 23714 29202 23726
rect 29150 23650 29202 23662
rect 29374 23714 29426 23726
rect 29374 23650 29426 23662
rect 33518 23714 33570 23726
rect 33518 23650 33570 23662
rect 33742 23714 33794 23726
rect 33742 23650 33794 23662
rect 34526 23714 34578 23726
rect 34526 23650 34578 23662
rect 38446 23714 38498 23726
rect 38446 23650 38498 23662
rect 39454 23714 39506 23726
rect 39454 23650 39506 23662
rect 40350 23714 40402 23726
rect 40350 23650 40402 23662
rect 1344 23546 49616 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 49616 23546
rect 1344 23460 49616 23494
rect 11790 23378 11842 23390
rect 16494 23378 16546 23390
rect 10434 23326 10446 23378
rect 10498 23326 10510 23378
rect 15810 23326 15822 23378
rect 15874 23326 15886 23378
rect 11790 23314 11842 23326
rect 16494 23314 16546 23326
rect 25342 23378 25394 23390
rect 25342 23314 25394 23326
rect 29150 23378 29202 23390
rect 29150 23314 29202 23326
rect 29822 23378 29874 23390
rect 29822 23314 29874 23326
rect 30270 23378 30322 23390
rect 30270 23314 30322 23326
rect 30382 23378 30434 23390
rect 31502 23378 31554 23390
rect 31154 23326 31166 23378
rect 31218 23326 31230 23378
rect 30382 23314 30434 23326
rect 31502 23314 31554 23326
rect 32622 23378 32674 23390
rect 35086 23378 35138 23390
rect 36990 23378 37042 23390
rect 33282 23326 33294 23378
rect 33346 23326 33358 23378
rect 36530 23326 36542 23378
rect 36594 23326 36606 23378
rect 32622 23314 32674 23326
rect 35086 23314 35138 23326
rect 36990 23314 37042 23326
rect 37214 23378 37266 23390
rect 37214 23314 37266 23326
rect 38894 23378 38946 23390
rect 38894 23314 38946 23326
rect 41022 23378 41074 23390
rect 41022 23314 41074 23326
rect 41134 23378 41186 23390
rect 41134 23314 41186 23326
rect 41806 23378 41858 23390
rect 41806 23314 41858 23326
rect 42030 23378 42082 23390
rect 42030 23314 42082 23326
rect 3390 23266 3442 23278
rect 3390 23202 3442 23214
rect 4286 23266 4338 23278
rect 4286 23202 4338 23214
rect 5742 23266 5794 23278
rect 11678 23266 11730 23278
rect 6850 23214 6862 23266
rect 6914 23214 6926 23266
rect 5742 23202 5794 23214
rect 11678 23202 11730 23214
rect 12014 23266 12066 23278
rect 12014 23202 12066 23214
rect 12238 23266 12290 23278
rect 16606 23266 16658 23278
rect 13346 23214 13358 23266
rect 13410 23214 13422 23266
rect 12238 23202 12290 23214
rect 16606 23202 16658 23214
rect 19182 23266 19234 23278
rect 19182 23202 19234 23214
rect 19630 23266 19682 23278
rect 28926 23266 28978 23278
rect 23426 23214 23438 23266
rect 23490 23214 23502 23266
rect 26450 23214 26462 23266
rect 26514 23214 26526 23266
rect 19630 23202 19682 23214
rect 28926 23202 28978 23214
rect 30494 23266 30546 23278
rect 30494 23202 30546 23214
rect 31950 23266 32002 23278
rect 36878 23266 36930 23278
rect 38222 23266 38274 23278
rect 35410 23214 35422 23266
rect 35474 23214 35486 23266
rect 37538 23214 37550 23266
rect 37602 23214 37614 23266
rect 31950 23202 32002 23214
rect 36878 23202 36930 23214
rect 38222 23202 38274 23214
rect 40910 23266 40962 23278
rect 44930 23214 44942 23266
rect 44994 23214 45006 23266
rect 40910 23202 40962 23214
rect 3614 23154 3666 23166
rect 3614 23090 3666 23102
rect 4062 23154 4114 23166
rect 4062 23090 4114 23102
rect 4398 23154 4450 23166
rect 4398 23090 4450 23102
rect 4622 23154 4674 23166
rect 5070 23154 5122 23166
rect 4834 23102 4846 23154
rect 4898 23102 4910 23154
rect 4622 23090 4674 23102
rect 5070 23090 5122 23102
rect 5294 23154 5346 23166
rect 5294 23090 5346 23102
rect 5406 23154 5458 23166
rect 10782 23154 10834 23166
rect 6178 23102 6190 23154
rect 6242 23102 6254 23154
rect 5406 23090 5458 23102
rect 10782 23090 10834 23102
rect 11006 23154 11058 23166
rect 18958 23154 19010 23166
rect 19966 23154 20018 23166
rect 12674 23102 12686 23154
rect 12738 23102 12750 23154
rect 16034 23102 16046 23154
rect 16098 23102 16110 23154
rect 19394 23102 19406 23154
rect 19458 23102 19470 23154
rect 11006 23090 11058 23102
rect 18958 23090 19010 23102
rect 19966 23090 20018 23102
rect 20190 23154 20242 23166
rect 20190 23090 20242 23102
rect 20638 23154 20690 23166
rect 29486 23154 29538 23166
rect 24210 23102 24222 23154
rect 24274 23102 24286 23154
rect 25666 23102 25678 23154
rect 25730 23102 25742 23154
rect 20638 23090 20690 23102
rect 29486 23090 29538 23102
rect 30942 23154 30994 23166
rect 37886 23154 37938 23166
rect 34178 23102 34190 23154
rect 34242 23102 34254 23154
rect 30942 23090 30994 23102
rect 37886 23090 37938 23102
rect 38334 23154 38386 23166
rect 43362 23102 43374 23154
rect 43426 23102 43438 23154
rect 38334 23090 38386 23102
rect 3502 23042 3554 23054
rect 18062 23042 18114 23054
rect 8978 22990 8990 23042
rect 9042 22990 9054 23042
rect 15474 22990 15486 23042
rect 15538 22990 15550 23042
rect 3502 22978 3554 22990
rect 18062 22978 18114 22990
rect 18510 23042 18562 23054
rect 18510 22978 18562 22990
rect 20078 23042 20130 23054
rect 20078 22978 20130 22990
rect 20974 23042 21026 23054
rect 24670 23042 24722 23054
rect 33630 23042 33682 23054
rect 21298 22990 21310 23042
rect 21362 22990 21374 23042
rect 28578 22990 28590 23042
rect 28642 22990 28654 23042
rect 20974 22978 21026 22990
rect 24670 22978 24722 22990
rect 33630 22978 33682 22990
rect 33854 23042 33906 23054
rect 33854 22978 33906 22990
rect 34750 23042 34802 23054
rect 34750 22978 34802 22990
rect 35982 23042 36034 23054
rect 35982 22978 36034 22990
rect 39230 23042 39282 23054
rect 39230 22978 39282 22990
rect 39678 23042 39730 23054
rect 39678 22978 39730 22990
rect 40126 23042 40178 23054
rect 40126 22978 40178 22990
rect 42590 23042 42642 23054
rect 42590 22978 42642 22990
rect 48862 23042 48914 23054
rect 48862 22978 48914 22990
rect 19070 22930 19122 22942
rect 19070 22866 19122 22878
rect 29262 22930 29314 22942
rect 34526 22930 34578 22942
rect 31938 22878 31950 22930
rect 32002 22927 32014 22930
rect 32610 22927 32622 22930
rect 32002 22881 32622 22927
rect 32002 22878 32014 22881
rect 32610 22878 32622 22881
rect 32674 22878 32686 22930
rect 29262 22866 29314 22878
rect 34526 22866 34578 22878
rect 36206 22930 36258 22942
rect 36206 22866 36258 22878
rect 48750 22930 48802 22942
rect 48750 22866 48802 22878
rect 1344 22762 49616 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 49616 22762
rect 1344 22676 49616 22710
rect 33282 22591 33294 22594
rect 32401 22545 33294 22591
rect 17054 22482 17106 22494
rect 20638 22482 20690 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 9090 22430 9102 22482
rect 9154 22430 9166 22482
rect 17266 22430 17278 22482
rect 17330 22430 17342 22482
rect 17054 22418 17106 22430
rect 20638 22418 20690 22430
rect 21422 22482 21474 22494
rect 29262 22482 29314 22494
rect 21746 22430 21758 22482
rect 21810 22430 21822 22482
rect 28130 22430 28142 22482
rect 28194 22430 28206 22482
rect 21422 22418 21474 22430
rect 29262 22418 29314 22430
rect 30382 22482 30434 22494
rect 30382 22418 30434 22430
rect 32062 22482 32114 22494
rect 32401 22482 32447 22545
rect 33282 22542 33294 22545
rect 33346 22542 33358 22594
rect 33618 22542 33630 22594
rect 33682 22542 33694 22594
rect 37762 22542 37774 22594
rect 37826 22542 37838 22594
rect 38882 22542 38894 22594
rect 38946 22542 38958 22594
rect 34638 22482 34690 22494
rect 43374 22482 43426 22494
rect 44942 22482 44994 22494
rect 32386 22430 32398 22482
rect 32450 22430 32462 22482
rect 41682 22430 41694 22482
rect 41746 22430 41758 22482
rect 42578 22430 42590 22482
rect 42642 22430 42654 22482
rect 44146 22430 44158 22482
rect 44210 22430 44222 22482
rect 47058 22430 47070 22482
rect 47122 22430 47134 22482
rect 49186 22430 49198 22482
rect 49250 22430 49262 22482
rect 32062 22418 32114 22430
rect 34638 22418 34690 22430
rect 43374 22418 43426 22430
rect 44942 22418 44994 22430
rect 11342 22370 11394 22382
rect 29934 22370 29986 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 6626 22318 6638 22370
rect 6690 22318 6702 22370
rect 20178 22318 20190 22370
rect 20242 22318 20254 22370
rect 24658 22318 24670 22370
rect 24722 22318 24734 22370
rect 25330 22318 25342 22370
rect 25394 22318 25406 22370
rect 11342 22306 11394 22318
rect 29934 22306 29986 22318
rect 31838 22370 31890 22382
rect 31838 22306 31890 22318
rect 33966 22370 34018 22382
rect 33966 22306 34018 22318
rect 34190 22370 34242 22382
rect 34190 22306 34242 22318
rect 35198 22370 35250 22382
rect 35198 22306 35250 22318
rect 38334 22370 38386 22382
rect 38334 22306 38386 22318
rect 38558 22370 38610 22382
rect 38558 22306 38610 22318
rect 39566 22370 39618 22382
rect 42142 22370 42194 22382
rect 45166 22370 45218 22382
rect 40674 22318 40686 22370
rect 40738 22318 40750 22370
rect 41346 22318 41358 22370
rect 41410 22318 41422 22370
rect 43810 22318 43822 22370
rect 43874 22318 43886 22370
rect 39566 22306 39618 22318
rect 42142 22306 42194 22318
rect 45166 22306 45218 22318
rect 45950 22370 46002 22382
rect 46274 22318 46286 22370
rect 46338 22318 46350 22370
rect 45950 22306 46002 22318
rect 29598 22258 29650 22270
rect 2482 22206 2494 22258
rect 2546 22206 2558 22258
rect 19394 22206 19406 22258
rect 19458 22206 19470 22258
rect 23874 22206 23886 22258
rect 23938 22206 23950 22258
rect 26002 22206 26014 22258
rect 26066 22206 26078 22258
rect 29598 22194 29650 22206
rect 31390 22258 31442 22270
rect 31390 22194 31442 22206
rect 31614 22258 31666 22270
rect 31614 22194 31666 22206
rect 32174 22258 32226 22270
rect 32174 22194 32226 22206
rect 32622 22258 32674 22270
rect 32622 22194 32674 22206
rect 33070 22258 33122 22270
rect 37102 22258 37154 22270
rect 35522 22206 35534 22258
rect 35586 22206 35598 22258
rect 33070 22194 33122 22206
rect 37102 22194 37154 22206
rect 37214 22258 37266 22270
rect 37214 22194 37266 22206
rect 37326 22258 37378 22270
rect 37326 22194 37378 22206
rect 39230 22258 39282 22270
rect 39230 22194 39282 22206
rect 40014 22258 40066 22270
rect 40014 22194 40066 22206
rect 43262 22258 43314 22270
rect 43262 22194 43314 22206
rect 28590 22146 28642 22158
rect 28590 22082 28642 22094
rect 30942 22146 30994 22158
rect 30942 22082 30994 22094
rect 36094 22146 36146 22158
rect 39902 22146 39954 22158
rect 36418 22094 36430 22146
rect 36482 22094 36494 22146
rect 36094 22082 36146 22094
rect 39902 22082 39954 22094
rect 40910 22146 40962 22158
rect 45490 22094 45502 22146
rect 45554 22094 45566 22146
rect 40910 22082 40962 22094
rect 1344 21978 49616 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 49616 21978
rect 1344 21892 49616 21926
rect 2718 21810 2770 21822
rect 2718 21746 2770 21758
rect 8766 21810 8818 21822
rect 8766 21746 8818 21758
rect 9662 21810 9714 21822
rect 9662 21746 9714 21758
rect 14030 21810 14082 21822
rect 14030 21746 14082 21758
rect 20862 21810 20914 21822
rect 20862 21746 20914 21758
rect 26350 21810 26402 21822
rect 26350 21746 26402 21758
rect 26462 21810 26514 21822
rect 26462 21746 26514 21758
rect 27470 21810 27522 21822
rect 33070 21810 33122 21822
rect 27906 21758 27918 21810
rect 27970 21758 27982 21810
rect 30594 21758 30606 21810
rect 30658 21758 30670 21810
rect 27470 21746 27522 21758
rect 2830 21698 2882 21710
rect 2830 21634 2882 21646
rect 10222 21698 10274 21710
rect 10222 21634 10274 21646
rect 10558 21698 10610 21710
rect 21198 21698 21250 21710
rect 10882 21646 10894 21698
rect 10946 21646 10958 21698
rect 19506 21646 19518 21698
rect 19570 21646 19582 21698
rect 10558 21634 10610 21646
rect 21198 21634 21250 21646
rect 27694 21698 27746 21710
rect 27694 21634 27746 21646
rect 8542 21586 8594 21598
rect 5506 21534 5518 21586
rect 5570 21534 5582 21586
rect 8542 21522 8594 21534
rect 8878 21586 8930 21598
rect 8878 21522 8930 21534
rect 9774 21586 9826 21598
rect 9774 21522 9826 21534
rect 11454 21586 11506 21598
rect 13358 21586 13410 21598
rect 16046 21586 16098 21598
rect 21086 21586 21138 21598
rect 12450 21534 12462 21586
rect 12514 21534 12526 21586
rect 14242 21534 14254 21586
rect 14306 21534 14318 21586
rect 20290 21534 20302 21586
rect 20354 21534 20366 21586
rect 11454 21522 11506 21534
rect 13358 21522 13410 21534
rect 16046 21522 16098 21534
rect 21086 21522 21138 21534
rect 21310 21586 21362 21598
rect 25342 21586 25394 21598
rect 21746 21534 21758 21586
rect 21810 21534 21822 21586
rect 21310 21522 21362 21534
rect 25342 21522 25394 21534
rect 25790 21586 25842 21598
rect 25790 21522 25842 21534
rect 26014 21586 26066 21598
rect 26014 21522 26066 21534
rect 26574 21586 26626 21598
rect 26574 21522 26626 21534
rect 27022 21586 27074 21598
rect 27022 21522 27074 21534
rect 27134 21586 27186 21598
rect 27134 21522 27186 21534
rect 11230 21474 11282 21486
rect 6178 21422 6190 21474
rect 6242 21422 6254 21474
rect 8306 21422 8318 21474
rect 8370 21422 8382 21474
rect 11230 21410 11282 21422
rect 11790 21474 11842 21486
rect 13134 21474 13186 21486
rect 12114 21422 12126 21474
rect 12178 21422 12190 21474
rect 11790 21410 11842 21422
rect 13134 21410 13186 21422
rect 16494 21474 16546 21486
rect 16494 21410 16546 21422
rect 16830 21474 16882 21486
rect 25902 21474 25954 21486
rect 17378 21422 17390 21474
rect 17442 21422 17454 21474
rect 22418 21422 22430 21474
rect 22482 21422 22494 21474
rect 24546 21422 24558 21474
rect 24610 21422 24622 21474
rect 16830 21410 16882 21422
rect 25902 21410 25954 21422
rect 9662 21362 9714 21374
rect 27358 21362 27410 21374
rect 27921 21362 27967 21758
rect 33070 21746 33122 21758
rect 33294 21810 33346 21822
rect 33294 21746 33346 21758
rect 34078 21810 34130 21822
rect 34078 21746 34130 21758
rect 35982 21810 36034 21822
rect 35982 21746 36034 21758
rect 36654 21810 36706 21822
rect 36654 21746 36706 21758
rect 46846 21810 46898 21822
rect 46846 21746 46898 21758
rect 47294 21810 47346 21822
rect 47294 21746 47346 21758
rect 47742 21810 47794 21822
rect 47742 21746 47794 21758
rect 29598 21698 29650 21710
rect 29598 21634 29650 21646
rect 29710 21698 29762 21710
rect 36206 21698 36258 21710
rect 46958 21698 47010 21710
rect 31938 21646 31950 21698
rect 32002 21646 32014 21698
rect 46050 21646 46062 21698
rect 46114 21646 46126 21698
rect 29710 21634 29762 21646
rect 36206 21634 36258 21646
rect 46958 21634 47010 21646
rect 28254 21586 28306 21598
rect 28254 21522 28306 21534
rect 28478 21586 28530 21598
rect 28478 21522 28530 21534
rect 28702 21586 28754 21598
rect 28702 21522 28754 21534
rect 29822 21586 29874 21598
rect 29822 21522 29874 21534
rect 30270 21586 30322 21598
rect 30270 21522 30322 21534
rect 31278 21586 31330 21598
rect 31278 21522 31330 21534
rect 31390 21586 31442 21598
rect 31390 21522 31442 21534
rect 31502 21586 31554 21598
rect 31502 21522 31554 21534
rect 33742 21586 33794 21598
rect 33742 21522 33794 21534
rect 34190 21586 34242 21598
rect 34190 21522 34242 21534
rect 35086 21586 35138 21598
rect 35086 21522 35138 21534
rect 35534 21586 35586 21598
rect 35534 21522 35586 21534
rect 36542 21586 36594 21598
rect 36542 21522 36594 21534
rect 36766 21586 36818 21598
rect 41358 21586 41410 21598
rect 46398 21586 46450 21598
rect 37090 21534 37102 21586
rect 37154 21534 37166 21586
rect 37538 21534 37550 21586
rect 37602 21534 37614 21586
rect 42466 21534 42478 21586
rect 42530 21534 42542 21586
rect 45826 21534 45838 21586
rect 45890 21534 45902 21586
rect 36766 21522 36818 21534
rect 41358 21522 41410 21534
rect 46398 21522 46450 21534
rect 46734 21586 46786 21598
rect 46734 21522 46786 21534
rect 47518 21586 47570 21598
rect 48738 21534 48750 21586
rect 48802 21534 48814 21586
rect 47518 21522 47570 21534
rect 28366 21474 28418 21486
rect 28366 21410 28418 21422
rect 32398 21474 32450 21486
rect 32398 21410 32450 21422
rect 33182 21474 33234 21486
rect 33182 21410 33234 21422
rect 34638 21474 34690 21486
rect 41022 21474 41074 21486
rect 47406 21474 47458 21486
rect 38210 21422 38222 21474
rect 38274 21422 38286 21474
rect 40338 21422 40350 21474
rect 40402 21422 40414 21474
rect 41794 21422 41806 21474
rect 41858 21422 41870 21474
rect 43250 21422 43262 21474
rect 43314 21422 43326 21474
rect 45378 21422 45390 21474
rect 45442 21422 45454 21474
rect 34638 21410 34690 21422
rect 41022 21410 41074 21422
rect 47406 21410 47458 21422
rect 34078 21362 34130 21374
rect 13682 21310 13694 21362
rect 13746 21310 13758 21362
rect 27906 21310 27918 21362
rect 27970 21310 27982 21362
rect 29138 21310 29150 21362
rect 29202 21310 29214 21362
rect 9662 21298 9714 21310
rect 27358 21298 27410 21310
rect 34078 21298 34130 21310
rect 35422 21362 35474 21374
rect 35422 21298 35474 21310
rect 35870 21362 35922 21374
rect 35870 21298 35922 21310
rect 40910 21362 40962 21374
rect 40910 21298 40962 21310
rect 48750 21362 48802 21374
rect 48750 21298 48802 21310
rect 49086 21362 49138 21374
rect 49086 21298 49138 21310
rect 1344 21194 49616 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 49616 21194
rect 1344 21108 49616 21142
rect 17950 21026 18002 21038
rect 35086 21026 35138 21038
rect 34402 20974 34414 21026
rect 34466 21023 34478 21026
rect 34850 21023 34862 21026
rect 34466 20977 34862 21023
rect 34466 20974 34478 20977
rect 34850 20974 34862 20977
rect 34914 20974 34926 21026
rect 17950 20962 18002 20974
rect 35086 20962 35138 20974
rect 35422 21026 35474 21038
rect 38322 20974 38334 21026
rect 38386 20974 38398 21026
rect 35422 20962 35474 20974
rect 18174 20914 18226 20926
rect 22318 20914 22370 20926
rect 4610 20862 4622 20914
rect 4674 20862 4686 20914
rect 9650 20862 9662 20914
rect 9714 20862 9726 20914
rect 10770 20862 10782 20914
rect 10834 20862 10846 20914
rect 12898 20862 12910 20914
rect 12962 20862 12974 20914
rect 17042 20862 17054 20914
rect 17106 20862 17118 20914
rect 19282 20862 19294 20914
rect 19346 20862 19358 20914
rect 21410 20862 21422 20914
rect 21474 20862 21486 20914
rect 18174 20850 18226 20862
rect 22318 20850 22370 20862
rect 22766 20914 22818 20926
rect 39454 20914 39506 20926
rect 24546 20862 24558 20914
rect 24610 20862 24622 20914
rect 26674 20862 26686 20914
rect 26738 20862 26750 20914
rect 30706 20862 30718 20914
rect 30770 20862 30782 20914
rect 32834 20862 32846 20914
rect 32898 20862 32910 20914
rect 22766 20850 22818 20862
rect 39454 20850 39506 20862
rect 40126 20914 40178 20926
rect 47058 20862 47070 20914
rect 47122 20862 47134 20914
rect 49186 20862 49198 20914
rect 49250 20862 49262 20914
rect 40126 20850 40178 20862
rect 6526 20802 6578 20814
rect 17390 20802 17442 20814
rect 1810 20750 1822 20802
rect 1874 20750 1886 20802
rect 6738 20750 6750 20802
rect 6802 20750 6814 20802
rect 10098 20750 10110 20802
rect 10162 20750 10174 20802
rect 14130 20750 14142 20802
rect 14194 20750 14206 20802
rect 6526 20738 6578 20750
rect 17390 20738 17442 20750
rect 18398 20802 18450 20814
rect 18398 20738 18450 20750
rect 18734 20802 18786 20814
rect 18734 20738 18786 20750
rect 18958 20802 19010 20814
rect 18958 20738 19010 20750
rect 19742 20802 19794 20814
rect 22654 20802 22706 20814
rect 21522 20750 21534 20802
rect 21586 20750 21598 20802
rect 21746 20750 21758 20802
rect 21810 20750 21822 20802
rect 19742 20738 19794 20750
rect 22654 20738 22706 20750
rect 22878 20802 22930 20814
rect 27246 20802 27298 20814
rect 29486 20802 29538 20814
rect 34190 20802 34242 20814
rect 23874 20750 23886 20802
rect 23938 20750 23950 20802
rect 28018 20750 28030 20802
rect 28082 20750 28094 20802
rect 30034 20750 30046 20802
rect 30098 20750 30110 20802
rect 33618 20750 33630 20802
rect 33682 20750 33694 20802
rect 22878 20738 22930 20750
rect 27246 20738 27298 20750
rect 29486 20738 29538 20750
rect 34190 20738 34242 20750
rect 35982 20802 36034 20814
rect 35982 20738 36034 20750
rect 36318 20802 36370 20814
rect 37326 20802 37378 20814
rect 39230 20802 39282 20814
rect 37090 20750 37102 20802
rect 37154 20750 37166 20802
rect 38322 20750 38334 20802
rect 38386 20750 38398 20802
rect 38658 20750 38670 20802
rect 38722 20750 38734 20802
rect 36318 20738 36370 20750
rect 37326 20738 37378 20750
rect 39230 20738 39282 20750
rect 39678 20802 39730 20814
rect 39678 20738 39730 20750
rect 39790 20802 39842 20814
rect 39790 20738 39842 20750
rect 40350 20802 40402 20814
rect 43150 20802 43202 20814
rect 42018 20750 42030 20802
rect 42082 20750 42094 20802
rect 40350 20738 40402 20750
rect 43150 20738 43202 20750
rect 45726 20802 45778 20814
rect 46274 20750 46286 20802
rect 46338 20750 46350 20802
rect 45726 20738 45778 20750
rect 5854 20690 5906 20702
rect 2482 20638 2494 20690
rect 2546 20638 2558 20690
rect 5854 20626 5906 20638
rect 6078 20690 6130 20702
rect 20750 20690 20802 20702
rect 7522 20638 7534 20690
rect 7586 20638 7598 20690
rect 14914 20638 14926 20690
rect 14978 20638 14990 20690
rect 17714 20638 17726 20690
rect 17778 20638 17790 20690
rect 20402 20638 20414 20690
rect 20466 20638 20478 20690
rect 6078 20626 6130 20638
rect 20750 20626 20802 20638
rect 27022 20690 27074 20702
rect 27022 20626 27074 20638
rect 27582 20690 27634 20702
rect 27582 20626 27634 20638
rect 35198 20690 35250 20702
rect 35198 20626 35250 20638
rect 35758 20690 35810 20702
rect 35758 20626 35810 20638
rect 37438 20690 37490 20702
rect 42366 20690 42418 20702
rect 40450 20638 40462 20690
rect 40514 20638 40526 20690
rect 41010 20638 41022 20690
rect 41074 20638 41086 20690
rect 37438 20626 37490 20638
rect 42366 20626 42418 20638
rect 42702 20690 42754 20702
rect 42702 20626 42754 20638
rect 43710 20690 43762 20702
rect 43710 20626 43762 20638
rect 44046 20690 44098 20702
rect 44046 20626 44098 20638
rect 44942 20690 44994 20702
rect 44942 20626 44994 20638
rect 45950 20690 46002 20702
rect 45950 20626 46002 20638
rect 6190 20578 6242 20590
rect 19630 20578 19682 20590
rect 17826 20526 17838 20578
rect 17890 20526 17902 20578
rect 6190 20514 6242 20526
rect 19630 20514 19682 20526
rect 21310 20578 21362 20590
rect 21310 20514 21362 20526
rect 23102 20578 23154 20590
rect 23102 20514 23154 20526
rect 27358 20578 27410 20590
rect 29598 20578 29650 20590
rect 28242 20526 28254 20578
rect 28306 20526 28318 20578
rect 27358 20514 27410 20526
rect 29598 20514 29650 20526
rect 29710 20578 29762 20590
rect 29710 20514 29762 20526
rect 33854 20578 33906 20590
rect 33854 20514 33906 20526
rect 34078 20578 34130 20590
rect 34078 20514 34130 20526
rect 34750 20578 34802 20590
rect 34750 20514 34802 20526
rect 35870 20578 35922 20590
rect 42254 20578 42306 20590
rect 37874 20526 37886 20578
rect 37938 20526 37950 20578
rect 35870 20514 35922 20526
rect 42254 20514 42306 20526
rect 42478 20578 42530 20590
rect 42478 20514 42530 20526
rect 43262 20578 43314 20590
rect 43262 20514 43314 20526
rect 43374 20578 43426 20590
rect 43374 20514 43426 20526
rect 43486 20578 43538 20590
rect 43486 20514 43538 20526
rect 44158 20578 44210 20590
rect 44158 20514 44210 20526
rect 45054 20578 45106 20590
rect 45378 20526 45390 20578
rect 45442 20526 45454 20578
rect 45054 20514 45106 20526
rect 1344 20410 49616 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 49616 20410
rect 1344 20324 49616 20358
rect 3054 20242 3106 20254
rect 9662 20242 9714 20254
rect 8306 20190 8318 20242
rect 8370 20190 8382 20242
rect 3054 20178 3106 20190
rect 9662 20178 9714 20190
rect 23998 20242 24050 20254
rect 23998 20178 24050 20190
rect 41246 20242 41298 20254
rect 41246 20178 41298 20190
rect 2494 20130 2546 20142
rect 2494 20066 2546 20078
rect 2718 20130 2770 20142
rect 13470 20130 13522 20142
rect 7410 20078 7422 20130
rect 7474 20078 7486 20130
rect 8866 20078 8878 20130
rect 8930 20078 8942 20130
rect 2718 20066 2770 20078
rect 13470 20066 13522 20078
rect 15374 20130 15426 20142
rect 15374 20066 15426 20078
rect 16270 20130 16322 20142
rect 16270 20066 16322 20078
rect 16382 20130 16434 20142
rect 16382 20066 16434 20078
rect 22654 20130 22706 20142
rect 22654 20066 22706 20078
rect 23774 20130 23826 20142
rect 24670 20130 24722 20142
rect 24322 20078 24334 20130
rect 24386 20078 24398 20130
rect 23774 20066 23826 20078
rect 24670 20066 24722 20078
rect 41582 20130 41634 20142
rect 44370 20078 44382 20130
rect 44434 20078 44446 20130
rect 46722 20078 46734 20130
rect 46786 20078 46798 20130
rect 47394 20078 47406 20130
rect 47458 20078 47470 20130
rect 49074 20078 49086 20130
rect 49138 20078 49150 20130
rect 41582 20066 41634 20078
rect 2382 20018 2434 20030
rect 2382 19954 2434 19966
rect 2830 20018 2882 20030
rect 2830 19954 2882 19966
rect 3166 20018 3218 20030
rect 3166 19954 3218 19966
rect 3502 20018 3554 20030
rect 9438 20018 9490 20030
rect 3938 19966 3950 20018
rect 4002 19966 4014 20018
rect 7298 19966 7310 20018
rect 7362 19966 7374 20018
rect 8418 19966 8430 20018
rect 8482 19966 8494 20018
rect 3502 19954 3554 19966
rect 9438 19954 9490 19966
rect 9774 20018 9826 20030
rect 9774 19954 9826 19966
rect 14366 20018 14418 20030
rect 14366 19954 14418 19966
rect 14478 20018 14530 20030
rect 15934 20018 15986 20030
rect 14690 19966 14702 20018
rect 14754 19966 14766 20018
rect 15586 19966 15598 20018
rect 15650 19966 15662 20018
rect 14478 19954 14530 19966
rect 15934 19954 15986 19966
rect 16046 20018 16098 20030
rect 22878 20018 22930 20030
rect 21970 19966 21982 20018
rect 22034 19966 22046 20018
rect 16046 19954 16098 19966
rect 22878 19954 22930 19966
rect 23326 20018 23378 20030
rect 23326 19954 23378 19966
rect 23438 20018 23490 20030
rect 34190 20018 34242 20030
rect 25554 19966 25566 20018
rect 25618 19966 25630 20018
rect 23438 19954 23490 19966
rect 34190 19954 34242 19966
rect 34414 20018 34466 20030
rect 41134 20018 41186 20030
rect 35074 19966 35086 20018
rect 35138 19966 35150 20018
rect 40898 19966 40910 20018
rect 40962 19966 40974 20018
rect 34414 19954 34466 19966
rect 41134 19954 41186 19966
rect 41358 20018 41410 20030
rect 45502 20018 45554 20030
rect 45154 19966 45166 20018
rect 45218 19966 45230 20018
rect 41358 19954 41410 19966
rect 45502 19954 45554 19966
rect 45726 20018 45778 20030
rect 45726 19954 45778 19966
rect 46174 20018 46226 20030
rect 48750 20018 48802 20030
rect 46610 19966 46622 20018
rect 46674 19966 46686 20018
rect 47842 19966 47854 20018
rect 47906 19966 47918 20018
rect 48178 19966 48190 20018
rect 48242 19966 48254 20018
rect 46174 19954 46226 19966
rect 48750 19954 48802 19966
rect 16830 19906 16882 19918
rect 4610 19854 4622 19906
rect 4674 19854 4686 19906
rect 6738 19854 6750 19906
rect 6802 19854 6814 19906
rect 15362 19854 15374 19906
rect 15426 19854 15438 19906
rect 16830 19842 16882 19854
rect 17502 19906 17554 19918
rect 17502 19842 17554 19854
rect 18062 19906 18114 19918
rect 18062 19842 18114 19854
rect 18734 19906 18786 19918
rect 22766 19906 22818 19918
rect 19058 19854 19070 19906
rect 19122 19854 19134 19906
rect 21186 19854 21198 19906
rect 21250 19854 21262 19906
rect 18734 19842 18786 19854
rect 22766 19842 22818 19854
rect 23662 19906 23714 19918
rect 31166 19906 31218 19918
rect 27346 19854 27358 19906
rect 27410 19854 27422 19906
rect 23662 19842 23714 19854
rect 31166 19842 31218 19854
rect 31614 19906 31666 19918
rect 31614 19842 31666 19854
rect 32062 19906 32114 19918
rect 32062 19842 32114 19854
rect 32510 19906 32562 19918
rect 32510 19842 32562 19854
rect 33182 19906 33234 19918
rect 45614 19906 45666 19918
rect 40114 19854 40126 19906
rect 40178 19854 40190 19906
rect 42242 19854 42254 19906
rect 42306 19854 42318 19906
rect 33182 19842 33234 19854
rect 45614 19842 45666 19854
rect 13582 19794 13634 19806
rect 16718 19794 16770 19806
rect 13906 19742 13918 19794
rect 13970 19742 13982 19794
rect 13582 19730 13634 19742
rect 16718 19730 16770 19742
rect 17838 19794 17890 19806
rect 17838 19730 17890 19742
rect 31054 19794 31106 19806
rect 33842 19742 33854 19794
rect 33906 19742 33918 19794
rect 31054 19730 31106 19742
rect 1344 19626 49616 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 49616 19626
rect 1344 19540 49616 19574
rect 25666 19406 25678 19458
rect 25730 19406 25742 19458
rect 21422 19346 21474 19358
rect 4610 19294 4622 19346
rect 4674 19294 4686 19346
rect 18386 19294 18398 19346
rect 18450 19294 18462 19346
rect 21422 19282 21474 19294
rect 25006 19346 25058 19358
rect 30494 19346 30546 19358
rect 28242 19294 28254 19346
rect 28306 19294 28318 19346
rect 29698 19294 29710 19346
rect 29762 19294 29774 19346
rect 25006 19282 25058 19294
rect 30494 19282 30546 19294
rect 31278 19346 31330 19358
rect 34290 19294 34302 19346
rect 34354 19294 34366 19346
rect 36418 19294 36430 19346
rect 36482 19294 36494 19346
rect 42914 19294 42926 19346
rect 42978 19294 42990 19346
rect 45042 19294 45054 19346
rect 45106 19294 45118 19346
rect 47058 19294 47070 19346
rect 47122 19294 47134 19346
rect 49186 19294 49198 19346
rect 49250 19294 49262 19346
rect 31278 19282 31330 19294
rect 7422 19234 7474 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 7422 19170 7474 19182
rect 8318 19234 8370 19246
rect 8318 19170 8370 19182
rect 8542 19234 8594 19246
rect 8542 19170 8594 19182
rect 8990 19234 9042 19246
rect 8990 19170 9042 19182
rect 13694 19234 13746 19246
rect 13694 19170 13746 19182
rect 14030 19234 14082 19246
rect 14030 19170 14082 19182
rect 14702 19234 14754 19246
rect 14702 19170 14754 19182
rect 14814 19234 14866 19246
rect 14814 19170 14866 19182
rect 14926 19234 14978 19246
rect 21310 19234 21362 19246
rect 20066 19182 20078 19234
rect 20130 19182 20142 19234
rect 14926 19170 14978 19182
rect 21310 19170 21362 19182
rect 21534 19234 21586 19246
rect 22094 19234 22146 19246
rect 22766 19234 22818 19246
rect 23998 19234 24050 19246
rect 21858 19182 21870 19234
rect 21922 19182 21934 19234
rect 22418 19182 22430 19234
rect 22482 19182 22494 19234
rect 23202 19182 23214 19234
rect 23266 19182 23278 19234
rect 21534 19170 21586 19182
rect 22094 19170 22146 19182
rect 22766 19170 22818 19182
rect 23998 19170 24050 19182
rect 26126 19234 26178 19246
rect 26126 19170 26178 19182
rect 26238 19234 26290 19246
rect 26798 19234 26850 19246
rect 29598 19234 29650 19246
rect 30606 19234 30658 19246
rect 26450 19182 26462 19234
rect 26514 19182 26526 19234
rect 27234 19182 27246 19234
rect 27298 19182 27310 19234
rect 27906 19182 27918 19234
rect 27970 19182 27982 19234
rect 29138 19182 29150 19234
rect 29202 19182 29214 19234
rect 30146 19182 30158 19234
rect 30210 19182 30222 19234
rect 26238 19170 26290 19182
rect 26798 19170 26850 19182
rect 29598 19170 29650 19182
rect 30606 19170 30658 19182
rect 32622 19234 32674 19246
rect 43038 19234 43090 19246
rect 33618 19182 33630 19234
rect 33682 19182 33694 19234
rect 41906 19182 41918 19234
rect 41970 19182 41982 19234
rect 32622 19170 32674 19182
rect 43038 19170 43090 19182
rect 43262 19234 43314 19246
rect 43262 19170 43314 19182
rect 44046 19234 44098 19246
rect 45490 19182 45502 19234
rect 45554 19182 45566 19234
rect 46274 19182 46286 19234
rect 46338 19182 46350 19234
rect 44046 19170 44098 19182
rect 5630 19122 5682 19134
rect 2482 19070 2494 19122
rect 2546 19070 2558 19122
rect 5630 19058 5682 19070
rect 5854 19122 5906 19134
rect 5854 19058 5906 19070
rect 6190 19122 6242 19134
rect 6190 19058 6242 19070
rect 6414 19122 6466 19134
rect 6414 19058 6466 19070
rect 6638 19122 6690 19134
rect 6638 19058 6690 19070
rect 6750 19122 6802 19134
rect 6750 19058 6802 19070
rect 7646 19122 7698 19134
rect 7646 19058 7698 19070
rect 7758 19122 7810 19134
rect 7758 19058 7810 19070
rect 9326 19122 9378 19134
rect 9326 19058 9378 19070
rect 9438 19122 9490 19134
rect 9438 19058 9490 19070
rect 12126 19122 12178 19134
rect 12126 19058 12178 19070
rect 13806 19122 13858 19134
rect 23662 19122 23714 19134
rect 22978 19070 22990 19122
rect 23042 19070 23054 19122
rect 13806 19058 13858 19070
rect 23662 19058 23714 19070
rect 25342 19122 25394 19134
rect 30830 19122 30882 19134
rect 28242 19070 28254 19122
rect 28306 19070 28318 19122
rect 25342 19058 25394 19070
rect 30830 19058 30882 19070
rect 31166 19122 31218 19134
rect 31166 19058 31218 19070
rect 31390 19122 31442 19134
rect 31390 19058 31442 19070
rect 33070 19122 33122 19134
rect 43486 19122 43538 19134
rect 39554 19070 39566 19122
rect 39618 19070 39630 19122
rect 33070 19058 33122 19070
rect 43486 19058 43538 19070
rect 45950 19122 46002 19134
rect 45950 19058 46002 19070
rect 5966 19010 6018 19022
rect 5966 18946 6018 18958
rect 8654 19010 8706 19022
rect 8654 18946 8706 18958
rect 9102 19010 9154 19022
rect 9102 18946 9154 18958
rect 9998 19010 10050 19022
rect 9998 18946 10050 18958
rect 11790 19010 11842 19022
rect 11790 18946 11842 18958
rect 12686 19010 12738 19022
rect 22206 19010 22258 19022
rect 14242 18958 14254 19010
rect 14306 18958 14318 19010
rect 12686 18946 12738 18958
rect 22206 18946 22258 18958
rect 24446 19010 24498 19022
rect 24446 18946 24498 18958
rect 29374 19010 29426 19022
rect 29374 18946 29426 18958
rect 29710 19010 29762 19022
rect 29710 18946 29762 18958
rect 30382 19010 30434 19022
rect 32174 19010 32226 19022
rect 31826 18958 31838 19010
rect 31890 18958 31902 19010
rect 30382 18946 30434 18958
rect 32174 18946 32226 18958
rect 33182 19010 33234 19022
rect 33182 18946 33234 18958
rect 42926 19010 42978 19022
rect 42926 18946 42978 18958
rect 44158 19010 44210 19022
rect 44158 18946 44210 18958
rect 44382 19010 44434 19022
rect 44382 18946 44434 18958
rect 1344 18842 49616 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 49616 18842
rect 1344 18756 49616 18790
rect 5070 18674 5122 18686
rect 5070 18610 5122 18622
rect 5294 18674 5346 18686
rect 16606 18674 16658 18686
rect 6626 18622 6638 18674
rect 6690 18622 6702 18674
rect 14242 18622 14254 18674
rect 14306 18622 14318 18674
rect 5294 18610 5346 18622
rect 16606 18610 16658 18622
rect 17390 18674 17442 18686
rect 17390 18610 17442 18622
rect 17614 18674 17666 18686
rect 17614 18610 17666 18622
rect 19406 18674 19458 18686
rect 19406 18610 19458 18622
rect 21086 18674 21138 18686
rect 21086 18610 21138 18622
rect 31390 18674 31442 18686
rect 31390 18610 31442 18622
rect 41022 18674 41074 18686
rect 48738 18622 48750 18674
rect 48802 18622 48814 18674
rect 41022 18610 41074 18622
rect 2494 18562 2546 18574
rect 2494 18498 2546 18510
rect 2606 18562 2658 18574
rect 2606 18498 2658 18510
rect 2942 18562 2994 18574
rect 2942 18498 2994 18510
rect 3054 18562 3106 18574
rect 3054 18498 3106 18510
rect 3278 18562 3330 18574
rect 3278 18498 3330 18510
rect 4510 18562 4562 18574
rect 4510 18498 4562 18510
rect 4622 18562 4674 18574
rect 4622 18498 4674 18510
rect 4958 18562 5010 18574
rect 4958 18498 5010 18510
rect 5518 18562 5570 18574
rect 8318 18562 8370 18574
rect 7746 18510 7758 18562
rect 7810 18510 7822 18562
rect 5518 18498 5570 18510
rect 8318 18498 8370 18510
rect 8542 18562 8594 18574
rect 8542 18498 8594 18510
rect 9662 18562 9714 18574
rect 9662 18498 9714 18510
rect 9774 18562 9826 18574
rect 17726 18562 17778 18574
rect 11778 18510 11790 18562
rect 11842 18510 11854 18562
rect 9774 18498 9826 18510
rect 17726 18498 17778 18510
rect 18510 18562 18562 18574
rect 18510 18498 18562 18510
rect 18622 18562 18674 18574
rect 18622 18498 18674 18510
rect 19182 18562 19234 18574
rect 19182 18498 19234 18510
rect 31278 18562 31330 18574
rect 42590 18562 42642 18574
rect 32050 18510 32062 18562
rect 32114 18510 32126 18562
rect 37538 18510 37550 18562
rect 37602 18510 37614 18562
rect 38658 18510 38670 18562
rect 38722 18510 38734 18562
rect 31278 18498 31330 18510
rect 42590 18498 42642 18510
rect 46510 18562 46562 18574
rect 46510 18498 46562 18510
rect 47518 18562 47570 18574
rect 47518 18498 47570 18510
rect 2270 18450 2322 18462
rect 2270 18386 2322 18398
rect 3390 18450 3442 18462
rect 3390 18386 3442 18398
rect 3726 18450 3778 18462
rect 3726 18386 3778 18398
rect 3950 18450 4002 18462
rect 3950 18386 4002 18398
rect 5854 18450 5906 18462
rect 7422 18450 7474 18462
rect 6850 18398 6862 18450
rect 6914 18398 6926 18450
rect 5854 18386 5906 18398
rect 7422 18386 7474 18398
rect 8990 18450 9042 18462
rect 8990 18386 9042 18398
rect 9438 18450 9490 18462
rect 14590 18450 14642 18462
rect 11106 18398 11118 18450
rect 11170 18398 11182 18450
rect 9438 18386 9490 18398
rect 14590 18386 14642 18398
rect 14814 18450 14866 18462
rect 14814 18386 14866 18398
rect 15262 18450 15314 18462
rect 15262 18386 15314 18398
rect 15374 18450 15426 18462
rect 15374 18386 15426 18398
rect 15598 18450 15650 18462
rect 16270 18450 16322 18462
rect 15810 18398 15822 18450
rect 15874 18398 15886 18450
rect 15598 18386 15650 18398
rect 16270 18386 16322 18398
rect 16382 18450 16434 18462
rect 16382 18386 16434 18398
rect 16494 18450 16546 18462
rect 19294 18450 19346 18462
rect 25342 18450 25394 18462
rect 16818 18398 16830 18450
rect 16882 18398 16894 18450
rect 18050 18398 18062 18450
rect 18114 18398 18126 18450
rect 19730 18398 19742 18450
rect 19794 18398 19806 18450
rect 24210 18398 24222 18450
rect 24274 18398 24286 18450
rect 16494 18386 16546 18398
rect 19294 18386 19346 18398
rect 25342 18386 25394 18398
rect 25790 18450 25842 18462
rect 30718 18450 30770 18462
rect 27346 18398 27358 18450
rect 27410 18398 27422 18450
rect 28018 18398 28030 18450
rect 28082 18398 28094 18450
rect 25790 18386 25842 18398
rect 30718 18386 30770 18398
rect 31166 18450 31218 18462
rect 31166 18386 31218 18398
rect 31502 18450 31554 18462
rect 36430 18450 36482 18462
rect 40910 18450 40962 18462
rect 42030 18450 42082 18462
rect 31714 18398 31726 18450
rect 31778 18398 31790 18450
rect 32274 18398 32286 18450
rect 32338 18398 32350 18450
rect 33282 18398 33294 18450
rect 33346 18398 33358 18450
rect 33954 18398 33966 18450
rect 34018 18398 34030 18450
rect 36978 18398 36990 18450
rect 37042 18398 37054 18450
rect 40226 18398 40238 18450
rect 40290 18398 40302 18450
rect 41122 18398 41134 18450
rect 41186 18398 41198 18450
rect 46162 18398 46174 18450
rect 46226 18398 46238 18450
rect 46722 18398 46734 18450
rect 46786 18398 46798 18450
rect 47954 18398 47966 18450
rect 48018 18398 48030 18450
rect 48962 18398 48974 18450
rect 49026 18398 49038 18450
rect 31502 18386 31554 18398
rect 36430 18386 36482 18398
rect 40910 18386 40962 18398
rect 42030 18386 42082 18398
rect 3614 18338 3666 18350
rect 3614 18274 3666 18286
rect 8766 18338 8818 18350
rect 8766 18274 8818 18286
rect 10222 18338 10274 18350
rect 10222 18274 10274 18286
rect 10670 18338 10722 18350
rect 20190 18338 20242 18350
rect 24670 18338 24722 18350
rect 13906 18286 13918 18338
rect 13970 18286 13982 18338
rect 15698 18286 15710 18338
rect 15762 18286 15774 18338
rect 18162 18286 18174 18338
rect 18226 18286 18238 18338
rect 21298 18286 21310 18338
rect 21362 18286 21374 18338
rect 23426 18286 23438 18338
rect 23490 18286 23502 18338
rect 10670 18274 10722 18286
rect 20190 18274 20242 18286
rect 24670 18274 24722 18286
rect 26462 18338 26514 18350
rect 26462 18274 26514 18286
rect 26574 18338 26626 18350
rect 30606 18338 30658 18350
rect 42142 18338 42194 18350
rect 30146 18286 30158 18338
rect 30210 18286 30222 18338
rect 36082 18286 36094 18338
rect 36146 18286 36158 18338
rect 26574 18274 26626 18286
rect 30606 18274 30658 18286
rect 42142 18274 42194 18286
rect 42478 18338 42530 18350
rect 43250 18286 43262 18338
rect 43314 18286 43326 18338
rect 45378 18286 45390 18338
rect 45442 18286 45454 18338
rect 42478 18274 42530 18286
rect 4510 18226 4562 18238
rect 18622 18226 18674 18238
rect 9986 18174 9998 18226
rect 10050 18223 10062 18226
rect 10658 18223 10670 18226
rect 10050 18177 10670 18223
rect 10050 18174 10062 18177
rect 10658 18174 10670 18177
rect 10722 18174 10734 18226
rect 4510 18162 4562 18174
rect 18622 18162 18674 18174
rect 20078 18226 20130 18238
rect 20078 18162 20130 18174
rect 25230 18226 25282 18238
rect 25230 18162 25282 18174
rect 25678 18226 25730 18238
rect 25678 18162 25730 18174
rect 36542 18226 36594 18238
rect 36542 18162 36594 18174
rect 37102 18226 37154 18238
rect 47058 18174 47070 18226
rect 47122 18174 47134 18226
rect 37102 18162 37154 18174
rect 1344 18058 49616 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 49616 18058
rect 1344 17972 49616 18006
rect 19070 17890 19122 17902
rect 19070 17826 19122 17838
rect 33182 17890 33234 17902
rect 33182 17826 33234 17838
rect 44942 17890 44994 17902
rect 44942 17826 44994 17838
rect 19406 17778 19458 17790
rect 4610 17726 4622 17778
rect 4674 17726 4686 17778
rect 8642 17726 8654 17778
rect 8706 17726 8718 17778
rect 10770 17726 10782 17778
rect 10834 17726 10846 17778
rect 13682 17726 13694 17778
rect 13746 17726 13758 17778
rect 19406 17714 19458 17726
rect 19630 17778 19682 17790
rect 19630 17714 19682 17726
rect 21422 17778 21474 17790
rect 21422 17714 21474 17726
rect 22206 17778 22258 17790
rect 27694 17778 27746 17790
rect 26898 17726 26910 17778
rect 26962 17726 26974 17778
rect 22206 17714 22258 17726
rect 27694 17714 27746 17726
rect 28366 17778 28418 17790
rect 28366 17714 28418 17726
rect 29262 17778 29314 17790
rect 42926 17778 42978 17790
rect 30706 17726 30718 17778
rect 30770 17726 30782 17778
rect 32834 17726 32846 17778
rect 32898 17726 32910 17778
rect 33954 17726 33966 17778
rect 34018 17726 34030 17778
rect 37090 17726 37102 17778
rect 37154 17726 37166 17778
rect 40338 17726 40350 17778
rect 40402 17726 40414 17778
rect 42466 17726 42478 17778
rect 42530 17726 42542 17778
rect 29262 17714 29314 17726
rect 42926 17714 42978 17726
rect 43374 17778 43426 17790
rect 44830 17778 44882 17790
rect 43810 17726 43822 17778
rect 43874 17726 43886 17778
rect 49186 17726 49198 17778
rect 49250 17726 49262 17778
rect 43374 17714 43426 17726
rect 44830 17714 44882 17726
rect 6302 17666 6354 17678
rect 20190 17666 20242 17678
rect 1810 17614 1822 17666
rect 1874 17614 1886 17666
rect 7970 17614 7982 17666
rect 8034 17614 8046 17666
rect 12674 17614 12686 17666
rect 12738 17614 12750 17666
rect 18386 17614 18398 17666
rect 18450 17614 18462 17666
rect 6302 17602 6354 17614
rect 20190 17602 20242 17614
rect 20414 17666 20466 17678
rect 20414 17602 20466 17614
rect 20862 17666 20914 17678
rect 20862 17602 20914 17614
rect 22094 17666 22146 17678
rect 22094 17602 22146 17614
rect 22318 17666 22370 17678
rect 22878 17666 22930 17678
rect 27582 17666 27634 17678
rect 34078 17666 34130 17678
rect 38334 17666 38386 17678
rect 22642 17614 22654 17666
rect 22706 17614 22718 17666
rect 23202 17614 23214 17666
rect 23266 17614 23278 17666
rect 24098 17614 24110 17666
rect 24162 17614 24174 17666
rect 24770 17614 24782 17666
rect 24834 17614 24846 17666
rect 28018 17614 28030 17666
rect 28082 17614 28094 17666
rect 30034 17614 30046 17666
rect 30098 17614 30110 17666
rect 33506 17614 33518 17666
rect 33570 17614 33582 17666
rect 33842 17614 33854 17666
rect 33906 17614 33918 17666
rect 34514 17614 34526 17666
rect 34578 17614 34590 17666
rect 37314 17614 37326 17666
rect 37378 17614 37390 17666
rect 37538 17614 37550 17666
rect 37602 17614 37614 17666
rect 22318 17602 22370 17614
rect 22878 17602 22930 17614
rect 27582 17602 27634 17614
rect 34078 17602 34130 17614
rect 38334 17602 38386 17614
rect 38446 17666 38498 17678
rect 38446 17602 38498 17614
rect 38894 17666 38946 17678
rect 38894 17602 38946 17614
rect 39006 17666 39058 17678
rect 45502 17666 45554 17678
rect 39554 17614 39566 17666
rect 39618 17614 39630 17666
rect 44146 17614 44158 17666
rect 44210 17614 44222 17666
rect 39006 17602 39058 17614
rect 45502 17602 45554 17614
rect 45726 17666 45778 17678
rect 46274 17614 46286 17666
rect 46338 17614 46350 17666
rect 45726 17602 45778 17614
rect 6862 17554 6914 17566
rect 2482 17502 2494 17554
rect 2546 17502 2558 17554
rect 6862 17490 6914 17502
rect 7198 17554 7250 17566
rect 7198 17490 7250 17502
rect 7534 17554 7586 17566
rect 7534 17490 7586 17502
rect 11118 17554 11170 17566
rect 11118 17490 11170 17502
rect 11902 17554 11954 17566
rect 11902 17490 11954 17502
rect 21310 17554 21362 17566
rect 21310 17490 21362 17502
rect 23438 17554 23490 17566
rect 23438 17490 23490 17502
rect 27358 17554 27410 17566
rect 27358 17490 27410 17502
rect 28478 17554 28530 17566
rect 28478 17490 28530 17502
rect 33294 17554 33346 17566
rect 33294 17490 33346 17502
rect 34302 17554 34354 17566
rect 45278 17554 45330 17566
rect 35410 17502 35422 17554
rect 35474 17502 35486 17554
rect 36082 17502 36094 17554
rect 36146 17502 36158 17554
rect 47058 17502 47070 17554
rect 47122 17502 47134 17554
rect 34302 17490 34354 17502
rect 45278 17490 45330 17502
rect 6526 17442 6578 17454
rect 5954 17390 5966 17442
rect 6018 17390 6030 17442
rect 6526 17378 6578 17390
rect 6750 17442 6802 17454
rect 6750 17378 6802 17390
rect 11230 17442 11282 17454
rect 11230 17378 11282 17390
rect 11454 17442 11506 17454
rect 11454 17378 11506 17390
rect 11566 17442 11618 17454
rect 11566 17378 11618 17390
rect 11790 17442 11842 17454
rect 11790 17378 11842 17390
rect 12910 17442 12962 17454
rect 12910 17378 12962 17390
rect 20302 17442 20354 17454
rect 20302 17378 20354 17390
rect 21534 17442 21586 17454
rect 21534 17378 21586 17390
rect 21758 17442 21810 17454
rect 21758 17378 21810 17390
rect 22990 17442 23042 17454
rect 22990 17378 23042 17390
rect 27806 17442 27858 17454
rect 27806 17378 27858 17390
rect 35086 17442 35138 17454
rect 35086 17378 35138 17390
rect 35758 17442 35810 17454
rect 35758 17378 35810 17390
rect 39118 17442 39170 17454
rect 39118 17378 39170 17390
rect 45614 17442 45666 17454
rect 45614 17378 45666 17390
rect 45838 17442 45890 17454
rect 45838 17378 45890 17390
rect 1344 17274 49616 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 49616 17274
rect 1344 17188 49616 17222
rect 9662 17106 9714 17118
rect 9662 17042 9714 17054
rect 16718 17106 16770 17118
rect 16718 17042 16770 17054
rect 17838 17106 17890 17118
rect 17838 17042 17890 17054
rect 21422 17106 21474 17118
rect 23438 17106 23490 17118
rect 22306 17054 22318 17106
rect 22370 17054 22382 17106
rect 21422 17042 21474 17054
rect 23438 17042 23490 17054
rect 23886 17106 23938 17118
rect 23886 17042 23938 17054
rect 24334 17106 24386 17118
rect 24334 17042 24386 17054
rect 24782 17106 24834 17118
rect 24782 17042 24834 17054
rect 25454 17106 25506 17118
rect 25454 17042 25506 17054
rect 26238 17106 26290 17118
rect 26238 17042 26290 17054
rect 31726 17106 31778 17118
rect 31726 17042 31778 17054
rect 31838 17106 31890 17118
rect 31838 17042 31890 17054
rect 33406 17106 33458 17118
rect 33406 17042 33458 17054
rect 35534 17106 35586 17118
rect 35534 17042 35586 17054
rect 47966 17106 48018 17118
rect 47966 17042 48018 17054
rect 48862 17106 48914 17118
rect 48862 17042 48914 17054
rect 1710 16994 1762 17006
rect 1710 16930 1762 16942
rect 2270 16994 2322 17006
rect 9550 16994 9602 17006
rect 17726 16994 17778 17006
rect 21870 16994 21922 17006
rect 30270 16994 30322 17006
rect 2818 16942 2830 16994
rect 2882 16942 2894 16994
rect 14130 16942 14142 16994
rect 14194 16942 14206 16994
rect 20290 16942 20302 16994
rect 20354 16942 20366 16994
rect 27682 16942 27694 16994
rect 27746 16942 27758 16994
rect 2270 16930 2322 16942
rect 9550 16930 9602 16942
rect 17726 16930 17778 16942
rect 21870 16930 21922 16942
rect 30270 16930 30322 16942
rect 30942 16994 30994 17006
rect 30942 16930 30994 16942
rect 33518 16994 33570 17006
rect 33518 16930 33570 16942
rect 33966 16994 34018 17006
rect 33966 16930 34018 16942
rect 34078 16994 34130 17006
rect 34078 16930 34130 16942
rect 34526 16994 34578 17006
rect 34526 16930 34578 16942
rect 34638 16994 34690 17006
rect 34638 16930 34690 16942
rect 35086 16994 35138 17006
rect 35086 16930 35138 16942
rect 35758 16994 35810 17006
rect 35758 16930 35810 16942
rect 40910 16994 40962 17006
rect 49086 16994 49138 17006
rect 42130 16942 42142 16994
rect 42194 16942 42206 16994
rect 45378 16942 45390 16994
rect 45442 16942 45454 16994
rect 40910 16930 40962 16942
rect 49086 16930 49138 16942
rect 1934 16882 1986 16894
rect 8094 16882 8146 16894
rect 7858 16830 7870 16882
rect 7922 16830 7934 16882
rect 1934 16818 1986 16830
rect 8094 16818 8146 16830
rect 8542 16882 8594 16894
rect 8542 16818 8594 16830
rect 8654 16882 8706 16894
rect 8654 16818 8706 16830
rect 9886 16882 9938 16894
rect 16830 16882 16882 16894
rect 21646 16882 21698 16894
rect 26574 16882 26626 16894
rect 31502 16882 31554 16894
rect 12226 16830 12238 16882
rect 12290 16830 12302 16882
rect 13010 16830 13022 16882
rect 13074 16830 13086 16882
rect 13346 16830 13358 16882
rect 13410 16830 13422 16882
rect 21074 16830 21086 16882
rect 21138 16830 21150 16882
rect 22530 16830 22542 16882
rect 22594 16830 22606 16882
rect 27010 16830 27022 16882
rect 27074 16830 27086 16882
rect 9886 16818 9938 16830
rect 16830 16818 16882 16830
rect 21646 16818 21698 16830
rect 26574 16818 26626 16830
rect 31502 16818 31554 16830
rect 31614 16882 31666 16894
rect 36654 16882 36706 16894
rect 41022 16882 41074 16894
rect 32050 16830 32062 16882
rect 32114 16830 32126 16882
rect 36530 16830 36542 16882
rect 36594 16830 36606 16882
rect 36978 16830 36990 16882
rect 37042 16830 37054 16882
rect 40338 16830 40350 16882
rect 40402 16830 40414 16882
rect 41458 16830 41470 16882
rect 41522 16830 41534 16882
rect 44706 16830 44718 16882
rect 44770 16830 44782 16882
rect 31614 16818 31666 16830
rect 36654 16818 36706 16830
rect 41022 16818 41074 16830
rect 2158 16770 2210 16782
rect 2158 16706 2210 16718
rect 8318 16770 8370 16782
rect 21534 16770 21586 16782
rect 30158 16770 30210 16782
rect 10098 16718 10110 16770
rect 10162 16718 10174 16770
rect 16258 16718 16270 16770
rect 16322 16718 16334 16770
rect 18162 16718 18174 16770
rect 18226 16718 18238 16770
rect 29810 16718 29822 16770
rect 29874 16718 29886 16770
rect 8318 16706 8370 16718
rect 21534 16706 21586 16718
rect 30158 16706 30210 16718
rect 32398 16770 32450 16782
rect 37426 16718 37438 16770
rect 37490 16718 37502 16770
rect 39554 16718 39566 16770
rect 39618 16718 39630 16770
rect 44258 16718 44270 16770
rect 44322 16718 44334 16770
rect 47506 16718 47518 16770
rect 47570 16718 47582 16770
rect 47842 16718 47854 16770
rect 47906 16718 47918 16770
rect 48738 16718 48750 16770
rect 48802 16718 48814 16770
rect 32398 16706 32450 16718
rect 30830 16658 30882 16670
rect 30830 16594 30882 16606
rect 32510 16658 32562 16670
rect 32510 16594 32562 16606
rect 33406 16658 33458 16670
rect 33406 16594 33458 16606
rect 33966 16658 34018 16670
rect 33966 16594 34018 16606
rect 34526 16658 34578 16670
rect 34526 16594 34578 16606
rect 34974 16658 35026 16670
rect 34974 16594 35026 16606
rect 48190 16658 48242 16670
rect 48190 16594 48242 16606
rect 1344 16490 49616 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 49616 16490
rect 1344 16404 49616 16438
rect 9550 16322 9602 16334
rect 9550 16258 9602 16270
rect 9998 16322 10050 16334
rect 48190 16322 48242 16334
rect 37538 16270 37550 16322
rect 37602 16270 37614 16322
rect 9998 16258 10050 16270
rect 48190 16258 48242 16270
rect 11678 16210 11730 16222
rect 4610 16158 4622 16210
rect 4674 16158 4686 16210
rect 5954 16158 5966 16210
rect 6018 16158 6030 16210
rect 8082 16158 8094 16210
rect 8146 16158 8158 16210
rect 11678 16146 11730 16158
rect 17166 16210 17218 16222
rect 23550 16210 23602 16222
rect 27358 16210 27410 16222
rect 29150 16210 29202 16222
rect 17826 16158 17838 16210
rect 17890 16158 17902 16210
rect 19954 16158 19966 16210
rect 20018 16158 20030 16210
rect 21746 16158 21758 16210
rect 21810 16158 21822 16210
rect 24658 16158 24670 16210
rect 24722 16158 24734 16210
rect 26786 16158 26798 16210
rect 26850 16158 26862 16210
rect 28354 16158 28366 16210
rect 28418 16158 28430 16210
rect 17166 16146 17218 16158
rect 23550 16146 23602 16158
rect 27358 16146 27410 16158
rect 29150 16146 29202 16158
rect 30158 16210 30210 16222
rect 30158 16146 30210 16158
rect 30606 16210 30658 16222
rect 44270 16210 44322 16222
rect 48414 16210 48466 16222
rect 37202 16158 37214 16210
rect 37266 16158 37278 16210
rect 42354 16158 42366 16210
rect 42418 16158 42430 16210
rect 45938 16158 45950 16210
rect 46002 16158 46014 16210
rect 30606 16146 30658 16158
rect 44270 16146 44322 16158
rect 48414 16146 48466 16158
rect 9774 16098 9826 16110
rect 10894 16098 10946 16110
rect 11566 16098 11618 16110
rect 1810 16046 1822 16098
rect 1874 16046 1886 16098
rect 8866 16046 8878 16098
rect 8930 16046 8942 16098
rect 9314 16046 9326 16098
rect 9378 16046 9390 16098
rect 10658 16046 10670 16098
rect 10722 16046 10734 16098
rect 11218 16046 11230 16098
rect 11282 16046 11294 16098
rect 9774 16034 9826 16046
rect 10894 16034 10946 16046
rect 11566 16034 11618 16046
rect 11790 16098 11842 16110
rect 11790 16034 11842 16046
rect 13358 16098 13410 16110
rect 13358 16034 13410 16046
rect 13694 16098 13746 16110
rect 17278 16098 17330 16110
rect 16818 16046 16830 16098
rect 16882 16046 16894 16098
rect 13694 16034 13746 16046
rect 17278 16034 17330 16046
rect 17390 16098 17442 16110
rect 23102 16098 23154 16110
rect 38894 16098 38946 16110
rect 42702 16098 42754 16110
rect 48862 16098 48914 16110
rect 20738 16046 20750 16098
rect 20802 16046 20814 16098
rect 21298 16046 21310 16098
rect 21362 16046 21374 16098
rect 21522 16046 21534 16098
rect 21586 16046 21598 16098
rect 23986 16046 23998 16098
rect 24050 16046 24062 16098
rect 27458 16046 27470 16098
rect 27522 16046 27534 16098
rect 28018 16046 28030 16098
rect 28082 16046 28094 16098
rect 28242 16046 28254 16098
rect 28306 16046 28318 16098
rect 35298 16046 35310 16098
rect 35362 16046 35374 16098
rect 37314 16046 37326 16098
rect 37378 16046 37390 16098
rect 37538 16046 37550 16098
rect 37602 16046 37614 16098
rect 39442 16046 39454 16098
rect 39506 16046 39518 16098
rect 46274 16046 46286 16098
rect 46338 16046 46350 16098
rect 47058 16046 47070 16098
rect 47122 16046 47134 16098
rect 47282 16046 47294 16098
rect 47346 16046 47358 16098
rect 17390 16034 17442 16046
rect 23102 16034 23154 16046
rect 38894 16034 38946 16046
rect 42702 16034 42754 16046
rect 48862 16034 48914 16046
rect 10110 15986 10162 15998
rect 2482 15934 2494 15986
rect 2546 15934 2558 15986
rect 10110 15922 10162 15934
rect 10446 15986 10498 15998
rect 10446 15922 10498 15934
rect 12126 15986 12178 15998
rect 12126 15922 12178 15934
rect 12686 15986 12738 15998
rect 12686 15922 12738 15934
rect 12798 15986 12850 15998
rect 12798 15922 12850 15934
rect 13022 15986 13074 15998
rect 13022 15922 13074 15934
rect 14030 15986 14082 15998
rect 14030 15922 14082 15934
rect 15486 15986 15538 15998
rect 15486 15922 15538 15934
rect 15822 15986 15874 15998
rect 15822 15922 15874 15934
rect 16158 15986 16210 15998
rect 16158 15922 16210 15934
rect 21758 15986 21810 15998
rect 21758 15922 21810 15934
rect 22542 15986 22594 15998
rect 22542 15922 22594 15934
rect 27246 15986 27298 15998
rect 27246 15922 27298 15934
rect 27694 15986 27746 15998
rect 27694 15922 27746 15934
rect 28478 15986 28530 15998
rect 38558 15986 38610 15998
rect 33506 15934 33518 15986
rect 33570 15934 33582 15986
rect 28478 15922 28530 15934
rect 38558 15922 38610 15934
rect 39118 15986 39170 15998
rect 46846 15986 46898 15998
rect 40226 15934 40238 15986
rect 40290 15934 40302 15986
rect 42914 15934 42926 15986
rect 42978 15934 42990 15986
rect 43586 15934 43598 15986
rect 43650 15934 43662 15986
rect 39118 15922 39170 15934
rect 46846 15922 46898 15934
rect 48638 15986 48690 15998
rect 48638 15922 48690 15934
rect 10558 15874 10610 15886
rect 10558 15810 10610 15822
rect 13582 15874 13634 15886
rect 13582 15810 13634 15822
rect 14478 15874 14530 15886
rect 15150 15874 15202 15886
rect 14802 15822 14814 15874
rect 14866 15822 14878 15874
rect 14478 15810 14530 15822
rect 15150 15810 15202 15822
rect 17054 15874 17106 15886
rect 17054 15810 17106 15822
rect 22206 15874 22258 15886
rect 22206 15810 22258 15822
rect 29262 15874 29314 15886
rect 29262 15810 29314 15822
rect 38670 15874 38722 15886
rect 45054 15874 45106 15886
rect 42802 15822 42814 15874
rect 42866 15822 42878 15874
rect 38670 15810 38722 15822
rect 45054 15810 45106 15822
rect 48750 15874 48802 15886
rect 48750 15810 48802 15822
rect 1344 15706 49616 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 49616 15706
rect 1344 15620 49616 15654
rect 2046 15538 2098 15550
rect 2046 15474 2098 15486
rect 2270 15538 2322 15550
rect 2270 15474 2322 15486
rect 3390 15538 3442 15550
rect 7758 15538 7810 15550
rect 5618 15486 5630 15538
rect 5682 15486 5694 15538
rect 3390 15474 3442 15486
rect 7758 15474 7810 15486
rect 8654 15538 8706 15550
rect 8654 15474 8706 15486
rect 16718 15538 16770 15550
rect 16718 15474 16770 15486
rect 17614 15538 17666 15550
rect 17614 15474 17666 15486
rect 19406 15538 19458 15550
rect 19406 15474 19458 15486
rect 20078 15538 20130 15550
rect 20078 15474 20130 15486
rect 20526 15538 20578 15550
rect 21198 15538 21250 15550
rect 25790 15538 25842 15550
rect 20850 15486 20862 15538
rect 20914 15486 20926 15538
rect 24546 15486 24558 15538
rect 24610 15486 24622 15538
rect 20526 15474 20578 15486
rect 21198 15474 21250 15486
rect 25790 15474 25842 15486
rect 26126 15538 26178 15550
rect 26126 15474 26178 15486
rect 26462 15538 26514 15550
rect 26462 15474 26514 15486
rect 26686 15538 26738 15550
rect 38670 15538 38722 15550
rect 37874 15486 37886 15538
rect 37938 15486 37950 15538
rect 26686 15474 26738 15486
rect 38670 15474 38722 15486
rect 38894 15538 38946 15550
rect 38894 15474 38946 15486
rect 41470 15538 41522 15550
rect 41470 15474 41522 15486
rect 2382 15426 2434 15438
rect 2382 15362 2434 15374
rect 2830 15426 2882 15438
rect 6190 15426 6242 15438
rect 4274 15374 4286 15426
rect 4338 15374 4350 15426
rect 5730 15374 5742 15426
rect 5794 15374 5806 15426
rect 2830 15362 2882 15374
rect 6190 15362 6242 15374
rect 6974 15426 7026 15438
rect 6974 15362 7026 15374
rect 7086 15426 7138 15438
rect 8430 15426 8482 15438
rect 8082 15374 8094 15426
rect 8146 15374 8158 15426
rect 7086 15362 7138 15374
rect 8430 15362 8482 15374
rect 8766 15426 8818 15438
rect 8766 15362 8818 15374
rect 8990 15426 9042 15438
rect 8990 15362 9042 15374
rect 16606 15426 16658 15438
rect 32286 15426 32338 15438
rect 28242 15374 28254 15426
rect 28306 15374 28318 15426
rect 29586 15374 29598 15426
rect 29650 15374 29662 15426
rect 30594 15374 30606 15426
rect 30658 15374 30670 15426
rect 16606 15362 16658 15374
rect 32286 15362 32338 15374
rect 32398 15426 32450 15438
rect 32398 15362 32450 15374
rect 33182 15426 33234 15438
rect 33182 15362 33234 15374
rect 38558 15426 38610 15438
rect 38558 15362 38610 15374
rect 39230 15426 39282 15438
rect 39230 15362 39282 15374
rect 39342 15426 39394 15438
rect 39342 15362 39394 15374
rect 39678 15426 39730 15438
rect 39678 15362 39730 15374
rect 39902 15426 39954 15438
rect 41918 15426 41970 15438
rect 41122 15374 41134 15426
rect 41186 15374 41198 15426
rect 48850 15374 48862 15426
rect 48914 15374 48926 15426
rect 39902 15362 39954 15374
rect 41918 15362 41970 15374
rect 2606 15314 2658 15326
rect 2606 15250 2658 15262
rect 2942 15314 2994 15326
rect 2942 15250 2994 15262
rect 3278 15314 3330 15326
rect 3278 15250 3330 15262
rect 3614 15314 3666 15326
rect 3614 15250 3666 15262
rect 3838 15314 3890 15326
rect 6526 15314 6578 15326
rect 4162 15262 4174 15314
rect 4226 15262 4238 15314
rect 5842 15262 5854 15314
rect 5906 15262 5918 15314
rect 3838 15250 3890 15262
rect 6526 15250 6578 15262
rect 6750 15314 6802 15326
rect 15486 15314 15538 15326
rect 15026 15262 15038 15314
rect 15090 15262 15102 15314
rect 6750 15250 6802 15262
rect 15486 15250 15538 15262
rect 15710 15314 15762 15326
rect 15710 15250 15762 15262
rect 16046 15314 16098 15326
rect 16046 15250 16098 15262
rect 18062 15314 18114 15326
rect 18062 15250 18114 15262
rect 18398 15314 18450 15326
rect 27134 15314 27186 15326
rect 32622 15314 32674 15326
rect 37774 15314 37826 15326
rect 18834 15262 18846 15314
rect 18898 15262 18910 15314
rect 21634 15262 21646 15314
rect 21698 15262 21710 15314
rect 22306 15262 22318 15314
rect 22370 15262 22382 15314
rect 27570 15262 27582 15314
rect 27634 15262 27646 15314
rect 29026 15262 29038 15314
rect 29090 15262 29102 15314
rect 30818 15262 30830 15314
rect 30882 15262 30894 15314
rect 33506 15262 33518 15314
rect 33570 15262 33582 15314
rect 37538 15262 37550 15314
rect 37602 15262 37614 15314
rect 18398 15250 18450 15262
rect 27134 15250 27186 15262
rect 32622 15250 32674 15262
rect 37774 15250 37826 15262
rect 42030 15314 42082 15326
rect 42030 15250 42082 15262
rect 42142 15314 42194 15326
rect 43026 15262 43038 15314
rect 43090 15262 43102 15314
rect 49074 15262 49086 15314
rect 49138 15262 49150 15314
rect 42142 15250 42194 15262
rect 15822 15202 15874 15214
rect 10098 15150 10110 15202
rect 10162 15150 10174 15202
rect 15822 15138 15874 15150
rect 26574 15202 26626 15214
rect 26574 15138 26626 15150
rect 31838 15202 31890 15214
rect 31838 15138 31890 15150
rect 33070 15202 33122 15214
rect 34290 15150 34302 15202
rect 34354 15150 34366 15202
rect 36418 15150 36430 15202
rect 36482 15150 36494 15202
rect 37202 15150 37214 15202
rect 37266 15150 37278 15202
rect 40002 15150 40014 15202
rect 40066 15150 40078 15202
rect 46050 15150 46062 15202
rect 46114 15150 46126 15202
rect 33070 15138 33122 15150
rect 31950 15090 32002 15102
rect 17378 15038 17390 15090
rect 17442 15087 17454 15090
rect 18162 15087 18174 15090
rect 17442 15041 18174 15087
rect 17442 15038 17454 15041
rect 18162 15038 18174 15041
rect 18226 15038 18238 15090
rect 31950 15026 32002 15038
rect 39230 15090 39282 15102
rect 42578 15038 42590 15090
rect 42642 15038 42654 15090
rect 39230 15026 39282 15038
rect 1344 14922 49616 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 49616 14922
rect 1344 14836 49616 14870
rect 8654 14754 8706 14766
rect 8654 14690 8706 14702
rect 9214 14642 9266 14654
rect 13582 14642 13634 14654
rect 17278 14642 17330 14654
rect 4610 14590 4622 14642
rect 4674 14590 4686 14642
rect 12898 14590 12910 14642
rect 12962 14590 12974 14642
rect 14690 14590 14702 14642
rect 14754 14590 14766 14642
rect 16818 14590 16830 14642
rect 16882 14590 16894 14642
rect 9214 14578 9266 14590
rect 13582 14578 13634 14590
rect 17278 14578 17330 14590
rect 17950 14642 18002 14654
rect 17950 14578 18002 14590
rect 26910 14642 26962 14654
rect 26910 14578 26962 14590
rect 27918 14642 27970 14654
rect 36094 14642 36146 14654
rect 30034 14590 30046 14642
rect 30098 14590 30110 14642
rect 32162 14590 32174 14642
rect 32226 14590 32238 14642
rect 35522 14590 35534 14642
rect 35586 14590 35598 14642
rect 27918 14578 27970 14590
rect 36094 14578 36146 14590
rect 36430 14642 36482 14654
rect 38110 14642 38162 14654
rect 37426 14590 37438 14642
rect 37490 14590 37502 14642
rect 36430 14578 36482 14590
rect 38110 14578 38162 14590
rect 40798 14642 40850 14654
rect 44942 14642 44994 14654
rect 41346 14590 41358 14642
rect 41410 14590 41422 14642
rect 40798 14578 40850 14590
rect 44942 14578 44994 14590
rect 45502 14642 45554 14654
rect 49186 14590 49198 14642
rect 49250 14590 49262 14642
rect 45502 14578 45554 14590
rect 6862 14530 6914 14542
rect 9438 14530 9490 14542
rect 19854 14530 19906 14542
rect 1810 14478 1822 14530
rect 1874 14478 1886 14530
rect 8306 14478 8318 14530
rect 8370 14478 8382 14530
rect 10098 14478 10110 14530
rect 10162 14478 10174 14530
rect 13906 14478 13918 14530
rect 13970 14478 13982 14530
rect 6862 14466 6914 14478
rect 9438 14466 9490 14478
rect 19854 14466 19906 14478
rect 20078 14530 20130 14542
rect 20078 14466 20130 14478
rect 20414 14530 20466 14542
rect 28030 14530 28082 14542
rect 37998 14530 38050 14542
rect 25554 14478 25566 14530
rect 25618 14478 25630 14530
rect 28354 14478 28366 14530
rect 28418 14478 28430 14530
rect 29362 14478 29374 14530
rect 29426 14478 29438 14530
rect 32722 14478 32734 14530
rect 32786 14478 32798 14530
rect 37538 14478 37550 14530
rect 37602 14478 37614 14530
rect 20414 14466 20466 14478
rect 28030 14466 28082 14478
rect 37998 14466 38050 14478
rect 38222 14530 38274 14542
rect 38222 14466 38274 14478
rect 38558 14530 38610 14542
rect 38558 14466 38610 14478
rect 39006 14530 39058 14542
rect 39006 14466 39058 14478
rect 39118 14530 39170 14542
rect 39118 14466 39170 14478
rect 39566 14530 39618 14542
rect 45390 14530 45442 14542
rect 44258 14478 44270 14530
rect 44322 14478 44334 14530
rect 39566 14466 39618 14478
rect 45390 14466 45442 14478
rect 45726 14530 45778 14542
rect 45726 14466 45778 14478
rect 45950 14530 46002 14542
rect 46274 14478 46286 14530
rect 46338 14478 46350 14530
rect 45950 14466 46002 14478
rect 7086 14418 7138 14430
rect 2482 14366 2494 14418
rect 2546 14366 2558 14418
rect 7086 14354 7138 14366
rect 7198 14418 7250 14430
rect 7198 14354 7250 14366
rect 9550 14418 9602 14430
rect 27806 14418 27858 14430
rect 38894 14418 38946 14430
rect 10770 14366 10782 14418
rect 10834 14366 10846 14418
rect 23650 14366 23662 14418
rect 23714 14366 23726 14418
rect 33394 14366 33406 14418
rect 33458 14366 33470 14418
rect 37426 14366 37438 14418
rect 37490 14366 37502 14418
rect 43474 14366 43486 14418
rect 43538 14366 43550 14418
rect 47058 14366 47070 14418
rect 47122 14366 47134 14418
rect 9550 14354 9602 14366
rect 27806 14354 27858 14366
rect 38894 14354 38946 14366
rect 5966 14306 6018 14318
rect 6638 14306 6690 14318
rect 5618 14254 5630 14306
rect 5682 14254 5694 14306
rect 6290 14254 6302 14306
rect 6354 14254 6366 14306
rect 5966 14242 6018 14254
rect 6638 14242 6690 14254
rect 8094 14306 8146 14318
rect 8094 14242 8146 14254
rect 8542 14306 8594 14318
rect 8542 14242 8594 14254
rect 9774 14306 9826 14318
rect 9774 14242 9826 14254
rect 18174 14306 18226 14318
rect 19294 14306 19346 14318
rect 20750 14306 20802 14318
rect 18498 14254 18510 14306
rect 18562 14254 18574 14306
rect 19506 14254 19518 14306
rect 19570 14254 19582 14306
rect 18174 14242 18226 14254
rect 19294 14242 19346 14254
rect 20750 14242 20802 14254
rect 27470 14306 27522 14318
rect 27470 14242 27522 14254
rect 39790 14306 39842 14318
rect 39790 14242 39842 14254
rect 39902 14306 39954 14318
rect 39902 14242 39954 14254
rect 40014 14306 40066 14318
rect 40014 14242 40066 14254
rect 40238 14306 40290 14318
rect 40238 14242 40290 14254
rect 45054 14306 45106 14318
rect 45054 14242 45106 14254
rect 1344 14138 49616 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 49616 14138
rect 1344 14052 49616 14086
rect 3502 13970 3554 13982
rect 3502 13906 3554 13918
rect 6190 13970 6242 13982
rect 6190 13906 6242 13918
rect 6414 13970 6466 13982
rect 6414 13906 6466 13918
rect 7310 13970 7362 13982
rect 7310 13906 7362 13918
rect 8206 13970 8258 13982
rect 8206 13906 8258 13918
rect 9774 13970 9826 13982
rect 9774 13906 9826 13918
rect 9998 13970 10050 13982
rect 9998 13906 10050 13918
rect 10782 13970 10834 13982
rect 12574 13970 12626 13982
rect 11890 13918 11902 13970
rect 11954 13918 11966 13970
rect 10782 13906 10834 13918
rect 12574 13906 12626 13918
rect 12798 13970 12850 13982
rect 12798 13906 12850 13918
rect 16830 13970 16882 13982
rect 16830 13906 16882 13918
rect 23998 13970 24050 13982
rect 23998 13906 24050 13918
rect 24334 13970 24386 13982
rect 24334 13906 24386 13918
rect 26686 13970 26738 13982
rect 33518 13970 33570 13982
rect 27234 13918 27246 13970
rect 27298 13918 27310 13970
rect 26686 13906 26738 13918
rect 33518 13906 33570 13918
rect 34638 13970 34690 13982
rect 34638 13906 34690 13918
rect 34862 13970 34914 13982
rect 34862 13906 34914 13918
rect 35534 13970 35586 13982
rect 35534 13906 35586 13918
rect 41022 13970 41074 13982
rect 41022 13906 41074 13918
rect 41246 13970 41298 13982
rect 41246 13906 41298 13918
rect 41470 13970 41522 13982
rect 41470 13906 41522 13918
rect 42814 13970 42866 13982
rect 42814 13906 42866 13918
rect 46622 13970 46674 13982
rect 46622 13906 46674 13918
rect 48302 13970 48354 13982
rect 48302 13906 48354 13918
rect 3166 13858 3218 13870
rect 3166 13794 3218 13806
rect 3278 13858 3330 13870
rect 3278 13794 3330 13806
rect 3838 13858 3890 13870
rect 3838 13794 3890 13806
rect 4062 13858 4114 13870
rect 4062 13794 4114 13806
rect 4398 13858 4450 13870
rect 4398 13794 4450 13806
rect 4846 13858 4898 13870
rect 4846 13794 4898 13806
rect 5518 13858 5570 13870
rect 5518 13794 5570 13806
rect 5630 13858 5682 13870
rect 8318 13858 8370 13870
rect 6626 13806 6638 13858
rect 6690 13806 6702 13858
rect 5630 13794 5682 13806
rect 8318 13794 8370 13806
rect 10334 13858 10386 13870
rect 10334 13794 10386 13806
rect 11566 13858 11618 13870
rect 11566 13794 11618 13806
rect 12462 13858 12514 13870
rect 18622 13858 18674 13870
rect 33742 13858 33794 13870
rect 13906 13806 13918 13858
rect 13970 13806 13982 13858
rect 24658 13806 24670 13858
rect 24722 13806 24734 13858
rect 12462 13794 12514 13806
rect 18622 13794 18674 13806
rect 33742 13794 33794 13806
rect 39342 13858 39394 13870
rect 39342 13794 39394 13806
rect 39678 13858 39730 13870
rect 39678 13794 39730 13806
rect 40014 13858 40066 13870
rect 48862 13858 48914 13870
rect 46946 13806 46958 13858
rect 47010 13806 47022 13858
rect 47730 13806 47742 13858
rect 47794 13806 47806 13858
rect 40014 13794 40066 13806
rect 48862 13794 48914 13806
rect 48974 13858 49026 13870
rect 48974 13794 49026 13806
rect 3726 13746 3778 13758
rect 3726 13682 3778 13694
rect 4174 13746 4226 13758
rect 4174 13682 4226 13694
rect 4510 13746 4562 13758
rect 4510 13682 4562 13694
rect 5854 13746 5906 13758
rect 5854 13682 5906 13694
rect 6078 13746 6130 13758
rect 6078 13682 6130 13694
rect 6974 13746 7026 13758
rect 6974 13682 7026 13694
rect 7646 13746 7698 13758
rect 7646 13682 7698 13694
rect 7982 13746 8034 13758
rect 10558 13746 10610 13758
rect 8642 13694 8654 13746
rect 8706 13694 8718 13746
rect 7982 13682 8034 13694
rect 10558 13682 10610 13694
rect 10894 13746 10946 13758
rect 10894 13682 10946 13694
rect 11118 13746 11170 13758
rect 17278 13746 17330 13758
rect 13234 13694 13246 13746
rect 13298 13694 13310 13746
rect 11118 13682 11170 13694
rect 17278 13682 17330 13694
rect 17614 13746 17666 13758
rect 17614 13682 17666 13694
rect 17950 13746 18002 13758
rect 17950 13682 18002 13694
rect 19518 13746 19570 13758
rect 19518 13682 19570 13694
rect 19742 13746 19794 13758
rect 28814 13746 28866 13758
rect 32510 13746 32562 13758
rect 20066 13694 20078 13746
rect 20130 13694 20142 13746
rect 20402 13694 20414 13746
rect 20466 13694 20478 13746
rect 23762 13694 23774 13746
rect 23826 13694 23838 13746
rect 27010 13694 27022 13746
rect 27074 13694 27086 13746
rect 29250 13694 29262 13746
rect 29314 13694 29326 13746
rect 19742 13682 19794 13694
rect 28814 13682 28866 13694
rect 32510 13682 32562 13694
rect 33070 13746 33122 13758
rect 33070 13682 33122 13694
rect 33294 13746 33346 13758
rect 33294 13682 33346 13694
rect 34190 13746 34242 13758
rect 34190 13682 34242 13694
rect 34414 13746 34466 13758
rect 40238 13746 40290 13758
rect 35746 13694 35758 13746
rect 35810 13694 35822 13746
rect 39106 13694 39118 13746
rect 39170 13694 39182 13746
rect 34414 13682 34466 13694
rect 40238 13682 40290 13694
rect 41358 13746 41410 13758
rect 41358 13682 41410 13694
rect 41694 13746 41746 13758
rect 41694 13682 41746 13694
rect 42142 13746 42194 13758
rect 42142 13682 42194 13694
rect 42254 13746 42306 13758
rect 47518 13746 47570 13758
rect 43474 13694 43486 13746
rect 43538 13694 43550 13746
rect 42254 13682 42306 13694
rect 47518 13682 47570 13694
rect 48078 13746 48130 13758
rect 48078 13682 48130 13694
rect 48750 13746 48802 13758
rect 48750 13682 48802 13694
rect 8878 13634 8930 13646
rect 17502 13634 17554 13646
rect 16034 13582 16046 13634
rect 16098 13582 16110 13634
rect 8878 13570 8930 13582
rect 17502 13570 17554 13582
rect 19630 13634 19682 13646
rect 26014 13634 26066 13646
rect 21186 13582 21198 13634
rect 21250 13582 21262 13634
rect 23314 13582 23326 13634
rect 23378 13582 23390 13634
rect 19630 13570 19682 13582
rect 26014 13570 26066 13582
rect 28030 13634 28082 13646
rect 28030 13570 28082 13582
rect 28366 13634 28418 13646
rect 33630 13634 33682 13646
rect 29922 13582 29934 13634
rect 29986 13582 29998 13634
rect 32050 13582 32062 13634
rect 32114 13582 32126 13634
rect 28366 13570 28418 13582
rect 33630 13570 33682 13582
rect 34750 13634 34802 13646
rect 39790 13634 39842 13646
rect 36530 13582 36542 13634
rect 36594 13582 36606 13634
rect 38658 13582 38670 13634
rect 38722 13582 38734 13634
rect 34750 13570 34802 13582
rect 39790 13570 39842 13582
rect 41918 13634 41970 13646
rect 47294 13634 47346 13646
rect 44146 13582 44158 13634
rect 44210 13582 44222 13634
rect 46274 13582 46286 13634
rect 46338 13582 46350 13634
rect 41918 13570 41970 13582
rect 47294 13570 47346 13582
rect 8990 13522 9042 13534
rect 8990 13458 9042 13470
rect 18510 13522 18562 13534
rect 18510 13458 18562 13470
rect 18846 13522 18898 13534
rect 25790 13522 25842 13534
rect 42702 13522 42754 13534
rect 25442 13470 25454 13522
rect 25506 13470 25518 13522
rect 27906 13470 27918 13522
rect 27970 13519 27982 13522
rect 28354 13519 28366 13522
rect 27970 13473 28366 13519
rect 27970 13470 27982 13473
rect 28354 13470 28366 13473
rect 28418 13470 28430 13522
rect 18846 13458 18898 13470
rect 25790 13458 25842 13470
rect 42702 13458 42754 13470
rect 43038 13522 43090 13534
rect 43038 13458 43090 13470
rect 1344 13354 49616 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 49616 13354
rect 1344 13268 49616 13302
rect 21646 13186 21698 13198
rect 11330 13134 11342 13186
rect 11394 13134 11406 13186
rect 21646 13122 21698 13134
rect 32846 13186 32898 13198
rect 32846 13122 32898 13134
rect 45054 13186 45106 13198
rect 45054 13122 45106 13134
rect 45838 13186 45890 13198
rect 45838 13122 45890 13134
rect 11118 13074 11170 13086
rect 2482 13022 2494 13074
rect 2546 13022 2558 13074
rect 4610 13022 4622 13074
rect 4674 13022 4686 13074
rect 7634 13022 7646 13074
rect 7698 13022 7710 13074
rect 9762 13022 9774 13074
rect 9826 13022 9838 13074
rect 11118 13010 11170 13022
rect 11902 13074 11954 13086
rect 11902 13010 11954 13022
rect 14030 13074 14082 13086
rect 27246 13074 27298 13086
rect 33406 13074 33458 13086
rect 17266 13022 17278 13074
rect 17330 13022 17342 13074
rect 18498 13022 18510 13074
rect 18562 13022 18574 13074
rect 20626 13022 20638 13074
rect 20690 13022 20702 13074
rect 24434 13022 24446 13074
rect 24498 13022 24510 13074
rect 26562 13022 26574 13074
rect 26626 13022 26638 13074
rect 30258 13022 30270 13074
rect 30322 13022 30334 13074
rect 14030 13010 14082 13022
rect 27246 13010 27298 13022
rect 33406 13010 33458 13022
rect 36094 13074 36146 13086
rect 36094 13010 36146 13022
rect 36430 13074 36482 13086
rect 43150 13074 43202 13086
rect 39442 13022 39454 13074
rect 39506 13022 39518 13074
rect 41570 13022 41582 13074
rect 41634 13022 41646 13074
rect 42018 13022 42030 13074
rect 42082 13022 42094 13074
rect 36430 13010 36482 13022
rect 43150 13010 43202 13022
rect 45390 13074 45442 13086
rect 45390 13010 45442 13022
rect 5630 12962 5682 12974
rect 1810 12910 1822 12962
rect 1874 12910 1886 12962
rect 5630 12898 5682 12910
rect 5854 12962 5906 12974
rect 5854 12898 5906 12910
rect 6190 12962 6242 12974
rect 6190 12898 6242 12910
rect 6414 12962 6466 12974
rect 6414 12898 6466 12910
rect 7086 12962 7138 12974
rect 11678 12962 11730 12974
rect 10546 12910 10558 12962
rect 10610 12910 10622 12962
rect 7086 12898 7138 12910
rect 11678 12898 11730 12910
rect 12126 12962 12178 12974
rect 12126 12898 12178 12910
rect 12462 12962 12514 12974
rect 12462 12898 12514 12910
rect 12798 12962 12850 12974
rect 12798 12898 12850 12910
rect 13806 12962 13858 12974
rect 22990 12962 23042 12974
rect 29486 12962 29538 12974
rect 14354 12910 14366 12962
rect 14418 12910 14430 12962
rect 17714 12910 17726 12962
rect 17778 12910 17790 12962
rect 21634 12910 21646 12962
rect 21698 12910 21710 12962
rect 23650 12910 23662 12962
rect 23714 12910 23726 12962
rect 27682 12910 27694 12962
rect 27746 12910 27758 12962
rect 28578 12910 28590 12962
rect 28642 12910 28654 12962
rect 13806 12898 13858 12910
rect 22990 12898 23042 12910
rect 29486 12898 29538 12910
rect 29710 12962 29762 12974
rect 29710 12898 29762 12910
rect 29934 12962 29986 12974
rect 33070 12962 33122 12974
rect 30370 12910 30382 12962
rect 30434 12910 30446 12962
rect 31490 12910 31502 12962
rect 31554 12910 31566 12962
rect 32050 12910 32062 12962
rect 32114 12910 32126 12962
rect 29934 12898 29986 12910
rect 33070 12898 33122 12910
rect 33294 12962 33346 12974
rect 33294 12898 33346 12910
rect 33518 12962 33570 12974
rect 34862 12962 34914 12974
rect 34290 12910 34302 12962
rect 34354 12910 34366 12962
rect 33518 12898 33570 12910
rect 34862 12898 34914 12910
rect 36318 12962 36370 12974
rect 36318 12898 36370 12910
rect 37214 12962 37266 12974
rect 37214 12898 37266 12910
rect 37662 12962 37714 12974
rect 44046 12962 44098 12974
rect 38658 12910 38670 12962
rect 38722 12910 38734 12962
rect 42354 12910 42366 12962
rect 42418 12910 42430 12962
rect 42802 12910 42814 12962
rect 42866 12910 42878 12962
rect 43810 12910 43822 12962
rect 43874 12910 43886 12962
rect 37662 12898 37714 12910
rect 44046 12898 44098 12910
rect 46062 12962 46114 12974
rect 47518 12962 47570 12974
rect 46274 12910 46286 12962
rect 46338 12910 46350 12962
rect 47282 12910 47294 12962
rect 47346 12910 47358 12962
rect 46062 12898 46114 12910
rect 47518 12898 47570 12910
rect 48078 12962 48130 12974
rect 48078 12898 48130 12910
rect 48302 12962 48354 12974
rect 48302 12898 48354 12910
rect 49198 12962 49250 12974
rect 49198 12898 49250 12910
rect 6750 12850 6802 12862
rect 6750 12786 6802 12798
rect 7198 12850 7250 12862
rect 7198 12786 7250 12798
rect 12350 12850 12402 12862
rect 12350 12786 12402 12798
rect 12910 12850 12962 12862
rect 21982 12850 22034 12862
rect 15138 12798 15150 12850
rect 15202 12798 15214 12850
rect 12910 12786 12962 12798
rect 21982 12786 22034 12798
rect 22542 12850 22594 12862
rect 22542 12786 22594 12798
rect 22878 12850 22930 12862
rect 34974 12850 35026 12862
rect 27906 12798 27918 12850
rect 27970 12798 27982 12850
rect 30706 12798 30718 12850
rect 30770 12798 30782 12850
rect 31378 12798 31390 12850
rect 31442 12798 31454 12850
rect 22878 12786 22930 12798
rect 34974 12786 35026 12798
rect 35310 12850 35362 12862
rect 35310 12786 35362 12798
rect 35422 12850 35474 12862
rect 35422 12786 35474 12798
rect 36990 12850 37042 12862
rect 36990 12786 37042 12798
rect 46622 12850 46674 12862
rect 46622 12786 46674 12798
rect 48190 12850 48242 12862
rect 48190 12786 48242 12798
rect 49086 12850 49138 12862
rect 49086 12786 49138 12798
rect 5182 12738 5234 12750
rect 5182 12674 5234 12686
rect 5966 12738 6018 12750
rect 5966 12674 6018 12686
rect 6638 12738 6690 12750
rect 6638 12674 6690 12686
rect 7422 12738 7474 12750
rect 22766 12738 22818 12750
rect 13458 12686 13470 12738
rect 13522 12686 13534 12738
rect 7422 12674 7474 12686
rect 22766 12674 22818 12686
rect 23214 12738 23266 12750
rect 29262 12738 29314 12750
rect 28466 12686 28478 12738
rect 28530 12686 28542 12738
rect 23214 12674 23266 12686
rect 29262 12674 29314 12686
rect 29374 12738 29426 12750
rect 29374 12674 29426 12686
rect 35646 12738 35698 12750
rect 35646 12674 35698 12686
rect 37326 12738 37378 12750
rect 37326 12674 37378 12686
rect 37886 12738 37938 12750
rect 45166 12738 45218 12750
rect 38210 12686 38222 12738
rect 38274 12686 38286 12738
rect 37886 12674 37938 12686
rect 45166 12674 45218 12686
rect 46174 12738 46226 12750
rect 48738 12686 48750 12738
rect 48802 12686 48814 12738
rect 46174 12674 46226 12686
rect 1344 12570 49616 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 49616 12570
rect 1344 12484 49616 12518
rect 3502 12402 3554 12414
rect 3502 12338 3554 12350
rect 9550 12402 9602 12414
rect 9550 12338 9602 12350
rect 9662 12402 9714 12414
rect 9662 12338 9714 12350
rect 9774 12402 9826 12414
rect 9774 12338 9826 12350
rect 15822 12402 15874 12414
rect 15822 12338 15874 12350
rect 15934 12402 15986 12414
rect 15934 12338 15986 12350
rect 21086 12402 21138 12414
rect 21086 12338 21138 12350
rect 22430 12402 22482 12414
rect 24446 12402 24498 12414
rect 22754 12350 22766 12402
rect 22818 12350 22830 12402
rect 22430 12338 22482 12350
rect 24446 12338 24498 12350
rect 25454 12402 25506 12414
rect 25454 12338 25506 12350
rect 25678 12402 25730 12414
rect 25678 12338 25730 12350
rect 31838 12402 31890 12414
rect 31838 12338 31890 12350
rect 40014 12402 40066 12414
rect 40014 12338 40066 12350
rect 46510 12402 46562 12414
rect 46510 12338 46562 12350
rect 3390 12290 3442 12302
rect 3390 12226 3442 12238
rect 3726 12290 3778 12302
rect 3726 12226 3778 12238
rect 4510 12290 4562 12302
rect 4510 12226 4562 12238
rect 5630 12290 5682 12302
rect 5630 12226 5682 12238
rect 17950 12290 18002 12302
rect 17950 12226 18002 12238
rect 18062 12290 18114 12302
rect 18062 12226 18114 12238
rect 21422 12290 21474 12302
rect 21422 12226 21474 12238
rect 21758 12290 21810 12302
rect 30158 12290 30210 12302
rect 32398 12290 32450 12302
rect 22082 12238 22094 12290
rect 22146 12238 22158 12290
rect 31042 12238 31054 12290
rect 31106 12238 31118 12290
rect 21758 12226 21810 12238
rect 30158 12226 30210 12238
rect 32398 12226 32450 12238
rect 32510 12290 32562 12302
rect 42814 12290 42866 12302
rect 45838 12290 45890 12302
rect 35746 12238 35758 12290
rect 35810 12238 35822 12290
rect 45266 12238 45278 12290
rect 45330 12238 45342 12290
rect 32510 12226 32562 12238
rect 42814 12226 42866 12238
rect 45838 12226 45890 12238
rect 46734 12290 46786 12302
rect 46734 12226 46786 12238
rect 3838 12178 3890 12190
rect 3838 12114 3890 12126
rect 4286 12178 4338 12190
rect 5070 12178 5122 12190
rect 10222 12178 10274 12190
rect 14478 12178 14530 12190
rect 4834 12126 4846 12178
rect 4898 12126 4910 12178
rect 8754 12126 8766 12178
rect 8818 12126 8830 12178
rect 10770 12126 10782 12178
rect 10834 12126 10846 12178
rect 4286 12114 4338 12126
rect 5070 12114 5122 12126
rect 10222 12114 10274 12126
rect 14478 12114 14530 12126
rect 14814 12178 14866 12190
rect 14814 12114 14866 12126
rect 15038 12178 15090 12190
rect 15710 12178 15762 12190
rect 15362 12126 15374 12178
rect 15426 12126 15438 12178
rect 15038 12114 15090 12126
rect 15710 12114 15762 12126
rect 16382 12178 16434 12190
rect 16382 12114 16434 12126
rect 16606 12178 16658 12190
rect 16606 12114 16658 12126
rect 16718 12178 16770 12190
rect 17838 12178 17890 12190
rect 23102 12178 23154 12190
rect 17378 12126 17390 12178
rect 17442 12126 17454 12178
rect 19058 12126 19070 12178
rect 19122 12126 19134 12178
rect 19730 12126 19742 12178
rect 19794 12126 19806 12178
rect 16718 12114 16770 12126
rect 17838 12114 17890 12126
rect 23102 12114 23154 12126
rect 23326 12178 23378 12190
rect 23326 12114 23378 12126
rect 26126 12178 26178 12190
rect 26126 12114 26178 12126
rect 26462 12178 26514 12190
rect 39230 12178 39282 12190
rect 29698 12126 29710 12178
rect 29762 12126 29774 12178
rect 31154 12126 31166 12178
rect 31218 12126 31230 12178
rect 31602 12126 31614 12178
rect 31666 12126 31678 12178
rect 37090 12126 37102 12178
rect 37154 12126 37166 12178
rect 38770 12126 38782 12178
rect 38834 12126 38846 12178
rect 26462 12114 26514 12126
rect 39230 12114 39282 12126
rect 39566 12178 39618 12190
rect 39566 12114 39618 12126
rect 39790 12178 39842 12190
rect 39790 12114 39842 12126
rect 41246 12178 41298 12190
rect 41246 12114 41298 12126
rect 41470 12178 41522 12190
rect 41470 12114 41522 12126
rect 41694 12178 41746 12190
rect 41694 12114 41746 12126
rect 41918 12178 41970 12190
rect 41918 12114 41970 12126
rect 42478 12178 42530 12190
rect 42478 12114 42530 12126
rect 42702 12178 42754 12190
rect 42702 12114 42754 12126
rect 43262 12178 43314 12190
rect 43262 12114 43314 12126
rect 43486 12178 43538 12190
rect 43486 12114 43538 12126
rect 44942 12178 44994 12190
rect 44942 12114 44994 12126
rect 46062 12178 46114 12190
rect 47730 12126 47742 12178
rect 47794 12126 47806 12178
rect 49074 12126 49086 12178
rect 49138 12126 49150 12178
rect 46062 12114 46114 12126
rect 4062 12066 4114 12078
rect 14142 12066 14194 12078
rect 5954 12014 5966 12066
rect 6018 12014 6030 12066
rect 8082 12014 8094 12066
rect 8146 12014 8158 12066
rect 11554 12014 11566 12066
rect 11618 12014 11630 12066
rect 13682 12014 13694 12066
rect 13746 12014 13758 12066
rect 4062 12002 4114 12014
rect 14142 12002 14194 12014
rect 14590 12066 14642 12078
rect 14590 12002 14642 12014
rect 18846 12066 18898 12078
rect 18846 12002 18898 12014
rect 20302 12066 20354 12078
rect 20302 12002 20354 12014
rect 23998 12066 24050 12078
rect 24670 12066 24722 12078
rect 24434 12014 24446 12066
rect 24498 12014 24510 12066
rect 23998 12002 24050 12014
rect 24670 12002 24722 12014
rect 25566 12066 25618 12078
rect 39678 12066 39730 12078
rect 26786 12014 26798 12066
rect 26850 12014 26862 12066
rect 28914 12014 28926 12066
rect 28978 12014 28990 12066
rect 31266 12014 31278 12066
rect 31330 12014 31342 12066
rect 25566 12002 25618 12014
rect 39678 12002 39730 12014
rect 41022 12066 41074 12078
rect 41022 12002 41074 12014
rect 44046 12066 44098 12078
rect 44046 12002 44098 12014
rect 45950 12066 46002 12078
rect 47506 12014 47518 12066
rect 47570 12014 47582 12066
rect 45950 12002 46002 12014
rect 5294 11954 5346 11966
rect 5294 11890 5346 11902
rect 5518 11954 5570 11966
rect 5518 11890 5570 11902
rect 16270 11954 16322 11966
rect 16270 11890 16322 11902
rect 19070 11954 19122 11966
rect 19070 11890 19122 11902
rect 19406 11954 19458 11966
rect 19406 11890 19458 11902
rect 20078 11954 20130 11966
rect 20078 11890 20130 11902
rect 30270 11954 30322 11966
rect 30270 11890 30322 11902
rect 42366 11954 42418 11966
rect 42366 11890 42418 11902
rect 43150 11954 43202 11966
rect 43150 11890 43202 11902
rect 43598 11954 43650 11966
rect 43598 11890 43650 11902
rect 44270 11954 44322 11966
rect 46398 11954 46450 11966
rect 48750 11954 48802 11966
rect 44594 11902 44606 11954
rect 44658 11902 44670 11954
rect 47954 11902 47966 11954
rect 48018 11902 48030 11954
rect 44270 11890 44322 11902
rect 46398 11890 46450 11902
rect 48750 11890 48802 11902
rect 49086 11954 49138 11966
rect 49086 11890 49138 11902
rect 1344 11786 49616 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 49616 11786
rect 1344 11700 49616 11734
rect 49086 11618 49138 11630
rect 11330 11566 11342 11618
rect 11394 11615 11406 11618
rect 12338 11615 12350 11618
rect 11394 11569 12350 11615
rect 11394 11566 11406 11569
rect 12338 11566 12350 11569
rect 12402 11566 12414 11618
rect 44258 11566 44270 11618
rect 44322 11566 44334 11618
rect 49086 11554 49138 11566
rect 11342 11506 11394 11518
rect 2482 11454 2494 11506
rect 2546 11454 2558 11506
rect 4610 11454 4622 11506
rect 4674 11454 4686 11506
rect 8754 11454 8766 11506
rect 8818 11454 8830 11506
rect 11342 11442 11394 11454
rect 11790 11506 11842 11518
rect 11790 11442 11842 11454
rect 12238 11506 12290 11518
rect 12238 11442 12290 11454
rect 19182 11506 19234 11518
rect 19182 11442 19234 11454
rect 19854 11506 19906 11518
rect 19854 11442 19906 11454
rect 22430 11506 22482 11518
rect 22430 11442 22482 11454
rect 23326 11506 23378 11518
rect 48190 11506 48242 11518
rect 24434 11454 24446 11506
rect 24498 11454 24510 11506
rect 26562 11454 26574 11506
rect 26626 11454 26638 11506
rect 30930 11454 30942 11506
rect 30994 11454 31006 11506
rect 33058 11454 33070 11506
rect 33122 11454 33134 11506
rect 33506 11454 33518 11506
rect 33570 11454 33582 11506
rect 35634 11454 35646 11506
rect 35698 11454 35710 11506
rect 45602 11454 45614 11506
rect 45666 11454 45678 11506
rect 47730 11454 47742 11506
rect 47794 11454 47806 11506
rect 23326 11442 23378 11454
rect 48190 11442 48242 11454
rect 12910 11394 12962 11406
rect 19966 11394 20018 11406
rect 1810 11342 1822 11394
rect 1874 11342 1886 11394
rect 10770 11342 10782 11394
rect 10834 11342 10846 11394
rect 18274 11342 18286 11394
rect 18338 11342 18350 11394
rect 12910 11330 12962 11342
rect 19966 11330 20018 11342
rect 20414 11394 20466 11406
rect 28366 11394 28418 11406
rect 23650 11342 23662 11394
rect 23714 11342 23726 11394
rect 26898 11342 26910 11394
rect 26962 11342 26974 11394
rect 20414 11330 20466 11342
rect 28366 11330 28418 11342
rect 28590 11394 28642 11406
rect 28590 11330 28642 11342
rect 29150 11394 29202 11406
rect 36990 11394 37042 11406
rect 29586 11342 29598 11394
rect 29650 11342 29662 11394
rect 30258 11342 30270 11394
rect 30322 11342 30334 11394
rect 36418 11342 36430 11394
rect 36482 11342 36494 11394
rect 29150 11330 29202 11342
rect 36990 11330 37042 11342
rect 37550 11394 37602 11406
rect 47966 11394 48018 11406
rect 42914 11342 42926 11394
rect 42978 11342 42990 11394
rect 43474 11342 43486 11394
rect 43538 11342 43550 11394
rect 44818 11342 44830 11394
rect 44882 11342 44894 11394
rect 37550 11330 37602 11342
rect 47966 11330 48018 11342
rect 48302 11394 48354 11406
rect 48302 11330 48354 11342
rect 48638 11394 48690 11406
rect 48638 11330 48690 11342
rect 48974 11394 49026 11406
rect 48974 11330 49026 11342
rect 12574 11282 12626 11294
rect 20862 11282 20914 11294
rect 13682 11230 13694 11282
rect 13746 11230 13758 11282
rect 12574 11218 12626 11230
rect 20862 11218 20914 11230
rect 21646 11282 21698 11294
rect 43710 11282 43762 11294
rect 38098 11230 38110 11282
rect 38162 11230 38174 11282
rect 21646 11218 21698 11230
rect 43710 11218 43762 11230
rect 43822 11282 43874 11294
rect 43822 11218 43874 11230
rect 5070 11170 5122 11182
rect 5070 11106 5122 11118
rect 19742 11170 19794 11182
rect 19742 11106 19794 11118
rect 21982 11170 22034 11182
rect 21982 11106 22034 11118
rect 22990 11170 23042 11182
rect 22990 11106 23042 11118
rect 27246 11170 27298 11182
rect 27246 11106 27298 11118
rect 27358 11170 27410 11182
rect 27358 11106 27410 11118
rect 27470 11170 27522 11182
rect 49086 11170 49138 11182
rect 28018 11118 28030 11170
rect 28082 11118 28094 11170
rect 27470 11106 27522 11118
rect 49086 11106 49138 11118
rect 1344 11002 49616 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 49616 11002
rect 1344 10916 49616 10950
rect 5518 10834 5570 10846
rect 5518 10770 5570 10782
rect 5742 10834 5794 10846
rect 5742 10770 5794 10782
rect 6638 10834 6690 10846
rect 6638 10770 6690 10782
rect 9102 10834 9154 10846
rect 16718 10834 16770 10846
rect 10210 10782 10222 10834
rect 10274 10782 10286 10834
rect 9102 10770 9154 10782
rect 16718 10770 16770 10782
rect 16830 10834 16882 10846
rect 16830 10770 16882 10782
rect 20974 10834 21026 10846
rect 20974 10770 21026 10782
rect 31614 10834 31666 10846
rect 31614 10770 31666 10782
rect 31726 10834 31778 10846
rect 31726 10770 31778 10782
rect 31838 10834 31890 10846
rect 31838 10770 31890 10782
rect 32398 10834 32450 10846
rect 32398 10770 32450 10782
rect 37102 10834 37154 10846
rect 37102 10770 37154 10782
rect 42366 10834 42418 10846
rect 45826 10782 45838 10834
rect 45890 10782 45902 10834
rect 42366 10770 42418 10782
rect 5854 10722 5906 10734
rect 5854 10658 5906 10670
rect 6862 10722 6914 10734
rect 6862 10658 6914 10670
rect 7422 10722 7474 10734
rect 11790 10722 11842 10734
rect 32510 10722 32562 10734
rect 10882 10670 10894 10722
rect 10946 10670 10958 10722
rect 13794 10670 13806 10722
rect 13858 10670 13870 10722
rect 18386 10670 18398 10722
rect 18450 10670 18462 10722
rect 28802 10670 28814 10722
rect 28866 10670 28878 10722
rect 7422 10658 7474 10670
rect 11790 10658 11842 10670
rect 32510 10658 32562 10670
rect 34078 10722 34130 10734
rect 34078 10658 34130 10670
rect 34974 10722 35026 10734
rect 34974 10658 35026 10670
rect 35198 10722 35250 10734
rect 35198 10658 35250 10670
rect 36654 10722 36706 10734
rect 36654 10658 36706 10670
rect 41246 10722 41298 10734
rect 46734 10722 46786 10734
rect 44706 10670 44718 10722
rect 44770 10670 44782 10722
rect 41246 10658 41298 10670
rect 46734 10658 46786 10670
rect 47294 10722 47346 10734
rect 47294 10658 47346 10670
rect 48750 10722 48802 10734
rect 48750 10658 48802 10670
rect 48974 10722 49026 10734
rect 48974 10658 49026 10670
rect 6526 10610 6578 10622
rect 6526 10546 6578 10558
rect 6974 10610 7026 10622
rect 6974 10546 7026 10558
rect 7646 10610 7698 10622
rect 7646 10546 7698 10558
rect 10558 10610 10610 10622
rect 10558 10546 10610 10558
rect 11230 10610 11282 10622
rect 16158 10610 16210 10622
rect 13010 10558 13022 10610
rect 13074 10558 13086 10610
rect 11230 10546 11282 10558
rect 16158 10546 16210 10558
rect 16606 10610 16658 10622
rect 31166 10610 31218 10622
rect 17714 10558 17726 10610
rect 17778 10558 17790 10610
rect 21298 10558 21310 10610
rect 21362 10558 21374 10610
rect 25330 10558 25342 10610
rect 25394 10558 25406 10610
rect 29362 10558 29374 10610
rect 29426 10558 29438 10610
rect 30034 10558 30046 10610
rect 30098 10558 30110 10610
rect 16606 10546 16658 10558
rect 31166 10546 31218 10558
rect 31390 10610 31442 10622
rect 31390 10546 31442 10558
rect 32174 10610 32226 10622
rect 32174 10546 32226 10558
rect 33070 10610 33122 10622
rect 34414 10610 34466 10622
rect 33506 10558 33518 10610
rect 33570 10558 33582 10610
rect 33070 10546 33122 10558
rect 34414 10546 34466 10558
rect 34526 10610 34578 10622
rect 36094 10610 36146 10622
rect 35410 10558 35422 10610
rect 35474 10558 35486 10610
rect 35634 10558 35646 10610
rect 35698 10558 35710 10610
rect 34526 10546 34578 10558
rect 36094 10546 36146 10558
rect 36318 10610 36370 10622
rect 41918 10610 41970 10622
rect 37538 10558 37550 10610
rect 37602 10558 37614 10610
rect 45490 10558 45502 10610
rect 45554 10558 45566 10610
rect 46050 10558 46062 10610
rect 46114 10558 46126 10610
rect 48066 10558 48078 10610
rect 48130 10558 48142 10610
rect 36318 10546 36370 10558
rect 41918 10546 41970 10558
rect 5294 10498 5346 10510
rect 5294 10434 5346 10446
rect 7198 10498 7250 10510
rect 7198 10434 7250 10446
rect 7982 10498 8034 10510
rect 7982 10434 8034 10446
rect 9886 10498 9938 10510
rect 9886 10434 9938 10446
rect 12798 10498 12850 10510
rect 24670 10498 24722 10510
rect 30718 10498 30770 10510
rect 15922 10446 15934 10498
rect 15986 10446 15998 10498
rect 20514 10446 20526 10498
rect 20578 10446 20590 10498
rect 22082 10446 22094 10498
rect 22146 10446 22158 10498
rect 24210 10446 24222 10498
rect 24274 10446 24286 10498
rect 26002 10446 26014 10498
rect 26066 10446 26078 10498
rect 28130 10446 28142 10498
rect 28194 10446 28206 10498
rect 12798 10434 12850 10446
rect 24670 10434 24722 10446
rect 30718 10434 30770 10446
rect 34190 10498 34242 10510
rect 36542 10498 36594 10510
rect 47630 10498 47682 10510
rect 35746 10446 35758 10498
rect 35810 10446 35822 10498
rect 38210 10446 38222 10498
rect 38274 10446 38286 10498
rect 40338 10446 40350 10498
rect 40402 10446 40414 10498
rect 42578 10446 42590 10498
rect 42642 10446 42654 10498
rect 34190 10434 34242 10446
rect 36542 10434 36594 10446
rect 47630 10434 47682 10446
rect 48862 10498 48914 10510
rect 48862 10434 48914 10446
rect 8206 10386 8258 10398
rect 11566 10386 11618 10398
rect 8530 10334 8542 10386
rect 8594 10334 8606 10386
rect 8206 10322 8258 10334
rect 11566 10322 11618 10334
rect 11902 10386 11954 10398
rect 11902 10322 11954 10334
rect 41470 10386 41522 10398
rect 41470 10322 41522 10334
rect 41694 10386 41746 10398
rect 41694 10322 41746 10334
rect 46510 10386 46562 10398
rect 46510 10322 46562 10334
rect 46846 10386 46898 10398
rect 46846 10322 46898 10334
rect 1344 10218 49616 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 49616 10218
rect 1344 10132 49616 10166
rect 20302 10050 20354 10062
rect 11890 9998 11902 10050
rect 11954 9998 11966 10050
rect 20302 9986 20354 9998
rect 25790 10050 25842 10062
rect 25790 9986 25842 9998
rect 26462 10050 26514 10062
rect 45378 9998 45390 10050
rect 45442 9998 45454 10050
rect 26462 9986 26514 9998
rect 5854 9938 5906 9950
rect 12462 9938 12514 9950
rect 9426 9886 9438 9938
rect 9490 9886 9502 9938
rect 11554 9886 11566 9938
rect 11618 9886 11630 9938
rect 5854 9874 5906 9886
rect 12462 9874 12514 9886
rect 15262 9938 15314 9950
rect 20078 9938 20130 9950
rect 25678 9938 25730 9950
rect 19730 9886 19742 9938
rect 19794 9886 19806 9938
rect 21746 9886 21758 9938
rect 21810 9886 21822 9938
rect 15262 9874 15314 9886
rect 20078 9874 20130 9886
rect 25678 9874 25730 9886
rect 26686 9938 26738 9950
rect 37550 9938 37602 9950
rect 44830 9938 44882 9950
rect 35634 9886 35646 9938
rect 35698 9886 35710 9938
rect 41122 9886 41134 9938
rect 41186 9886 41198 9938
rect 47058 9886 47070 9938
rect 47122 9886 47134 9938
rect 49186 9886 49198 9938
rect 49250 9886 49262 9938
rect 26686 9874 26738 9886
rect 37550 9874 37602 9886
rect 44830 9874 44882 9886
rect 4734 9826 4786 9838
rect 4734 9762 4786 9774
rect 7310 9826 7362 9838
rect 7310 9762 7362 9774
rect 7758 9826 7810 9838
rect 7758 9762 7810 9774
rect 7870 9826 7922 9838
rect 7870 9762 7922 9774
rect 8318 9826 8370 9838
rect 12238 9826 12290 9838
rect 8754 9774 8766 9826
rect 8818 9774 8830 9826
rect 8318 9762 8370 9774
rect 12238 9762 12290 9774
rect 12910 9826 12962 9838
rect 15598 9826 15650 9838
rect 13682 9774 13694 9826
rect 13746 9774 13758 9826
rect 12910 9762 12962 9774
rect 15598 9762 15650 9774
rect 15710 9826 15762 9838
rect 15710 9762 15762 9774
rect 15822 9826 15874 9838
rect 21982 9826 22034 9838
rect 16818 9774 16830 9826
rect 16882 9774 16894 9826
rect 21634 9774 21646 9826
rect 21698 9774 21710 9826
rect 15822 9762 15874 9774
rect 21982 9762 22034 9774
rect 22878 9826 22930 9838
rect 22878 9762 22930 9774
rect 23550 9826 23602 9838
rect 23550 9762 23602 9774
rect 23774 9826 23826 9838
rect 23774 9762 23826 9774
rect 27134 9826 27186 9838
rect 27134 9762 27186 9774
rect 27806 9826 27858 9838
rect 36430 9826 36482 9838
rect 45054 9826 45106 9838
rect 28130 9774 28142 9826
rect 28194 9774 28206 9826
rect 29362 9774 29374 9826
rect 29426 9774 29438 9826
rect 30930 9774 30942 9826
rect 30994 9774 31006 9826
rect 31266 9774 31278 9826
rect 31330 9774 31342 9826
rect 32834 9774 32846 9826
rect 32898 9774 32910 9826
rect 37090 9774 37102 9826
rect 37154 9774 37166 9826
rect 38210 9774 38222 9826
rect 38274 9774 38286 9826
rect 41458 9774 41470 9826
rect 41522 9774 41534 9826
rect 46274 9774 46286 9826
rect 46338 9774 46350 9826
rect 27806 9762 27858 9774
rect 36430 9762 36482 9774
rect 45054 9762 45106 9774
rect 5182 9714 5234 9726
rect 22766 9714 22818 9726
rect 24446 9714 24498 9726
rect 17602 9662 17614 9714
rect 17666 9662 17678 9714
rect 23202 9662 23214 9714
rect 23266 9662 23278 9714
rect 5182 9650 5234 9662
rect 22766 9650 22818 9662
rect 24446 9650 24498 9662
rect 25566 9714 25618 9726
rect 27470 9714 27522 9726
rect 26114 9662 26126 9714
rect 26178 9662 26190 9714
rect 25566 9650 25618 9662
rect 27470 9650 27522 9662
rect 28590 9714 28642 9726
rect 29586 9662 29598 9714
rect 29650 9662 29662 9714
rect 33506 9662 33518 9714
rect 33570 9662 33582 9714
rect 36082 9662 36094 9714
rect 36146 9662 36158 9714
rect 38994 9662 39006 9714
rect 39058 9662 39070 9714
rect 28590 9650 28642 9662
rect 6302 9602 6354 9614
rect 6302 9538 6354 9550
rect 6638 9602 6690 9614
rect 6638 9538 6690 9550
rect 7086 9602 7138 9614
rect 7086 9538 7138 9550
rect 7198 9602 7250 9614
rect 7198 9538 7250 9550
rect 7646 9602 7698 9614
rect 14814 9602 14866 9614
rect 22430 9602 22482 9614
rect 13906 9550 13918 9602
rect 13970 9550 13982 9602
rect 16258 9550 16270 9602
rect 16322 9550 16334 9602
rect 20626 9550 20638 9602
rect 20690 9550 20702 9602
rect 7646 9538 7698 9550
rect 14814 9538 14866 9550
rect 22430 9538 22482 9550
rect 22654 9602 22706 9614
rect 22654 9538 22706 9550
rect 24222 9602 24274 9614
rect 24222 9538 24274 9550
rect 24334 9602 24386 9614
rect 24334 9538 24386 9550
rect 24782 9602 24834 9614
rect 42478 9602 42530 9614
rect 30258 9550 30270 9602
rect 30322 9550 30334 9602
rect 24782 9538 24834 9550
rect 42478 9538 42530 9550
rect 45838 9602 45890 9614
rect 45838 9538 45890 9550
rect 1344 9434 49616 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 49616 9434
rect 1344 9348 49616 9382
rect 8542 9266 8594 9278
rect 8542 9202 8594 9214
rect 8990 9266 9042 9278
rect 8990 9202 9042 9214
rect 9998 9266 10050 9278
rect 9998 9202 10050 9214
rect 10782 9266 10834 9278
rect 10782 9202 10834 9214
rect 11566 9266 11618 9278
rect 11566 9202 11618 9214
rect 11678 9266 11730 9278
rect 11678 9202 11730 9214
rect 12238 9266 12290 9278
rect 12238 9202 12290 9214
rect 14478 9266 14530 9278
rect 14478 9202 14530 9214
rect 16046 9266 16098 9278
rect 16046 9202 16098 9214
rect 18286 9266 18338 9278
rect 18286 9202 18338 9214
rect 18846 9266 18898 9278
rect 18846 9202 18898 9214
rect 19070 9266 19122 9278
rect 19070 9202 19122 9214
rect 22318 9266 22370 9278
rect 22318 9202 22370 9214
rect 23326 9266 23378 9278
rect 23326 9202 23378 9214
rect 25342 9266 25394 9278
rect 25342 9202 25394 9214
rect 25566 9266 25618 9278
rect 25566 9202 25618 9214
rect 27134 9266 27186 9278
rect 27134 9202 27186 9214
rect 28366 9266 28418 9278
rect 28366 9202 28418 9214
rect 31502 9266 31554 9278
rect 31502 9202 31554 9214
rect 39342 9266 39394 9278
rect 39342 9202 39394 9214
rect 40462 9266 40514 9278
rect 40462 9202 40514 9214
rect 41246 9266 41298 9278
rect 41246 9202 41298 9214
rect 41806 9266 41858 9278
rect 41806 9202 41858 9214
rect 42030 9266 42082 9278
rect 42030 9202 42082 9214
rect 46734 9266 46786 9278
rect 46734 9202 46786 9214
rect 47742 9266 47794 9278
rect 47742 9202 47794 9214
rect 13694 9154 13746 9166
rect 5954 9102 5966 9154
rect 6018 9102 6030 9154
rect 12898 9102 12910 9154
rect 12962 9102 12974 9154
rect 13694 9090 13746 9102
rect 15262 9154 15314 9166
rect 15262 9090 15314 9102
rect 16382 9154 16434 9166
rect 16382 9090 16434 9102
rect 16718 9154 16770 9166
rect 16718 9090 16770 9102
rect 20638 9154 20690 9166
rect 25902 9154 25954 9166
rect 21410 9102 21422 9154
rect 21474 9102 21486 9154
rect 20638 9090 20690 9102
rect 25902 9090 25954 9102
rect 30158 9154 30210 9166
rect 32510 9154 32562 9166
rect 31042 9102 31054 9154
rect 31106 9102 31118 9154
rect 30158 9090 30210 9102
rect 32510 9090 32562 9102
rect 33854 9154 33906 9166
rect 33854 9090 33906 9102
rect 33966 9154 34018 9166
rect 39566 9154 39618 9166
rect 36642 9102 36654 9154
rect 36706 9102 36718 9154
rect 45042 9102 45054 9154
rect 45106 9102 45118 9154
rect 48738 9102 48750 9154
rect 48802 9102 48814 9154
rect 33966 9090 34018 9102
rect 39566 9090 39618 9102
rect 11006 9042 11058 9054
rect 5282 8990 5294 9042
rect 5346 8990 5358 9042
rect 11006 8978 11058 8990
rect 11454 9042 11506 9054
rect 13582 9042 13634 9054
rect 13122 8990 13134 9042
rect 13186 8990 13198 9042
rect 11454 8978 11506 8990
rect 13582 8978 13634 8990
rect 13918 9042 13970 9054
rect 13918 8978 13970 8990
rect 15598 9042 15650 9054
rect 15598 8978 15650 8990
rect 19518 9042 19570 9054
rect 19518 8978 19570 8990
rect 20526 9042 20578 9054
rect 22878 9042 22930 9054
rect 21634 8990 21646 9042
rect 21698 8990 21710 9042
rect 20526 8978 20578 8990
rect 22878 8978 22930 8990
rect 23550 9042 23602 9054
rect 23550 8978 23602 8990
rect 23774 9042 23826 9054
rect 24446 9042 24498 9054
rect 24098 8990 24110 9042
rect 24162 8990 24174 9042
rect 23774 8978 23826 8990
rect 24446 8978 24498 8990
rect 24558 9042 24610 9054
rect 24558 8978 24610 8990
rect 24670 9042 24722 9054
rect 24670 8978 24722 8990
rect 25230 9042 25282 9054
rect 25230 8978 25282 8990
rect 25790 9042 25842 9054
rect 25790 8978 25842 8990
rect 28926 9042 28978 9054
rect 30046 9042 30098 9054
rect 29810 8990 29822 9042
rect 29874 8990 29886 9042
rect 28926 8978 28978 8990
rect 30046 8978 30098 8990
rect 30718 9042 30770 9054
rect 30718 8978 30770 8990
rect 31614 9042 31666 9054
rect 31614 8978 31666 8990
rect 32174 9042 32226 9054
rect 38334 9042 38386 9054
rect 34178 8990 34190 9042
rect 34242 8990 34254 9042
rect 37426 8990 37438 9042
rect 37490 8990 37502 9042
rect 37874 8990 37886 9042
rect 37938 8990 37950 9042
rect 32174 8978 32226 8990
rect 38334 8978 38386 8990
rect 38782 9042 38834 9054
rect 38782 8978 38834 8990
rect 39230 9042 39282 9054
rect 39230 8978 39282 8990
rect 39678 9042 39730 9054
rect 39678 8978 39730 8990
rect 41358 9042 41410 9054
rect 46622 9042 46674 9054
rect 45826 8990 45838 9042
rect 45890 8990 45902 9042
rect 46386 8990 46398 9042
rect 46450 8990 46462 9042
rect 41358 8978 41410 8990
rect 46622 8978 46674 8990
rect 46846 9042 46898 9054
rect 47630 9042 47682 9054
rect 47058 8990 47070 9042
rect 47122 8990 47134 9042
rect 47394 8990 47406 9042
rect 47458 8990 47470 9042
rect 46846 8978 46898 8990
rect 47630 8978 47682 8990
rect 47854 9042 47906 9054
rect 49086 9042 49138 9054
rect 48066 8990 48078 9042
rect 48130 8990 48142 9042
rect 47854 8978 47906 8990
rect 49086 8978 49138 8990
rect 10446 8930 10498 8942
rect 12574 8930 12626 8942
rect 8082 8878 8094 8930
rect 8146 8878 8158 8930
rect 10994 8878 11006 8930
rect 11058 8878 11070 8930
rect 10446 8866 10498 8878
rect 10210 8766 10222 8818
rect 10274 8815 10286 8818
rect 11009 8815 11055 8878
rect 12574 8866 12626 8878
rect 15038 8930 15090 8942
rect 15038 8866 15090 8878
rect 17502 8930 17554 8942
rect 18958 8930 19010 8942
rect 18162 8878 18174 8930
rect 18226 8878 18238 8930
rect 17502 8866 17554 8878
rect 18958 8866 19010 8878
rect 20078 8930 20130 8942
rect 20078 8866 20130 8878
rect 23662 8930 23714 8942
rect 23662 8866 23714 8878
rect 26462 8930 26514 8942
rect 28702 8930 28754 8942
rect 41918 8930 41970 8942
rect 27906 8878 27918 8930
rect 27970 8878 27982 8930
rect 34514 8878 34526 8930
rect 34578 8878 34590 8930
rect 26462 8866 26514 8878
rect 28702 8866 28754 8878
rect 41918 8866 41970 8878
rect 42590 8930 42642 8942
rect 42914 8878 42926 8930
rect 42978 8878 42990 8930
rect 42590 8866 42642 8878
rect 17390 8818 17442 8830
rect 10274 8769 11055 8815
rect 10274 8766 10286 8769
rect 11890 8766 11902 8818
rect 11954 8815 11966 8818
rect 12562 8815 12574 8818
rect 11954 8769 12574 8815
rect 11954 8766 11966 8769
rect 12562 8766 12574 8769
rect 12626 8766 12638 8818
rect 17390 8754 17442 8766
rect 18510 8818 18562 8830
rect 18510 8754 18562 8766
rect 20190 8818 20242 8830
rect 20190 8754 20242 8766
rect 20638 8818 20690 8830
rect 20638 8754 20690 8766
rect 25902 8818 25954 8830
rect 25902 8754 25954 8766
rect 26350 8818 26402 8830
rect 26350 8754 26402 8766
rect 29150 8818 29202 8830
rect 29150 8754 29202 8766
rect 29598 8818 29650 8830
rect 29598 8754 29650 8766
rect 31502 8818 31554 8830
rect 31502 8754 31554 8766
rect 32062 8818 32114 8830
rect 32062 8754 32114 8766
rect 32398 8818 32450 8830
rect 33394 8766 33406 8818
rect 33458 8766 33470 8818
rect 42354 8766 42366 8818
rect 42418 8815 42430 8818
rect 42690 8815 42702 8818
rect 42418 8769 42702 8815
rect 42418 8766 42430 8769
rect 42690 8766 42702 8769
rect 42754 8766 42766 8818
rect 32398 8754 32450 8766
rect 1344 8650 49616 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 49616 8650
rect 1344 8564 49616 8598
rect 36990 8482 37042 8494
rect 36990 8418 37042 8430
rect 8654 8370 8706 8382
rect 11342 8370 11394 8382
rect 20750 8370 20802 8382
rect 9538 8318 9550 8370
rect 9602 8318 9614 8370
rect 11666 8318 11678 8370
rect 11730 8318 11742 8370
rect 13906 8318 13918 8370
rect 13970 8318 13982 8370
rect 15474 8318 15486 8370
rect 15538 8318 15550 8370
rect 16930 8318 16942 8370
rect 16994 8318 17006 8370
rect 19058 8318 19070 8370
rect 19122 8318 19134 8370
rect 24098 8318 24110 8370
rect 24162 8318 24174 8370
rect 26226 8318 26238 8370
rect 26290 8318 26302 8370
rect 44258 8318 44270 8370
rect 44322 8318 44334 8370
rect 47058 8318 47070 8370
rect 47122 8318 47134 8370
rect 49186 8318 49198 8370
rect 49250 8318 49262 8370
rect 8654 8306 8706 8318
rect 11342 8306 11394 8318
rect 20750 8306 20802 8318
rect 7198 8258 7250 8270
rect 7198 8194 7250 8206
rect 7646 8258 7698 8270
rect 7646 8194 7698 8206
rect 7758 8258 7810 8270
rect 7758 8194 7810 8206
rect 8206 8258 8258 8270
rect 8206 8194 8258 8206
rect 8430 8258 8482 8270
rect 10782 8258 10834 8270
rect 10210 8206 10222 8258
rect 10274 8206 10286 8258
rect 8430 8194 8482 8206
rect 10782 8194 10834 8206
rect 11118 8258 11170 8270
rect 11118 8194 11170 8206
rect 12014 8258 12066 8270
rect 12014 8194 12066 8206
rect 12350 8258 12402 8270
rect 19406 8258 19458 8270
rect 21422 8258 21474 8270
rect 23102 8258 23154 8270
rect 28366 8258 28418 8270
rect 12674 8206 12686 8258
rect 12738 8206 12750 8258
rect 14130 8206 14142 8258
rect 14194 8206 14206 8258
rect 16146 8206 16158 8258
rect 16210 8206 16222 8258
rect 19842 8206 19854 8258
rect 19906 8206 19918 8258
rect 21746 8206 21758 8258
rect 21810 8206 21822 8258
rect 23426 8206 23438 8258
rect 23490 8206 23502 8258
rect 26786 8206 26798 8258
rect 26850 8206 26862 8258
rect 12350 8194 12402 8206
rect 19406 8194 19458 8206
rect 21422 8194 21474 8206
rect 23102 8194 23154 8206
rect 28366 8194 28418 8206
rect 28590 8258 28642 8270
rect 30942 8258 30994 8270
rect 33742 8258 33794 8270
rect 35870 8258 35922 8270
rect 29138 8206 29150 8258
rect 29202 8206 29214 8258
rect 32386 8206 32398 8258
rect 32450 8206 32462 8258
rect 34514 8206 34526 8258
rect 34578 8206 34590 8258
rect 28590 8194 28642 8206
rect 30942 8194 30994 8206
rect 33742 8194 33794 8206
rect 35870 8194 35922 8206
rect 37102 8258 37154 8270
rect 37102 8194 37154 8206
rect 37550 8258 37602 8270
rect 37550 8194 37602 8206
rect 37774 8258 37826 8270
rect 45502 8258 45554 8270
rect 38770 8206 38782 8258
rect 38834 8206 38846 8258
rect 41346 8206 41358 8258
rect 41410 8206 41422 8258
rect 45938 8206 45950 8258
rect 46002 8206 46014 8258
rect 46274 8206 46286 8258
rect 46338 8206 46350 8258
rect 37774 8194 37826 8206
rect 45502 8194 45554 8206
rect 6974 8146 7026 8158
rect 6974 8082 7026 8094
rect 9886 8146 9938 8158
rect 9886 8082 9938 8094
rect 10670 8146 10722 8158
rect 10670 8082 10722 8094
rect 12238 8146 12290 8158
rect 12238 8082 12290 8094
rect 13022 8146 13074 8158
rect 13022 8082 13074 8094
rect 14814 8146 14866 8158
rect 14814 8082 14866 8094
rect 15150 8146 15202 8158
rect 15150 8082 15202 8094
rect 20526 8146 20578 8158
rect 20526 8082 20578 8094
rect 21310 8146 21362 8158
rect 21310 8082 21362 8094
rect 22766 8146 22818 8158
rect 27694 8146 27746 8158
rect 26562 8094 26574 8146
rect 26626 8094 26638 8146
rect 22766 8082 22818 8094
rect 27694 8082 27746 8094
rect 28142 8146 28194 8158
rect 28142 8082 28194 8094
rect 30158 8146 30210 8158
rect 30158 8082 30210 8094
rect 33070 8146 33122 8158
rect 33070 8082 33122 8094
rect 33182 8146 33234 8158
rect 33182 8082 33234 8094
rect 34078 8146 34130 8158
rect 36318 8146 36370 8158
rect 45278 8146 45330 8158
rect 35074 8094 35086 8146
rect 35138 8094 35150 8146
rect 42130 8094 42142 8146
rect 42194 8094 42206 8146
rect 34078 8082 34130 8094
rect 36318 8082 36370 8094
rect 45278 8082 45330 8094
rect 5070 8034 5122 8046
rect 5070 7970 5122 7982
rect 6078 8034 6130 8046
rect 6078 7970 6130 7982
rect 6638 8034 6690 8046
rect 6638 7970 6690 7982
rect 7086 8034 7138 8046
rect 7086 7970 7138 7982
rect 7534 8034 7586 8046
rect 9662 8034 9714 8046
rect 8978 7982 8990 8034
rect 9042 7982 9054 8034
rect 7534 7970 7586 7982
rect 9662 7970 9714 7982
rect 10558 8034 10610 8046
rect 10558 7970 10610 7982
rect 15374 8034 15426 8046
rect 15374 7970 15426 7982
rect 20638 8034 20690 8046
rect 20638 7970 20690 7982
rect 22878 8034 22930 8046
rect 22878 7970 22930 7982
rect 27582 8034 27634 8046
rect 27582 7970 27634 7982
rect 28478 8034 28530 8046
rect 28478 7970 28530 7982
rect 29262 8034 29314 8046
rect 32846 8034 32898 8046
rect 32610 7982 32622 8034
rect 32674 7982 32686 8034
rect 29262 7970 29314 7982
rect 32846 7970 32898 7982
rect 33966 8034 34018 8046
rect 35422 8034 35474 8046
rect 34738 7982 34750 8034
rect 34802 7982 34814 8034
rect 33966 7970 34018 7982
rect 35422 7970 35474 7982
rect 35982 8034 36034 8046
rect 35982 7970 36034 7982
rect 36094 8034 36146 8046
rect 36094 7970 36146 7982
rect 36206 8034 36258 8046
rect 36206 7970 36258 7982
rect 37886 8034 37938 8046
rect 37886 7970 37938 7982
rect 39454 8034 39506 8046
rect 39454 7970 39506 7982
rect 44942 8034 44994 8046
rect 44942 7970 44994 7982
rect 45614 8034 45666 8046
rect 45614 7970 45666 7982
rect 45726 8034 45778 8046
rect 45726 7970 45778 7982
rect 1344 7866 49616 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 49616 7866
rect 1344 7780 49616 7814
rect 13022 7698 13074 7710
rect 13022 7634 13074 7646
rect 13246 7698 13298 7710
rect 13246 7634 13298 7646
rect 24334 7698 24386 7710
rect 24334 7634 24386 7646
rect 24446 7698 24498 7710
rect 24446 7634 24498 7646
rect 30270 7698 30322 7710
rect 30270 7634 30322 7646
rect 32286 7698 32338 7710
rect 32286 7634 32338 7646
rect 38894 7698 38946 7710
rect 42366 7698 42418 7710
rect 39554 7646 39566 7698
rect 39618 7646 39630 7698
rect 38894 7634 38946 7646
rect 42366 7634 42418 7646
rect 42478 7698 42530 7710
rect 42478 7634 42530 7646
rect 48862 7698 48914 7710
rect 48862 7634 48914 7646
rect 7758 7586 7810 7598
rect 5282 7534 5294 7586
rect 5346 7534 5358 7586
rect 7758 7522 7810 7534
rect 13470 7586 13522 7598
rect 23214 7586 23266 7598
rect 16034 7534 16046 7586
rect 16098 7534 16110 7586
rect 13470 7522 13522 7534
rect 23214 7522 23266 7534
rect 23326 7586 23378 7598
rect 23326 7522 23378 7534
rect 25230 7586 25282 7598
rect 25230 7522 25282 7534
rect 30046 7586 30098 7598
rect 30046 7522 30098 7534
rect 30494 7586 30546 7598
rect 30494 7522 30546 7534
rect 32510 7586 32562 7598
rect 32510 7522 32562 7534
rect 33182 7586 33234 7598
rect 33182 7522 33234 7534
rect 33630 7586 33682 7598
rect 33630 7522 33682 7534
rect 34078 7586 34130 7598
rect 40014 7586 40066 7598
rect 34962 7534 34974 7586
rect 35026 7534 35038 7586
rect 38546 7534 38558 7586
rect 38610 7534 38622 7586
rect 34078 7522 34130 7534
rect 40014 7522 40066 7534
rect 40910 7586 40962 7598
rect 40910 7522 40962 7534
rect 48974 7586 49026 7598
rect 48974 7522 49026 7534
rect 7982 7474 8034 7486
rect 8990 7474 9042 7486
rect 22990 7474 23042 7486
rect 4610 7422 4622 7474
rect 4674 7422 4686 7474
rect 8306 7422 8318 7474
rect 8370 7422 8382 7474
rect 9762 7422 9774 7474
rect 9826 7422 9838 7474
rect 16818 7422 16830 7474
rect 16882 7422 16894 7474
rect 22642 7422 22654 7474
rect 22706 7422 22718 7474
rect 7982 7410 8034 7422
rect 8990 7410 9042 7422
rect 22990 7410 23042 7422
rect 23774 7474 23826 7486
rect 23774 7410 23826 7422
rect 25342 7474 25394 7486
rect 25342 7410 25394 7422
rect 25566 7474 25618 7486
rect 27806 7474 27858 7486
rect 27570 7422 27582 7474
rect 27634 7422 27646 7474
rect 25566 7410 25618 7422
rect 27806 7410 27858 7422
rect 28030 7474 28082 7486
rect 30606 7474 30658 7486
rect 28466 7422 28478 7474
rect 28530 7422 28542 7474
rect 28030 7410 28082 7422
rect 30606 7410 30658 7422
rect 31054 7474 31106 7486
rect 31054 7410 31106 7422
rect 31614 7474 31666 7486
rect 31614 7410 31666 7422
rect 32958 7474 33010 7486
rect 32958 7410 33010 7422
rect 33294 7474 33346 7486
rect 41582 7474 41634 7486
rect 42590 7474 42642 7486
rect 34738 7422 34750 7474
rect 34802 7422 34814 7474
rect 38210 7422 38222 7474
rect 38274 7422 38286 7474
rect 39218 7422 39230 7474
rect 39282 7422 39294 7474
rect 39778 7422 39790 7474
rect 39842 7422 39854 7474
rect 41234 7422 41246 7474
rect 41298 7422 41310 7474
rect 42018 7422 42030 7474
rect 42082 7422 42094 7474
rect 43026 7422 43038 7474
rect 43090 7422 43102 7474
rect 33294 7410 33346 7422
rect 41582 7410 41634 7422
rect 42590 7410 42642 7422
rect 7870 7362 7922 7374
rect 13134 7362 13186 7374
rect 25678 7362 25730 7374
rect 39566 7362 39618 7374
rect 41694 7362 41746 7374
rect 7410 7310 7422 7362
rect 7474 7310 7486 7362
rect 10546 7310 10558 7362
rect 10610 7310 10622 7362
rect 12674 7310 12686 7362
rect 12738 7310 12750 7362
rect 13906 7310 13918 7362
rect 13970 7310 13982 7362
rect 17714 7310 17726 7362
rect 17778 7310 17790 7362
rect 30482 7310 30494 7362
rect 30546 7310 30558 7362
rect 33954 7310 33966 7362
rect 34018 7310 34030 7362
rect 35298 7310 35310 7362
rect 35362 7310 35374 7362
rect 37426 7310 37438 7362
rect 37490 7310 37502 7362
rect 41122 7310 41134 7362
rect 41186 7310 41198 7362
rect 45714 7310 45726 7362
rect 45778 7310 45790 7362
rect 7870 7298 7922 7310
rect 13134 7298 13186 7310
rect 25678 7298 25730 7310
rect 39566 7298 39618 7310
rect 41694 7298 41746 7310
rect 23998 7250 24050 7262
rect 23998 7186 24050 7198
rect 24558 7250 24610 7262
rect 32174 7250 32226 7262
rect 26450 7198 26462 7250
rect 26514 7198 26526 7250
rect 24558 7186 24610 7198
rect 32174 7186 32226 7198
rect 34302 7250 34354 7262
rect 34302 7186 34354 7198
rect 48750 7250 48802 7262
rect 48750 7186 48802 7198
rect 1344 7082 49616 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 49616 7082
rect 1344 6996 49616 7030
rect 7086 6914 7138 6926
rect 7086 6850 7138 6862
rect 7422 6914 7474 6926
rect 7422 6850 7474 6862
rect 8094 6914 8146 6926
rect 8094 6850 8146 6862
rect 30606 6914 30658 6926
rect 30606 6850 30658 6862
rect 30830 6914 30882 6926
rect 30830 6850 30882 6862
rect 34750 6914 34802 6926
rect 34750 6850 34802 6862
rect 5966 6802 6018 6814
rect 5966 6738 6018 6750
rect 8318 6802 8370 6814
rect 12014 6802 12066 6814
rect 30046 6802 30098 6814
rect 9538 6750 9550 6802
rect 9602 6750 9614 6802
rect 11666 6750 11678 6802
rect 11730 6750 11742 6802
rect 17378 6750 17390 6802
rect 17442 6750 17454 6802
rect 20626 6750 20638 6802
rect 20690 6750 20702 6802
rect 22642 6750 22654 6802
rect 22706 6799 22718 6802
rect 23314 6799 23326 6802
rect 22706 6753 23326 6799
rect 22706 6750 22718 6753
rect 23314 6750 23326 6753
rect 23378 6750 23390 6802
rect 25442 6750 25454 6802
rect 25506 6750 25518 6802
rect 32050 6750 32062 6802
rect 32114 6750 32126 6802
rect 34178 6750 34190 6802
rect 34242 6750 34254 6802
rect 35746 6750 35758 6802
rect 35810 6750 35822 6802
rect 37650 6750 37662 6802
rect 37714 6750 37726 6802
rect 39442 6750 39454 6802
rect 39506 6750 39518 6802
rect 41570 6750 41582 6802
rect 41634 6750 41646 6802
rect 42466 6750 42478 6802
rect 42530 6750 42542 6802
rect 43250 6750 43262 6802
rect 43314 6750 43326 6802
rect 45378 6750 45390 6802
rect 45442 6750 45454 6802
rect 49186 6750 49198 6802
rect 49250 6750 49262 6802
rect 8318 6738 8370 6750
rect 12014 6738 12066 6750
rect 30046 6738 30098 6750
rect 5182 6690 5234 6702
rect 5182 6626 5234 6638
rect 6302 6690 6354 6702
rect 6302 6626 6354 6638
rect 6750 6690 6802 6702
rect 12238 6690 12290 6702
rect 8866 6638 8878 6690
rect 8930 6638 8942 6690
rect 6750 6626 6802 6638
rect 12238 6626 12290 6638
rect 12350 6690 12402 6702
rect 13022 6690 13074 6702
rect 12674 6638 12686 6690
rect 12738 6638 12750 6690
rect 12350 6626 12402 6638
rect 13022 6626 13074 6638
rect 13358 6690 13410 6702
rect 13358 6626 13410 6638
rect 13582 6690 13634 6702
rect 13582 6626 13634 6638
rect 13694 6690 13746 6702
rect 13694 6626 13746 6638
rect 13918 6690 13970 6702
rect 29710 6690 29762 6702
rect 34526 6690 34578 6702
rect 36094 6690 36146 6702
rect 14578 6638 14590 6690
rect 14642 6638 14654 6690
rect 15250 6638 15262 6690
rect 15314 6638 15326 6690
rect 17714 6638 17726 6690
rect 17778 6638 17790 6690
rect 21410 6638 21422 6690
rect 21474 6638 21486 6690
rect 21858 6638 21870 6690
rect 21922 6638 21934 6690
rect 22418 6638 22430 6690
rect 22482 6638 22494 6690
rect 23314 6638 23326 6690
rect 23378 6638 23390 6690
rect 29474 6638 29486 6690
rect 29538 6638 29550 6690
rect 30370 6638 30382 6690
rect 30434 6638 30446 6690
rect 31266 6638 31278 6690
rect 31330 6638 31342 6690
rect 35074 6638 35086 6690
rect 35138 6638 35150 6690
rect 13918 6626 13970 6638
rect 29710 6626 29762 6638
rect 34526 6626 34578 6638
rect 36094 6626 36146 6638
rect 36990 6690 37042 6702
rect 37762 6638 37774 6690
rect 37826 6638 37838 6690
rect 38770 6638 38782 6690
rect 38834 6638 38846 6690
rect 41906 6638 41918 6690
rect 41970 6638 41982 6690
rect 42578 6638 42590 6690
rect 42642 6638 42654 6690
rect 43026 6638 43038 6690
rect 43090 6638 43102 6690
rect 46274 6638 46286 6690
rect 46338 6638 46350 6690
rect 47058 6638 47070 6690
rect 47122 6638 47134 6690
rect 36990 6626 37042 6638
rect 29038 6578 29090 6590
rect 36430 6578 36482 6590
rect 18498 6526 18510 6578
rect 18562 6526 18574 6578
rect 21746 6526 21758 6578
rect 21810 6526 21822 6578
rect 29922 6526 29934 6578
rect 29986 6526 29998 6578
rect 29038 6514 29090 6526
rect 36430 6514 36482 6526
rect 37102 6578 37154 6590
rect 37102 6514 37154 6526
rect 38334 6578 38386 6590
rect 38334 6514 38386 6526
rect 42142 6578 42194 6590
rect 43710 6578 43762 6590
rect 42690 6526 42702 6578
rect 42754 6575 42766 6578
rect 42914 6575 42926 6578
rect 42754 6529 42926 6575
rect 42754 6526 42766 6529
rect 42914 6526 42926 6529
rect 42978 6526 42990 6578
rect 42142 6514 42194 6526
rect 43710 6514 43762 6526
rect 44158 6578 44210 6590
rect 44158 6514 44210 6526
rect 45502 6578 45554 6590
rect 45502 6514 45554 6526
rect 45950 6578 46002 6590
rect 45950 6514 46002 6526
rect 4734 6466 4786 6478
rect 4734 6402 4786 6414
rect 7198 6466 7250 6478
rect 30494 6466 30546 6478
rect 7746 6414 7758 6466
rect 7810 6414 7822 6466
rect 7198 6402 7250 6414
rect 30494 6402 30546 6414
rect 42366 6466 42418 6478
rect 42366 6402 42418 6414
rect 43262 6466 43314 6478
rect 43262 6402 43314 6414
rect 43486 6466 43538 6478
rect 43486 6402 43538 6414
rect 44046 6466 44098 6478
rect 44046 6402 44098 6414
rect 44942 6466 44994 6478
rect 44942 6402 44994 6414
rect 45390 6466 45442 6478
rect 45390 6402 45442 6414
rect 45726 6466 45778 6478
rect 45726 6402 45778 6414
rect 1344 6298 49616 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 49616 6298
rect 1344 6212 49616 6246
rect 4734 6130 4786 6142
rect 4734 6066 4786 6078
rect 17726 6130 17778 6142
rect 17726 6066 17778 6078
rect 17838 6130 17890 6142
rect 39902 6130 39954 6142
rect 39106 6078 39118 6130
rect 39170 6078 39182 6130
rect 17838 6066 17890 6078
rect 39902 6066 39954 6078
rect 40014 6130 40066 6142
rect 40014 6066 40066 6078
rect 46734 6130 46786 6142
rect 46734 6066 46786 6078
rect 46846 6130 46898 6142
rect 46846 6066 46898 6078
rect 46958 6130 47010 6142
rect 47506 6078 47518 6130
rect 47570 6078 47582 6130
rect 48738 6078 48750 6130
rect 48802 6078 48814 6130
rect 46958 6066 47010 6078
rect 17950 6018 18002 6030
rect 24222 6018 24274 6030
rect 6178 5966 6190 6018
rect 6242 5966 6254 6018
rect 8978 5966 8990 6018
rect 9042 5966 9054 6018
rect 19618 5966 19630 6018
rect 19682 5966 19694 6018
rect 20738 5966 20750 6018
rect 20802 5966 20814 6018
rect 23538 5966 23550 6018
rect 23602 5966 23614 6018
rect 17950 5954 18002 5966
rect 24222 5954 24274 5966
rect 25454 6018 25506 6030
rect 25454 5954 25506 5966
rect 25790 6018 25842 6030
rect 25790 5954 25842 5966
rect 27134 6018 27186 6030
rect 39454 6018 39506 6030
rect 28578 5966 28590 6018
rect 28642 5966 28654 6018
rect 39218 5966 39230 6018
rect 39282 5966 39294 6018
rect 27134 5954 27186 5966
rect 39454 5954 39506 5966
rect 40126 6018 40178 6030
rect 40126 5954 40178 5966
rect 46510 6018 46562 6030
rect 46510 5954 46562 5966
rect 8654 5906 8706 5918
rect 25902 5906 25954 5918
rect 5506 5854 5518 5906
rect 5570 5854 5582 5906
rect 14354 5854 14366 5906
rect 14418 5854 14430 5906
rect 16146 5854 16158 5906
rect 16210 5854 16222 5906
rect 16930 5854 16942 5906
rect 16994 5854 17006 5906
rect 18610 5854 18622 5906
rect 18674 5854 18686 5906
rect 18946 5854 18958 5906
rect 19010 5854 19022 5906
rect 20066 5854 20078 5906
rect 20130 5854 20142 5906
rect 23650 5854 23662 5906
rect 23714 5854 23726 5906
rect 24434 5854 24446 5906
rect 24498 5854 24510 5906
rect 8654 5842 8706 5854
rect 25902 5842 25954 5854
rect 26910 5906 26962 5918
rect 39006 5906 39058 5918
rect 27794 5854 27806 5906
rect 27858 5854 27870 5906
rect 31826 5854 31838 5906
rect 31890 5854 31902 5906
rect 38322 5854 38334 5906
rect 38386 5854 38398 5906
rect 38658 5854 38670 5906
rect 38722 5854 38734 5906
rect 41234 5854 41246 5906
rect 41298 5854 41310 5906
rect 47170 5854 47182 5906
rect 47234 5854 47246 5906
rect 47730 5854 47742 5906
rect 47794 5854 47806 5906
rect 48962 5854 48974 5906
rect 49026 5854 49038 5906
rect 26910 5842 26962 5854
rect 39006 5842 39058 5854
rect 4286 5794 4338 5806
rect 4286 5730 4338 5742
rect 5182 5794 5234 5806
rect 25566 5794 25618 5806
rect 8306 5742 8318 5794
rect 8370 5742 8382 5794
rect 9986 5742 9998 5794
rect 10050 5742 10062 5794
rect 16258 5742 16270 5794
rect 16322 5742 16334 5794
rect 19058 5742 19070 5794
rect 19122 5742 19134 5794
rect 22866 5742 22878 5794
rect 22930 5742 22942 5794
rect 23202 5742 23214 5794
rect 23266 5742 23278 5794
rect 30706 5742 30718 5794
rect 30770 5742 30782 5794
rect 31938 5742 31950 5794
rect 32002 5742 32014 5794
rect 33730 5742 33742 5794
rect 33794 5742 33806 5794
rect 42914 5742 42926 5794
rect 42978 5742 42990 5794
rect 5182 5730 5234 5742
rect 25566 5730 25618 5742
rect 16718 5682 16770 5694
rect 4274 5630 4286 5682
rect 4338 5679 4350 5682
rect 5058 5679 5070 5682
rect 4338 5633 5070 5679
rect 4338 5630 4350 5633
rect 5058 5630 5070 5633
rect 5122 5630 5134 5682
rect 16718 5618 16770 5630
rect 26574 5682 26626 5694
rect 32386 5630 32398 5682
rect 32450 5630 32462 5682
rect 26574 5618 26626 5630
rect 1344 5514 49616 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 49616 5514
rect 1344 5428 49616 5462
rect 7198 5346 7250 5358
rect 7198 5282 7250 5294
rect 19070 5346 19122 5358
rect 19070 5282 19122 5294
rect 27470 5346 27522 5358
rect 27470 5282 27522 5294
rect 30382 5346 30434 5358
rect 30382 5282 30434 5294
rect 34078 5346 34130 5358
rect 34078 5282 34130 5294
rect 36430 5346 36482 5358
rect 36430 5282 36482 5294
rect 5182 5234 5234 5246
rect 5182 5170 5234 5182
rect 6078 5234 6130 5246
rect 6078 5170 6130 5182
rect 6526 5234 6578 5246
rect 18958 5234 19010 5246
rect 22318 5234 22370 5246
rect 12898 5182 12910 5234
rect 12962 5182 12974 5234
rect 15250 5182 15262 5234
rect 15314 5182 15326 5234
rect 15586 5182 15598 5234
rect 15650 5182 15662 5234
rect 20402 5182 20414 5234
rect 20466 5182 20478 5234
rect 24994 5182 25006 5234
rect 25058 5182 25070 5234
rect 27122 5182 27134 5234
rect 27186 5182 27198 5234
rect 30818 5182 30830 5234
rect 30882 5182 30894 5234
rect 35746 5182 35758 5234
rect 35810 5182 35822 5234
rect 36978 5182 36990 5234
rect 37042 5182 37054 5234
rect 39106 5182 39118 5234
rect 39170 5182 39182 5234
rect 43138 5182 43150 5234
rect 43202 5182 43214 5234
rect 46050 5182 46062 5234
rect 46114 5182 46126 5234
rect 48178 5182 48190 5234
rect 48242 5182 48254 5234
rect 48738 5182 48750 5234
rect 48802 5182 48814 5234
rect 6526 5170 6578 5182
rect 18958 5170 19010 5182
rect 22318 5170 22370 5182
rect 7422 5122 7474 5134
rect 7422 5058 7474 5070
rect 7982 5122 8034 5134
rect 7982 5058 8034 5070
rect 8430 5122 8482 5134
rect 8430 5058 8482 5070
rect 8766 5122 8818 5134
rect 8766 5058 8818 5070
rect 8990 5122 9042 5134
rect 13694 5122 13746 5134
rect 14590 5122 14642 5134
rect 9986 5070 9998 5122
rect 10050 5070 10062 5122
rect 13906 5070 13918 5122
rect 13970 5070 13982 5122
rect 8990 5058 9042 5070
rect 13694 5058 13746 5070
rect 14590 5058 14642 5070
rect 14926 5122 14978 5134
rect 27582 5122 27634 5134
rect 30494 5122 30546 5134
rect 34190 5122 34242 5134
rect 34750 5122 34802 5134
rect 35422 5122 35474 5134
rect 43598 5122 43650 5134
rect 18498 5070 18510 5122
rect 18562 5070 18574 5122
rect 19730 5070 19742 5122
rect 19794 5070 19806 5122
rect 20178 5070 20190 5122
rect 20242 5070 20254 5122
rect 21298 5070 21310 5122
rect 21362 5070 21374 5122
rect 24322 5070 24334 5122
rect 24386 5070 24398 5122
rect 29250 5070 29262 5122
rect 29314 5070 29326 5122
rect 32946 5070 32958 5122
rect 33010 5070 33022 5122
rect 33730 5070 33742 5122
rect 33794 5070 33806 5122
rect 34402 5070 34414 5122
rect 34466 5070 34478 5122
rect 35074 5070 35086 5122
rect 35138 5070 35150 5122
rect 36418 5070 36430 5122
rect 36482 5070 36494 5122
rect 39890 5070 39902 5122
rect 39954 5070 39966 5122
rect 40338 5070 40350 5122
rect 40402 5070 40414 5122
rect 14926 5058 14978 5070
rect 27582 5058 27634 5070
rect 30494 5058 30546 5070
rect 34190 5058 34242 5070
rect 34750 5058 34802 5070
rect 35422 5058 35474 5070
rect 43598 5058 43650 5070
rect 43710 5122 43762 5134
rect 43710 5058 43762 5070
rect 43822 5122 43874 5134
rect 43822 5058 43874 5070
rect 44046 5122 44098 5134
rect 49198 5122 49250 5134
rect 45266 5070 45278 5122
rect 45330 5070 45342 5122
rect 44046 5058 44098 5070
rect 49198 5058 49250 5070
rect 15150 5010 15202 5022
rect 27694 5010 27746 5022
rect 10770 4958 10782 5010
rect 10834 4958 10846 5010
rect 17714 4958 17726 5010
rect 17778 4958 17790 5010
rect 20738 4958 20750 5010
rect 20802 4958 20814 5010
rect 15150 4946 15202 4958
rect 27694 4946 27746 4958
rect 29598 5010 29650 5022
rect 29598 4946 29650 4958
rect 35646 5010 35698 5022
rect 35646 4946 35698 4958
rect 36094 5010 36146 5022
rect 41010 4958 41022 5010
rect 41074 4958 41086 5010
rect 36094 4946 36146 4958
rect 7758 4898 7810 4910
rect 6850 4846 6862 4898
rect 6914 4846 6926 4898
rect 7758 4834 7810 4846
rect 7870 4898 7922 4910
rect 7870 4834 7922 4846
rect 9438 4898 9490 4910
rect 9438 4834 9490 4846
rect 9550 4898 9602 4910
rect 9550 4834 9602 4846
rect 9662 4898 9714 4910
rect 9662 4834 9714 4846
rect 28142 4898 28194 4910
rect 28142 4834 28194 4846
rect 29710 4898 29762 4910
rect 29710 4834 29762 4846
rect 29822 4898 29874 4910
rect 29822 4834 29874 4846
rect 34862 4898 34914 4910
rect 34862 4834 34914 4846
rect 43934 4898 43986 4910
rect 43934 4834 43986 4846
rect 44830 4898 44882 4910
rect 44830 4834 44882 4846
rect 1344 4730 49616 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 49616 4730
rect 1344 4644 49616 4678
rect 4846 4562 4898 4574
rect 4846 4498 4898 4510
rect 8542 4562 8594 4574
rect 8542 4498 8594 4510
rect 12910 4562 12962 4574
rect 12910 4498 12962 4510
rect 13134 4562 13186 4574
rect 13134 4498 13186 4510
rect 20414 4562 20466 4574
rect 20414 4498 20466 4510
rect 24558 4562 24610 4574
rect 24558 4498 24610 4510
rect 32286 4562 32338 4574
rect 49086 4562 49138 4574
rect 33954 4510 33966 4562
rect 34018 4510 34030 4562
rect 48738 4510 48750 4562
rect 48802 4510 48814 4562
rect 32286 4498 32338 4510
rect 49086 4498 49138 4510
rect 24670 4450 24722 4462
rect 16034 4398 16046 4450
rect 16098 4398 16110 4450
rect 24670 4386 24722 4398
rect 25230 4450 25282 4462
rect 25230 4386 25282 4398
rect 25790 4450 25842 4462
rect 25790 4386 25842 4398
rect 26686 4450 26738 4462
rect 26686 4386 26738 4398
rect 26910 4450 26962 4462
rect 26910 4386 26962 4398
rect 27022 4450 27074 4462
rect 27022 4386 27074 4398
rect 30718 4450 30770 4462
rect 30718 4386 30770 4398
rect 31278 4450 31330 4462
rect 31278 4386 31330 4398
rect 31614 4450 31666 4462
rect 31614 4386 31666 4398
rect 32510 4450 32562 4462
rect 32510 4386 32562 4398
rect 33070 4450 33122 4462
rect 44158 4450 44210 4462
rect 35074 4398 35086 4450
rect 35138 4398 35150 4450
rect 41682 4398 41694 4450
rect 41746 4398 41758 4450
rect 33070 4386 33122 4398
rect 44158 4386 44210 4398
rect 44382 4450 44434 4462
rect 44382 4386 44434 4398
rect 48078 4450 48130 4462
rect 48078 4386 48130 4398
rect 25454 4338 25506 4350
rect 31054 4338 31106 4350
rect 5058 4286 5070 4338
rect 5122 4286 5134 4338
rect 9650 4286 9662 4338
rect 9714 4286 9726 4338
rect 13458 4286 13470 4338
rect 13522 4286 13534 4338
rect 16818 4286 16830 4338
rect 16882 4286 16894 4338
rect 17490 4286 17502 4338
rect 17554 4286 17566 4338
rect 24098 4286 24110 4338
rect 24162 4286 24174 4338
rect 26450 4286 26462 4338
rect 26514 4286 26526 4338
rect 27570 4286 27582 4338
rect 27634 4286 27646 4338
rect 33730 4286 33742 4338
rect 33794 4286 33806 4338
rect 34402 4286 34414 4338
rect 34466 4286 34478 4338
rect 37538 4286 37550 4338
rect 37602 4286 37614 4338
rect 40898 4286 40910 4338
rect 40962 4286 40974 4338
rect 44818 4286 44830 4338
rect 44882 4286 44894 4338
rect 25454 4274 25506 4286
rect 31054 4274 31106 4286
rect 8430 4226 8482 4238
rect 13022 4226 13074 4238
rect 20526 4226 20578 4238
rect 25342 4226 25394 4238
rect 5842 4174 5854 4226
rect 5906 4174 5918 4226
rect 7970 4174 7982 4226
rect 8034 4174 8046 4226
rect 10322 4174 10334 4226
rect 10386 4174 10398 4226
rect 12450 4174 12462 4226
rect 12514 4174 12526 4226
rect 13906 4174 13918 4226
rect 13970 4174 13982 4226
rect 21186 4174 21198 4226
rect 21250 4174 21262 4226
rect 23314 4174 23326 4226
rect 23378 4174 23390 4226
rect 8430 4162 8482 4174
rect 13022 4162 13074 4174
rect 20526 4162 20578 4174
rect 25342 4162 25394 4174
rect 26238 4226 26290 4238
rect 31166 4226 31218 4238
rect 44270 4226 44322 4238
rect 28242 4174 28254 4226
rect 28306 4174 28318 4226
rect 30370 4174 30382 4226
rect 30434 4174 30446 4226
rect 37202 4174 37214 4226
rect 37266 4174 37278 4226
rect 43810 4174 43822 4226
rect 43874 4174 43886 4226
rect 45602 4174 45614 4226
rect 45666 4174 45678 4226
rect 47730 4174 47742 4226
rect 47794 4174 47806 4226
rect 26238 4162 26290 4174
rect 31166 4162 31218 4174
rect 44270 4162 44322 4174
rect 8318 4114 8370 4126
rect 8318 4050 8370 4062
rect 18510 4114 18562 4126
rect 18510 4050 18562 4062
rect 24558 4114 24610 4126
rect 24558 4050 24610 4062
rect 26126 4114 26178 4126
rect 26126 4050 26178 4062
rect 32174 4114 32226 4126
rect 32174 4050 32226 4062
rect 38558 4114 38610 4126
rect 38558 4050 38610 4062
rect 1344 3946 49616 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 49616 3946
rect 1344 3860 49616 3894
rect 9550 3778 9602 3790
rect 9550 3714 9602 3726
rect 9886 3778 9938 3790
rect 9886 3714 9938 3726
rect 10446 3778 10498 3790
rect 11342 3778 11394 3790
rect 10770 3726 10782 3778
rect 10834 3726 10846 3778
rect 10446 3714 10498 3726
rect 11342 3714 11394 3726
rect 13246 3778 13298 3790
rect 13246 3714 13298 3726
rect 47406 3778 47458 3790
rect 47406 3714 47458 3726
rect 5070 3666 5122 3678
rect 5070 3602 5122 3614
rect 6526 3666 6578 3678
rect 6526 3602 6578 3614
rect 10222 3666 10274 3678
rect 10222 3602 10274 3614
rect 11230 3666 11282 3678
rect 11230 3602 11282 3614
rect 11790 3666 11842 3678
rect 40798 3666 40850 3678
rect 47518 3666 47570 3678
rect 20850 3614 20862 3666
rect 20914 3614 20926 3666
rect 22978 3614 22990 3666
rect 23042 3614 23054 3666
rect 25330 3614 25342 3666
rect 25394 3614 25406 3666
rect 27458 3614 27470 3666
rect 27522 3614 27534 3666
rect 30482 3614 30494 3666
rect 30546 3614 30558 3666
rect 32946 3614 32958 3666
rect 33010 3614 33022 3666
rect 35074 3614 35086 3666
rect 35138 3614 35150 3666
rect 36754 3614 36766 3666
rect 36818 3614 36830 3666
rect 38882 3614 38894 3666
rect 38946 3614 38958 3666
rect 44706 3614 44718 3666
rect 44770 3614 44782 3666
rect 46834 3614 46846 3666
rect 46898 3614 46910 3666
rect 48738 3614 48750 3666
rect 48802 3614 48814 3666
rect 11790 3602 11842 3614
rect 40798 3602 40850 3614
rect 47518 3602 47570 3614
rect 11678 3554 11730 3566
rect 11678 3490 11730 3502
rect 12014 3554 12066 3566
rect 12014 3490 12066 3502
rect 12238 3554 12290 3566
rect 49198 3554 49250 3566
rect 16370 3502 16382 3554
rect 16434 3502 16446 3554
rect 17042 3502 17054 3554
rect 17106 3502 17118 3554
rect 19730 3502 19742 3554
rect 19794 3502 19806 3554
rect 23762 3502 23774 3554
rect 23826 3502 23838 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 31378 3502 31390 3554
rect 31442 3502 31454 3554
rect 32274 3502 32286 3554
rect 32338 3502 32350 3554
rect 35970 3502 35982 3554
rect 36034 3502 36046 3554
rect 39778 3502 39790 3554
rect 39842 3502 39854 3554
rect 42802 3502 42814 3554
rect 42866 3502 42878 3554
rect 44034 3502 44046 3554
rect 44098 3502 44110 3554
rect 12238 3490 12290 3502
rect 49198 3490 49250 3502
rect 9774 3442 9826 3454
rect 13246 3442 13298 3454
rect 9774 3378 9826 3390
rect 13134 3386 13186 3398
rect 1710 3330 1762 3342
rect 1710 3266 1762 3278
rect 3166 3330 3218 3342
rect 3166 3266 3218 3278
rect 5518 3330 5570 3342
rect 5518 3266 5570 3278
rect 6750 3330 6802 3342
rect 6750 3266 6802 3278
rect 7422 3330 7474 3342
rect 7422 3266 7474 3278
rect 7870 3330 7922 3342
rect 7870 3266 7922 3278
rect 8318 3330 8370 3342
rect 8318 3266 8370 3278
rect 8766 3330 8818 3342
rect 13246 3378 13298 3390
rect 17278 3442 17330 3454
rect 47630 3442 47682 3454
rect 43026 3390 43038 3442
rect 43090 3390 43102 3442
rect 17278 3378 17330 3390
rect 47630 3378 47682 3390
rect 13134 3322 13186 3334
rect 15374 3330 15426 3342
rect 8766 3266 8818 3278
rect 15374 3266 15426 3278
rect 19182 3330 19234 3342
rect 19182 3266 19234 3278
rect 28366 3330 28418 3342
rect 28366 3266 28418 3278
rect 48078 3330 48130 3342
rect 48078 3266 48130 3278
rect 1344 3162 49616 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 49616 3162
rect 1344 3076 49616 3110
rect 7410 1710 7422 1762
rect 7474 1759 7486 1762
rect 8306 1759 8318 1762
rect 7474 1713 8318 1759
rect 7474 1710 7486 1713
rect 8306 1710 8318 1713
rect 8370 1710 8382 1762
<< via1 >>
rect 5518 47966 5570 48018
rect 6526 47966 6578 48018
rect 30830 47966 30882 48018
rect 31614 47966 31666 48018
rect 34078 47966 34130 48018
rect 35086 47966 35138 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 6526 47630 6578 47682
rect 42366 47630 42418 47682
rect 45390 47630 45442 47682
rect 19070 47518 19122 47570
rect 30830 47518 30882 47570
rect 35086 47518 35138 47570
rect 40574 47518 40626 47570
rect 44494 47518 44546 47570
rect 48750 47518 48802 47570
rect 19294 47406 19346 47458
rect 31614 47406 31666 47458
rect 32174 47406 32226 47458
rect 40014 47406 40066 47458
rect 41918 47406 41970 47458
rect 42142 47406 42194 47458
rect 42814 47406 42866 47458
rect 43710 47406 43762 47458
rect 44830 47406 44882 47458
rect 45614 47406 45666 47458
rect 45838 47406 45890 47458
rect 46398 47406 46450 47458
rect 47742 47406 47794 47458
rect 48190 47406 48242 47458
rect 49086 47406 49138 47458
rect 6862 47294 6914 47346
rect 19854 47294 19906 47346
rect 26574 47294 26626 47346
rect 29710 47294 29762 47346
rect 31054 47294 31106 47346
rect 32958 47294 33010 47346
rect 36318 47294 36370 47346
rect 38782 47294 38834 47346
rect 41582 47294 41634 47346
rect 45278 47294 45330 47346
rect 6638 47182 6690 47234
rect 26238 47182 26290 47234
rect 29374 47182 29426 47234
rect 35982 47182 36034 47234
rect 36878 47182 36930 47234
rect 37438 47182 37490 47234
rect 37774 47182 37826 47234
rect 38334 47182 38386 47234
rect 39230 47182 39282 47234
rect 41022 47182 41074 47234
rect 41358 47182 41410 47234
rect 41470 47182 41522 47234
rect 42030 47182 42082 47234
rect 42926 47182 42978 47234
rect 43934 47182 43986 47234
rect 46174 47182 46226 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 32398 46846 32450 46898
rect 33742 46846 33794 46898
rect 34190 46846 34242 46898
rect 5518 46734 5570 46786
rect 8430 46734 8482 46786
rect 26014 46734 26066 46786
rect 29598 46734 29650 46786
rect 35198 46734 35250 46786
rect 41694 46734 41746 46786
rect 45054 46734 45106 46786
rect 47518 46734 47570 46786
rect 48750 46734 48802 46786
rect 6302 46622 6354 46674
rect 7086 46622 7138 46674
rect 8094 46622 8146 46674
rect 21646 46622 21698 46674
rect 25230 46622 25282 46674
rect 28926 46622 28978 46674
rect 32062 46622 32114 46674
rect 34414 46622 34466 46674
rect 41022 46622 41074 46674
rect 44382 46622 44434 46674
rect 47854 46622 47906 46674
rect 48974 46622 49026 46674
rect 3390 46510 3442 46562
rect 6750 46510 6802 46562
rect 7310 46510 7362 46562
rect 8206 46510 8258 46562
rect 18846 46510 18898 46562
rect 20974 46510 21026 46562
rect 28142 46510 28194 46562
rect 31726 46510 31778 46562
rect 37326 46510 37378 46562
rect 37886 46510 37938 46562
rect 38334 46510 38386 46562
rect 38894 46510 38946 46562
rect 39342 46510 39394 46562
rect 39790 46510 39842 46562
rect 40462 46510 40514 46562
rect 43822 46510 43874 46562
rect 47182 46510 47234 46562
rect 37998 46398 38050 46450
rect 38446 46398 38498 46450
rect 38670 46398 38722 46450
rect 38894 46398 38946 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 27022 46062 27074 46114
rect 29710 46062 29762 46114
rect 30270 46062 30322 46114
rect 41246 46062 41298 46114
rect 44270 46062 44322 46114
rect 10558 45950 10610 46002
rect 31950 45950 32002 46002
rect 38446 45950 38498 46002
rect 40574 45950 40626 46002
rect 44158 45950 44210 46002
rect 46286 45950 46338 46002
rect 4510 45838 4562 45890
rect 4734 45838 4786 45890
rect 4958 45838 5010 45890
rect 5854 45838 5906 45890
rect 7086 45838 7138 45890
rect 7758 45838 7810 45890
rect 26574 45838 26626 45890
rect 27358 45838 27410 45890
rect 27582 45838 27634 45890
rect 29150 45838 29202 45890
rect 29374 45838 29426 45890
rect 30606 45838 30658 45890
rect 30830 45838 30882 45890
rect 36430 45838 36482 45890
rect 37326 45838 37378 45890
rect 37662 45838 37714 45890
rect 41582 45838 41634 45890
rect 41806 45838 41858 45890
rect 42702 45838 42754 45890
rect 43038 45838 43090 45890
rect 43934 45838 43986 45890
rect 45390 45838 45442 45890
rect 45726 45838 45778 45890
rect 45838 45838 45890 45890
rect 49086 45838 49138 45890
rect 4398 45726 4450 45778
rect 6750 45726 6802 45778
rect 7198 45726 7250 45778
rect 7310 45726 7362 45778
rect 8430 45726 8482 45778
rect 26686 45726 26738 45778
rect 27918 45726 27970 45778
rect 28030 45726 28082 45778
rect 28254 45726 28306 45778
rect 28478 45726 28530 45778
rect 36990 45726 37042 45778
rect 42590 45726 42642 45778
rect 44942 45726 44994 45778
rect 48414 45726 48466 45778
rect 6078 45614 6130 45666
rect 26462 45614 26514 45666
rect 37102 45614 37154 45666
rect 43262 45614 43314 45666
rect 43486 45614 43538 45666
rect 44830 45614 44882 45666
rect 45614 45614 45666 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 9662 45278 9714 45330
rect 28142 45278 28194 45330
rect 30046 45278 30098 45330
rect 30718 45278 30770 45330
rect 36430 45278 36482 45330
rect 41806 45278 41858 45330
rect 3054 45166 3106 45218
rect 8206 45166 8258 45218
rect 21646 45166 21698 45218
rect 25230 45166 25282 45218
rect 29934 45166 29986 45218
rect 31502 45166 31554 45218
rect 32958 45166 33010 45218
rect 35534 45166 35586 45218
rect 38110 45166 38162 45218
rect 41246 45166 41298 45218
rect 41694 45166 41746 45218
rect 42366 45166 42418 45218
rect 45278 45166 45330 45218
rect 48750 45166 48802 45218
rect 2270 45054 2322 45106
rect 8990 45054 9042 45106
rect 23550 45054 23602 45106
rect 25566 45054 25618 45106
rect 26910 45054 26962 45106
rect 27134 45054 27186 45106
rect 28590 45054 28642 45106
rect 28702 45054 28754 45106
rect 28814 45054 28866 45106
rect 30270 45054 30322 45106
rect 30606 45054 30658 45106
rect 30942 45054 30994 45106
rect 31166 45054 31218 45106
rect 32174 45054 32226 45106
rect 33406 45054 33458 45106
rect 33630 45054 33682 45106
rect 33742 45054 33794 45106
rect 33854 45054 33906 45106
rect 35086 45054 35138 45106
rect 36094 45054 36146 45106
rect 37438 45054 37490 45106
rect 47070 45054 47122 45106
rect 49086 45054 49138 45106
rect 5182 44942 5234 44994
rect 6078 44942 6130 44994
rect 9550 44942 9602 44994
rect 18734 44942 18786 44994
rect 27806 44942 27858 44994
rect 32398 44942 32450 44994
rect 35198 44942 35250 44994
rect 35870 44942 35922 44994
rect 37102 44942 37154 44994
rect 40238 44942 40290 44994
rect 41358 44942 41410 44994
rect 42478 44942 42530 44994
rect 9886 44830 9938 44882
rect 41806 44830 41858 44882
rect 42590 44830 42642 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 20414 44494 20466 44546
rect 27022 44494 27074 44546
rect 27358 44494 27410 44546
rect 48078 44494 48130 44546
rect 48414 44494 48466 44546
rect 48862 44494 48914 44546
rect 49310 44494 49362 44546
rect 4622 44382 4674 44434
rect 8990 44382 9042 44434
rect 19294 44382 19346 44434
rect 24558 44382 24610 44434
rect 26686 44382 26738 44434
rect 32062 44382 32114 44434
rect 32510 44382 32562 44434
rect 33406 44382 33458 44434
rect 34750 44382 34802 44434
rect 37214 44382 37266 44434
rect 38334 44382 38386 44434
rect 40462 44382 40514 44434
rect 41134 44382 41186 44434
rect 45614 44382 45666 44434
rect 47182 44382 47234 44434
rect 1822 44270 1874 44322
rect 5742 44270 5794 44322
rect 5854 44270 5906 44322
rect 6190 44270 6242 44322
rect 12238 44270 12290 44322
rect 16494 44270 16546 44322
rect 21982 44270 22034 44322
rect 23886 44270 23938 44322
rect 27582 44270 27634 44322
rect 27918 44270 27970 44322
rect 29150 44270 29202 44322
rect 33518 44270 33570 44322
rect 33966 44270 34018 44322
rect 34190 44270 34242 44322
rect 34862 44270 34914 44322
rect 35086 44270 35138 44322
rect 37550 44270 37602 44322
rect 41022 44270 41074 44322
rect 41358 44270 41410 44322
rect 42478 44270 42530 44322
rect 42702 44270 42754 44322
rect 43038 44270 43090 44322
rect 43262 44270 43314 44322
rect 43598 44270 43650 44322
rect 43822 44270 43874 44322
rect 45838 44270 45890 44322
rect 46062 44270 46114 44322
rect 46510 44270 46562 44322
rect 46622 44270 46674 44322
rect 46734 44270 46786 44322
rect 47406 44270 47458 44322
rect 48190 44270 48242 44322
rect 48526 44270 48578 44322
rect 2494 44158 2546 44210
rect 6078 44158 6130 44210
rect 17166 44158 17218 44210
rect 20302 44158 20354 44210
rect 22318 44158 22370 44210
rect 22990 44158 23042 44210
rect 29934 44158 29986 44210
rect 35870 44158 35922 44210
rect 37102 44158 37154 44210
rect 42142 44158 42194 44210
rect 44270 44158 44322 44210
rect 44830 44158 44882 44210
rect 45054 44158 45106 44210
rect 6638 44046 6690 44098
rect 12686 44046 12738 44098
rect 21646 44046 21698 44098
rect 22206 44046 22258 44098
rect 22430 44046 22482 44098
rect 22542 44046 22594 44098
rect 23102 44046 23154 44098
rect 28254 44046 28306 44098
rect 32398 44046 32450 44098
rect 32958 44046 33010 44098
rect 33406 44046 33458 44098
rect 33742 44046 33794 44098
rect 36206 44046 36258 44098
rect 40910 44046 40962 44098
rect 41246 44046 41298 44098
rect 42254 44046 42306 44098
rect 43150 44046 43202 44098
rect 43934 44046 43986 44098
rect 44046 44046 44098 44098
rect 44942 44046 44994 44098
rect 45502 44046 45554 44098
rect 47742 44046 47794 44098
rect 49198 44046 49250 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 7646 43710 7698 43762
rect 17390 43710 17442 43762
rect 30046 43710 30098 43762
rect 33966 43710 34018 43762
rect 2942 43598 2994 43650
rect 5630 43598 5682 43650
rect 6078 43598 6130 43650
rect 6190 43598 6242 43650
rect 6302 43598 6354 43650
rect 7086 43598 7138 43650
rect 7422 43598 7474 43650
rect 8206 43598 8258 43650
rect 8878 43598 8930 43650
rect 11454 43598 11506 43650
rect 23662 43598 23714 43650
rect 28254 43598 28306 43650
rect 33182 43598 33234 43650
rect 33630 43598 33682 43650
rect 35982 43598 36034 43650
rect 36094 43598 36146 43650
rect 36766 43598 36818 43650
rect 37102 43598 37154 43650
rect 46174 43598 46226 43650
rect 48974 43598 49026 43650
rect 3054 43486 3106 43538
rect 3502 43486 3554 43538
rect 6750 43486 6802 43538
rect 8766 43486 8818 43538
rect 10446 43486 10498 43538
rect 10894 43486 10946 43538
rect 11230 43486 11282 43538
rect 13918 43486 13970 43538
rect 17726 43486 17778 43538
rect 18398 43486 18450 43538
rect 24334 43486 24386 43538
rect 27246 43486 27298 43538
rect 27470 43486 27522 43538
rect 27694 43486 27746 43538
rect 27806 43486 27858 43538
rect 31166 43486 31218 43538
rect 31614 43486 31666 43538
rect 31838 43486 31890 43538
rect 34190 43486 34242 43538
rect 35198 43486 35250 43538
rect 36542 43486 36594 43538
rect 36654 43486 36706 43538
rect 36878 43486 36930 43538
rect 37550 43486 37602 43538
rect 41022 43486 41074 43538
rect 44494 43486 44546 43538
rect 44830 43486 44882 43538
rect 46734 43486 46786 43538
rect 47294 43486 47346 43538
rect 47518 43486 47570 43538
rect 3278 43374 3330 43426
rect 5294 43374 5346 43426
rect 7534 43374 7586 43426
rect 9774 43374 9826 43426
rect 14702 43374 14754 43426
rect 16830 43374 16882 43426
rect 19070 43374 19122 43426
rect 21198 43374 21250 43426
rect 21534 43374 21586 43426
rect 25902 43374 25954 43426
rect 26350 43374 26402 43426
rect 26910 43374 26962 43426
rect 27582 43374 27634 43426
rect 29150 43374 29202 43426
rect 30158 43374 30210 43426
rect 30830 43374 30882 43426
rect 31726 43374 31778 43426
rect 32174 43374 32226 43426
rect 33070 43374 33122 43426
rect 33518 43374 33570 43426
rect 34750 43374 34802 43426
rect 35646 43374 35698 43426
rect 38222 43374 38274 43426
rect 40350 43374 40402 43426
rect 41694 43374 41746 43426
rect 43822 43374 43874 43426
rect 44382 43374 44434 43426
rect 45838 43374 45890 43426
rect 47182 43374 47234 43426
rect 48078 43374 48130 43426
rect 48862 43374 48914 43426
rect 3838 43262 3890 43314
rect 3950 43262 4002 43314
rect 4174 43262 4226 43314
rect 4286 43262 4338 43314
rect 4734 43262 4786 43314
rect 5070 43262 5122 43314
rect 8094 43262 8146 43314
rect 8430 43262 8482 43314
rect 8878 43262 8930 43314
rect 9886 43262 9938 43314
rect 11118 43262 11170 43314
rect 26238 43262 26290 43314
rect 28478 43262 28530 43314
rect 28814 43262 28866 43314
rect 29374 43262 29426 43314
rect 29710 43262 29762 43314
rect 32286 43262 32338 43314
rect 44158 43262 44210 43314
rect 45054 43262 45106 43314
rect 45390 43262 45442 43314
rect 46510 43262 46562 43314
rect 47630 43262 47682 43314
rect 48750 43262 48802 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 6414 42926 6466 42978
rect 11566 42926 11618 42978
rect 19966 42926 20018 42978
rect 27358 42926 27410 42978
rect 29150 42926 29202 42978
rect 37214 42926 37266 42978
rect 37550 42926 37602 42978
rect 43374 42926 43426 42978
rect 44830 42926 44882 42978
rect 44942 42926 44994 42978
rect 45390 42926 45442 42978
rect 45614 42926 45666 42978
rect 2494 42814 2546 42866
rect 4622 42814 4674 42866
rect 6078 42814 6130 42866
rect 9886 42814 9938 42866
rect 18398 42814 18450 42866
rect 19182 42814 19234 42866
rect 23214 42814 23266 42866
rect 26910 42814 26962 42866
rect 28254 42814 28306 42866
rect 29262 42814 29314 42866
rect 30158 42814 30210 42866
rect 32734 42814 32786 42866
rect 35310 42814 35362 42866
rect 36990 42814 37042 42866
rect 42142 42814 42194 42866
rect 42590 42814 42642 42866
rect 44158 42814 44210 42866
rect 47070 42814 47122 42866
rect 49198 42814 49250 42866
rect 1822 42702 1874 42754
rect 6638 42702 6690 42754
rect 7086 42702 7138 42754
rect 10334 42702 10386 42754
rect 10782 42702 10834 42754
rect 12014 42702 12066 42754
rect 12126 42702 12178 42754
rect 12350 42702 12402 42754
rect 16830 42702 16882 42754
rect 17054 42702 17106 42754
rect 21870 42702 21922 42754
rect 22542 42702 22594 42754
rect 22878 42702 22930 42754
rect 24110 42702 24162 42754
rect 27806 42702 27858 42754
rect 27918 42702 27970 42754
rect 28142 42702 28194 42754
rect 28366 42702 28418 42754
rect 29934 42702 29986 42754
rect 30606 42702 30658 42754
rect 31950 42702 32002 42754
rect 32062 42702 32114 42754
rect 32622 42702 32674 42754
rect 33854 42702 33906 42754
rect 34862 42702 34914 42754
rect 35198 42702 35250 42754
rect 35422 42702 35474 42754
rect 35758 42702 35810 42754
rect 38334 42702 38386 42754
rect 38782 42702 38834 42754
rect 39230 42702 39282 42754
rect 42478 42702 42530 42754
rect 42814 42702 42866 42754
rect 42926 42702 42978 42754
rect 46286 42702 46338 42754
rect 7758 42590 7810 42642
rect 10222 42590 10274 42642
rect 14814 42590 14866 42642
rect 15150 42590 15202 42642
rect 16494 42590 16546 42642
rect 20078 42590 20130 42642
rect 22206 42590 22258 42642
rect 23438 42590 23490 42642
rect 24782 42590 24834 42642
rect 27246 42590 27298 42642
rect 30158 42590 30210 42642
rect 31054 42590 31106 42642
rect 33182 42590 33234 42642
rect 34190 42590 34242 42642
rect 40014 42590 40066 42642
rect 43598 42590 43650 42642
rect 44046 42590 44098 42642
rect 45054 42590 45106 42642
rect 18286 42478 18338 42530
rect 19070 42478 19122 42530
rect 21646 42478 21698 42530
rect 22094 42478 22146 42530
rect 22318 42478 22370 42530
rect 23102 42478 23154 42530
rect 23326 42478 23378 42530
rect 30382 42478 30434 42530
rect 31166 42478 31218 42530
rect 31614 42478 31666 42530
rect 31726 42478 31778 42530
rect 31838 42478 31890 42530
rect 32734 42478 32786 42530
rect 32958 42478 33010 42530
rect 33742 42478 33794 42530
rect 34414 42478 34466 42530
rect 34526 42478 34578 42530
rect 34638 42478 34690 42530
rect 35646 42478 35698 42530
rect 36430 42478 36482 42530
rect 38446 42478 38498 42530
rect 38558 42478 38610 42530
rect 38670 42478 38722 42530
rect 43486 42478 43538 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 7982 42142 8034 42194
rect 17950 42142 18002 42194
rect 22318 42142 22370 42194
rect 24670 42142 24722 42194
rect 32398 42142 32450 42194
rect 38558 42142 38610 42194
rect 39454 42142 39506 42194
rect 39678 42142 39730 42194
rect 47182 42142 47234 42194
rect 13806 42030 13858 42082
rect 16830 42030 16882 42082
rect 18958 42030 19010 42082
rect 31502 42030 31554 42082
rect 34414 42030 34466 42082
rect 39902 42030 39954 42082
rect 42702 42030 42754 42082
rect 43262 42030 43314 42082
rect 48862 42030 48914 42082
rect 6638 41918 6690 41970
rect 8206 41918 8258 41970
rect 8654 41918 8706 41970
rect 9998 41918 10050 41970
rect 13470 41918 13522 41970
rect 16382 41918 16434 41970
rect 16718 41918 16770 41970
rect 19182 41918 19234 41970
rect 23102 41918 23154 41970
rect 24558 41918 24610 41970
rect 25230 41918 25282 41970
rect 30830 41918 30882 41970
rect 31390 41918 31442 41970
rect 32510 41918 32562 41970
rect 33070 41918 33122 41970
rect 37438 41918 37490 41970
rect 38110 41918 38162 41970
rect 38894 41918 38946 41970
rect 39342 41918 39394 41970
rect 40350 41918 40402 41970
rect 41694 41918 41746 41970
rect 43038 41918 43090 41970
rect 43598 41918 43650 41970
rect 44494 41918 44546 41970
rect 44718 41918 44770 41970
rect 45726 41918 45778 41970
rect 47182 41918 47234 41970
rect 47518 41918 47570 41970
rect 49198 41918 49250 41970
rect 2270 41806 2322 41858
rect 7870 41806 7922 41858
rect 10670 41806 10722 41858
rect 12798 41806 12850 41858
rect 17390 41806 17442 41858
rect 18510 41806 18562 41858
rect 20078 41806 20130 41858
rect 22542 41806 22594 41858
rect 23550 41806 23602 41858
rect 24334 41806 24386 41858
rect 27246 41806 27298 41858
rect 31502 41806 31554 41858
rect 33518 41806 33570 41858
rect 34750 41806 34802 41858
rect 35198 41806 35250 41858
rect 39566 41806 39618 41858
rect 40238 41806 40290 41858
rect 41470 41806 41522 41858
rect 41806 41806 41858 41858
rect 43486 41806 43538 41858
rect 44942 41806 44994 41858
rect 45278 41806 45330 41858
rect 46734 41806 46786 41858
rect 48190 41806 48242 41858
rect 17614 41694 17666 41746
rect 18622 41694 18674 41746
rect 19966 41694 20018 41746
rect 22654 41694 22706 41746
rect 22878 41694 22930 41746
rect 23438 41694 23490 41746
rect 32398 41694 32450 41746
rect 33294 41694 33346 41746
rect 33966 41694 34018 41746
rect 42254 41694 42306 41746
rect 42366 41694 42418 41746
rect 42590 41694 42642 41746
rect 43822 41694 43874 41746
rect 44270 41694 44322 41746
rect 45502 41694 45554 41746
rect 45950 41694 46002 41746
rect 46398 41694 46450 41746
rect 47294 41694 47346 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 30718 41358 30770 41410
rect 36206 41358 36258 41410
rect 37102 41358 37154 41410
rect 4622 41246 4674 41298
rect 6414 41246 6466 41298
rect 9550 41246 9602 41298
rect 12910 41246 12962 41298
rect 14254 41246 14306 41298
rect 16382 41246 16434 41298
rect 17726 41246 17778 41298
rect 20078 41246 20130 41298
rect 20638 41246 20690 41298
rect 21310 41246 21362 41298
rect 23438 41246 23490 41298
rect 25566 41246 25618 41298
rect 27694 41246 27746 41298
rect 28478 41246 28530 41298
rect 30382 41246 30434 41298
rect 33966 41246 34018 41298
rect 38558 41246 38610 41298
rect 44046 41246 44098 41298
rect 47070 41246 47122 41298
rect 49198 41246 49250 41298
rect 1822 41134 1874 41186
rect 6750 41134 6802 41186
rect 6974 41134 7026 41186
rect 12462 41134 12514 41186
rect 13582 41134 13634 41186
rect 17054 41134 17106 41186
rect 17614 41134 17666 41186
rect 18174 41134 18226 41186
rect 18846 41134 18898 41186
rect 19518 41134 19570 41186
rect 20190 41134 20242 41186
rect 24110 41134 24162 41186
rect 24782 41134 24834 41186
rect 29150 41134 29202 41186
rect 29374 41134 29426 41186
rect 29486 41134 29538 41186
rect 31502 41134 31554 41186
rect 32286 41134 32338 41186
rect 33630 41134 33682 41186
rect 35198 41134 35250 41186
rect 35534 41134 35586 41186
rect 42142 41134 42194 41186
rect 44270 41134 44322 41186
rect 44830 41134 44882 41186
rect 45390 41134 45442 41186
rect 46398 41134 46450 41186
rect 2494 41022 2546 41074
rect 6526 41022 6578 41074
rect 8318 41022 8370 41074
rect 11678 41022 11730 41074
rect 18510 41022 18562 41074
rect 18734 41022 18786 41074
rect 19742 41022 19794 41074
rect 20526 41022 20578 41074
rect 28590 41022 28642 41074
rect 36318 41022 36370 41074
rect 36990 41022 37042 41074
rect 37662 41022 37714 41074
rect 43934 41022 43986 41074
rect 5742 40910 5794 40962
rect 6078 40910 6130 40962
rect 7422 40910 7474 40962
rect 7646 40910 7698 40962
rect 7982 40910 8034 40962
rect 8654 40910 8706 40962
rect 9102 40910 9154 40962
rect 12798 40910 12850 40962
rect 17950 40910 18002 40962
rect 19966 40910 20018 40962
rect 28142 40910 28194 40962
rect 29934 40910 29986 40962
rect 35310 40910 35362 40962
rect 35422 40910 35474 40962
rect 35646 40910 35698 40962
rect 36206 40910 36258 40962
rect 37998 40910 38050 40962
rect 44718 40910 44770 40962
rect 45054 40910 45106 40962
rect 45278 40910 45330 40962
rect 45950 40910 46002 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 6638 40574 6690 40626
rect 10670 40574 10722 40626
rect 17502 40574 17554 40626
rect 19854 40574 19906 40626
rect 20078 40574 20130 40626
rect 20974 40574 21026 40626
rect 21534 40574 21586 40626
rect 22990 40574 23042 40626
rect 23102 40574 23154 40626
rect 23214 40574 23266 40626
rect 23662 40574 23714 40626
rect 23998 40574 24050 40626
rect 25902 40574 25954 40626
rect 27470 40574 27522 40626
rect 27582 40574 27634 40626
rect 27694 40574 27746 40626
rect 33630 40574 33682 40626
rect 34526 40574 34578 40626
rect 39006 40574 39058 40626
rect 39902 40574 39954 40626
rect 40350 40574 40402 40626
rect 41022 40574 41074 40626
rect 42366 40574 42418 40626
rect 48974 40574 49026 40626
rect 2718 40462 2770 40514
rect 7758 40462 7810 40514
rect 8766 40462 8818 40514
rect 10894 40462 10946 40514
rect 13582 40462 13634 40514
rect 22094 40462 22146 40514
rect 22654 40462 22706 40514
rect 25454 40462 25506 40514
rect 29822 40462 29874 40514
rect 39454 40462 39506 40514
rect 41806 40462 41858 40514
rect 3726 40350 3778 40402
rect 4622 40350 4674 40402
rect 5070 40350 5122 40402
rect 5406 40350 5458 40402
rect 5742 40350 5794 40402
rect 6302 40350 6354 40402
rect 7646 40350 7698 40402
rect 8094 40350 8146 40402
rect 10334 40350 10386 40402
rect 10446 40350 10498 40402
rect 10558 40350 10610 40402
rect 16606 40350 16658 40402
rect 17726 40350 17778 40402
rect 18174 40350 18226 40402
rect 18398 40350 18450 40402
rect 19630 40350 19682 40402
rect 20302 40350 20354 40402
rect 20526 40350 20578 40402
rect 21198 40350 21250 40402
rect 21982 40350 22034 40402
rect 22878 40350 22930 40402
rect 24446 40350 24498 40402
rect 25678 40350 25730 40402
rect 26126 40350 26178 40402
rect 27358 40350 27410 40402
rect 27918 40350 27970 40402
rect 30158 40350 30210 40402
rect 31054 40350 31106 40402
rect 32174 40350 32226 40402
rect 32958 40350 33010 40402
rect 33406 40350 33458 40402
rect 34414 40350 34466 40402
rect 34638 40350 34690 40402
rect 37326 40350 37378 40402
rect 38110 40350 38162 40402
rect 38894 40350 38946 40402
rect 39230 40350 39282 40402
rect 42926 40350 42978 40402
rect 46398 40350 46450 40402
rect 2606 40238 2658 40290
rect 2942 40238 2994 40290
rect 4510 40238 4562 40290
rect 5294 40238 5346 40290
rect 6078 40238 6130 40290
rect 7982 40238 8034 40290
rect 18062 40238 18114 40290
rect 19966 40238 20018 40290
rect 21086 40238 21138 40290
rect 21646 40238 21698 40290
rect 25790 40238 25842 40290
rect 26686 40238 26738 40290
rect 28478 40238 28530 40290
rect 33518 40238 33570 40290
rect 33966 40238 34018 40290
rect 34190 40238 34242 40290
rect 35198 40238 35250 40290
rect 39118 40238 39170 40290
rect 39790 40238 39842 40290
rect 41470 40238 41522 40290
rect 42590 40238 42642 40290
rect 48974 40238 49026 40290
rect 8542 40126 8594 40178
rect 8878 40126 8930 40178
rect 24558 40126 24610 40178
rect 26798 40126 26850 40178
rect 28590 40126 28642 40178
rect 31838 40126 31890 40178
rect 41918 40126 41970 40178
rect 42254 40126 42306 40178
rect 48750 40126 48802 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 8990 39790 9042 39842
rect 13694 39790 13746 39842
rect 36430 39790 36482 39842
rect 46510 39790 46562 39842
rect 5070 39678 5122 39730
rect 9326 39678 9378 39730
rect 18734 39678 18786 39730
rect 19630 39678 19682 39730
rect 21646 39678 21698 39730
rect 22430 39678 22482 39730
rect 24558 39678 24610 39730
rect 25678 39678 25730 39730
rect 27806 39678 27858 39730
rect 42702 39678 42754 39730
rect 43374 39678 43426 39730
rect 44158 39678 44210 39730
rect 47742 39678 47794 39730
rect 48750 39678 48802 39730
rect 2158 39566 2210 39618
rect 5630 39566 5682 39618
rect 5854 39566 5906 39618
rect 6078 39566 6130 39618
rect 7310 39566 7362 39618
rect 7534 39566 7586 39618
rect 7646 39566 7698 39618
rect 7758 39566 7810 39618
rect 8206 39566 8258 39618
rect 12238 39566 12290 39618
rect 12686 39566 12738 39618
rect 14030 39566 14082 39618
rect 14254 39566 14306 39618
rect 15038 39566 15090 39618
rect 16382 39566 16434 39618
rect 16494 39566 16546 39618
rect 16942 39566 16994 39618
rect 19182 39566 19234 39618
rect 19518 39566 19570 39618
rect 19742 39566 19794 39618
rect 19966 39566 20018 39618
rect 20190 39566 20242 39618
rect 20526 39566 20578 39618
rect 21422 39566 21474 39618
rect 21870 39566 21922 39618
rect 25230 39566 25282 39618
rect 28590 39566 28642 39618
rect 34414 39566 34466 39618
rect 34862 39566 34914 39618
rect 35310 39566 35362 39618
rect 35422 39566 35474 39618
rect 36990 39566 37042 39618
rect 37214 39566 37266 39618
rect 37438 39566 37490 39618
rect 37662 39566 37714 39618
rect 37998 39566 38050 39618
rect 38670 39566 38722 39618
rect 39790 39566 39842 39618
rect 43150 39566 43202 39618
rect 43486 39566 43538 39618
rect 43710 39566 43762 39618
rect 45054 39566 45106 39618
rect 45278 39566 45330 39618
rect 45390 39566 45442 39618
rect 45726 39566 45778 39618
rect 47070 39566 47122 39618
rect 47182 39566 47234 39618
rect 47966 39566 48018 39618
rect 48190 39566 48242 39618
rect 2942 39454 2994 39506
rect 8430 39454 8482 39506
rect 8542 39454 8594 39506
rect 11454 39454 11506 39506
rect 14926 39454 14978 39506
rect 17726 39454 17778 39506
rect 18622 39454 18674 39506
rect 19070 39454 19122 39506
rect 20638 39454 20690 39506
rect 21758 39454 21810 39506
rect 29374 39454 29426 39506
rect 36318 39454 36370 39506
rect 37326 39454 37378 39506
rect 40574 39454 40626 39506
rect 43262 39454 43314 39506
rect 44830 39454 44882 39506
rect 46958 39454 47010 39506
rect 47630 39454 47682 39506
rect 48862 39454 48914 39506
rect 49086 39454 49138 39506
rect 5742 39342 5794 39394
rect 6862 39342 6914 39394
rect 12910 39342 12962 39394
rect 15150 39342 15202 39394
rect 15598 39342 15650 39394
rect 15934 39342 15986 39394
rect 16718 39342 16770 39394
rect 17502 39342 17554 39394
rect 17614 39342 17666 39394
rect 20862 39342 20914 39394
rect 21534 39342 21586 39394
rect 35534 39342 35586 39394
rect 35646 39342 35698 39394
rect 35758 39342 35810 39394
rect 38334 39342 38386 39394
rect 39006 39342 39058 39394
rect 39454 39342 39506 39394
rect 44718 39342 44770 39394
rect 46286 39342 46338 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 22990 39006 23042 39058
rect 24670 39006 24722 39058
rect 26574 39006 26626 39058
rect 26686 39006 26738 39058
rect 26910 39006 26962 39058
rect 27358 39006 27410 39058
rect 28478 39006 28530 39058
rect 32174 39006 32226 39058
rect 40350 39006 40402 39058
rect 41022 39006 41074 39058
rect 41134 39006 41186 39058
rect 41246 39006 41298 39058
rect 41358 39006 41410 39058
rect 42478 39006 42530 39058
rect 43598 39006 43650 39058
rect 44270 39006 44322 39058
rect 7646 38894 7698 38946
rect 8878 38894 8930 38946
rect 10110 38894 10162 38946
rect 13246 38894 13298 38946
rect 22654 38894 22706 38946
rect 23774 38894 23826 38946
rect 25790 38894 25842 38946
rect 26350 38894 26402 38946
rect 29934 38894 29986 38946
rect 33070 38894 33122 38946
rect 35422 38894 35474 38946
rect 36318 38894 36370 38946
rect 41582 38894 41634 38946
rect 45166 38894 45218 38946
rect 47630 38894 47682 38946
rect 48750 38894 48802 38946
rect 1822 38782 1874 38834
rect 5966 38782 6018 38834
rect 6862 38782 6914 38834
rect 7086 38782 7138 38834
rect 7534 38782 7586 38834
rect 8542 38782 8594 38834
rect 9550 38782 9602 38834
rect 9774 38782 9826 38834
rect 12462 38782 12514 38834
rect 16382 38782 16434 38834
rect 18062 38782 18114 38834
rect 20750 38782 20802 38834
rect 20974 38782 21026 38834
rect 21198 38782 21250 38834
rect 21646 38782 21698 38834
rect 21758 38782 21810 38834
rect 21982 38782 22034 38834
rect 22206 38782 22258 38834
rect 23326 38782 23378 38834
rect 23886 38782 23938 38834
rect 24334 38782 24386 38834
rect 25342 38782 25394 38834
rect 26798 38782 26850 38834
rect 27694 38782 27746 38834
rect 28142 38782 28194 38834
rect 28702 38782 28754 38834
rect 29262 38782 29314 38834
rect 34862 38782 34914 38834
rect 36654 38782 36706 38834
rect 38110 38782 38162 38834
rect 38782 38782 38834 38834
rect 43486 38782 43538 38834
rect 43934 38782 43986 38834
rect 44158 38782 44210 38834
rect 44382 38782 44434 38834
rect 44606 38782 44658 38834
rect 45838 38782 45890 38834
rect 46286 38782 46338 38834
rect 47070 38782 47122 38834
rect 47406 38782 47458 38834
rect 48078 38782 48130 38834
rect 49086 38782 49138 38834
rect 2494 38670 2546 38722
rect 4622 38670 4674 38722
rect 5294 38670 5346 38722
rect 5854 38670 5906 38722
rect 8430 38670 8482 38722
rect 15374 38670 15426 38722
rect 15710 38670 15762 38722
rect 16158 38670 16210 38722
rect 17838 38670 17890 38722
rect 18734 38670 18786 38722
rect 22094 38670 22146 38722
rect 22542 38670 22594 38722
rect 33742 38670 33794 38722
rect 34302 38670 34354 38722
rect 36206 38670 36258 38722
rect 39902 38670 39954 38722
rect 40238 38670 40290 38722
rect 42030 38670 42082 38722
rect 42926 38670 42978 38722
rect 45278 38670 45330 38722
rect 45726 38670 45778 38722
rect 48190 38670 48242 38722
rect 7534 38558 7586 38610
rect 8766 38558 8818 38610
rect 9998 38558 10050 38610
rect 18398 38558 18450 38610
rect 18846 38558 18898 38610
rect 20302 38558 20354 38610
rect 23998 38558 24050 38610
rect 33182 38558 33234 38610
rect 39790 38558 39842 38610
rect 44942 38558 44994 38610
rect 46062 38558 46114 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 2606 38222 2658 38274
rect 2942 38222 2994 38274
rect 13582 38222 13634 38274
rect 13918 38222 13970 38274
rect 21758 38222 21810 38274
rect 44942 38222 44994 38274
rect 45950 38222 46002 38274
rect 20302 38110 20354 38162
rect 22766 38110 22818 38162
rect 23326 38110 23378 38162
rect 27134 38110 27186 38162
rect 28590 38110 28642 38162
rect 29486 38110 29538 38162
rect 33966 38110 34018 38162
rect 36990 38110 37042 38162
rect 37550 38110 37602 38162
rect 39678 38110 39730 38162
rect 43710 38110 43762 38162
rect 44158 38110 44210 38162
rect 45390 38110 45442 38162
rect 47070 38110 47122 38162
rect 49198 38110 49250 38162
rect 10558 37998 10610 38050
rect 14142 37998 14194 38050
rect 14814 37998 14866 38050
rect 15150 37998 15202 38050
rect 15934 37998 15986 38050
rect 16046 37998 16098 38050
rect 16942 37998 16994 38050
rect 17166 37998 17218 38050
rect 17614 37998 17666 38050
rect 17950 37998 18002 38050
rect 18174 37998 18226 38050
rect 19518 37998 19570 38050
rect 20414 37998 20466 38050
rect 21870 37998 21922 38050
rect 22206 37998 22258 38050
rect 22430 37998 22482 38050
rect 26238 37998 26290 38050
rect 29374 37998 29426 38050
rect 29598 37998 29650 38050
rect 30046 37998 30098 38050
rect 30606 37998 30658 38050
rect 30942 37998 30994 38050
rect 35646 37998 35698 38050
rect 36206 37998 36258 38050
rect 40350 37998 40402 38050
rect 40910 37998 40962 38050
rect 45614 37998 45666 38050
rect 46286 37998 46338 38050
rect 2718 37886 2770 37938
rect 5630 37886 5682 37938
rect 10894 37886 10946 37938
rect 15374 37886 15426 37938
rect 15822 37886 15874 37938
rect 18286 37886 18338 37938
rect 18734 37886 18786 37938
rect 19070 37886 19122 37938
rect 20078 37886 20130 37938
rect 25454 37886 25506 37938
rect 26574 37886 26626 37938
rect 31726 37886 31778 37938
rect 34862 37886 34914 37938
rect 34974 37886 35026 37938
rect 35086 37886 35138 37938
rect 35758 37886 35810 37938
rect 41582 37886 41634 37938
rect 45054 37886 45106 37938
rect 5966 37774 6018 37826
rect 10782 37774 10834 37826
rect 15038 37774 15090 37826
rect 16494 37774 16546 37826
rect 17278 37774 17330 37826
rect 17390 37774 17442 37826
rect 21758 37774 21810 37826
rect 22654 37774 22706 37826
rect 22878 37774 22930 37826
rect 26686 37774 26738 37826
rect 27918 37774 27970 37826
rect 29822 37774 29874 37826
rect 34414 37774 34466 37826
rect 35870 37774 35922 37826
rect 35982 37774 36034 37826
rect 37102 37774 37154 37826
rect 44270 37774 44322 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 1934 37438 1986 37490
rect 3278 37438 3330 37490
rect 17950 37438 18002 37490
rect 18958 37438 19010 37490
rect 19182 37438 19234 37490
rect 24670 37438 24722 37490
rect 25454 37438 25506 37490
rect 26462 37438 26514 37490
rect 26574 37438 26626 37490
rect 27806 37438 27858 37490
rect 28254 37438 28306 37490
rect 28814 37438 28866 37490
rect 29934 37438 29986 37490
rect 31054 37438 31106 37490
rect 32062 37438 32114 37490
rect 32398 37438 32450 37490
rect 39678 37438 39730 37490
rect 41022 37438 41074 37490
rect 45726 37438 45778 37490
rect 3502 37326 3554 37378
rect 4622 37326 4674 37378
rect 6414 37326 6466 37378
rect 11790 37326 11842 37378
rect 16158 37326 16210 37378
rect 16382 37326 16434 37378
rect 17390 37326 17442 37378
rect 25678 37326 25730 37378
rect 29486 37326 29538 37378
rect 30494 37326 30546 37378
rect 32510 37326 32562 37378
rect 33854 37326 33906 37378
rect 37102 37326 37154 37378
rect 40238 37326 40290 37378
rect 42702 37326 42754 37378
rect 45166 37326 45218 37378
rect 45614 37326 45666 37378
rect 47966 37326 48018 37378
rect 48750 37326 48802 37378
rect 2270 37214 2322 37266
rect 3054 37214 3106 37266
rect 4958 37214 5010 37266
rect 6078 37214 6130 37266
rect 8094 37214 8146 37266
rect 8542 37214 8594 37266
rect 12462 37214 12514 37266
rect 12910 37214 12962 37266
rect 17614 37214 17666 37266
rect 18510 37214 18562 37266
rect 19742 37214 19794 37266
rect 21870 37214 21922 37266
rect 22542 37214 22594 37266
rect 23102 37214 23154 37266
rect 25230 37214 25282 37266
rect 25902 37214 25954 37266
rect 26238 37214 26290 37266
rect 26686 37214 26738 37266
rect 26798 37214 26850 37266
rect 27470 37214 27522 37266
rect 29150 37214 29202 37266
rect 31278 37214 31330 37266
rect 31726 37214 31778 37266
rect 33070 37214 33122 37266
rect 36430 37214 36482 37266
rect 39790 37214 39842 37266
rect 40014 37214 40066 37266
rect 41918 37214 41970 37266
rect 45390 37214 45442 37266
rect 46622 37214 46674 37266
rect 46846 37214 46898 37266
rect 47630 37214 47682 37266
rect 49086 37214 49138 37266
rect 9662 37102 9714 37154
rect 13694 37102 13746 37154
rect 15822 37102 15874 37154
rect 16270 37102 16322 37154
rect 19070 37102 19122 37154
rect 20750 37102 20802 37154
rect 24558 37102 24610 37154
rect 25566 37102 25618 37154
rect 35982 37102 36034 37154
rect 39230 37102 39282 37154
rect 39902 37102 39954 37154
rect 40910 37102 40962 37154
rect 41470 37102 41522 37154
rect 44830 37102 44882 37154
rect 3614 36990 3666 37042
rect 8318 36990 8370 37042
rect 8654 36990 8706 37042
rect 20638 36990 20690 37042
rect 30270 36990 30322 37042
rect 30606 36990 30658 37042
rect 46734 36990 46786 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 10894 36654 10946 36706
rect 14926 36654 14978 36706
rect 28590 36654 28642 36706
rect 46062 36654 46114 36706
rect 4622 36542 4674 36594
rect 6302 36542 6354 36594
rect 8430 36542 8482 36594
rect 10222 36542 10274 36594
rect 17614 36542 17666 36594
rect 19742 36542 19794 36594
rect 24670 36542 24722 36594
rect 26798 36542 26850 36594
rect 28030 36542 28082 36594
rect 29150 36542 29202 36594
rect 31278 36542 31330 36594
rect 32734 36542 32786 36594
rect 36430 36542 36482 36594
rect 38782 36542 38834 36594
rect 40014 36542 40066 36594
rect 45054 36542 45106 36594
rect 47070 36542 47122 36594
rect 49198 36542 49250 36594
rect 1822 36430 1874 36482
rect 9214 36430 9266 36482
rect 10558 36430 10610 36482
rect 11230 36430 11282 36482
rect 11566 36430 11618 36482
rect 11790 36430 11842 36482
rect 12686 36430 12738 36482
rect 14142 36430 14194 36482
rect 14366 36430 14418 36482
rect 14702 36430 14754 36482
rect 15262 36430 15314 36482
rect 15822 36430 15874 36482
rect 17838 36430 17890 36482
rect 19294 36430 19346 36482
rect 20078 36430 20130 36482
rect 22318 36430 22370 36482
rect 22878 36430 22930 36482
rect 23326 36430 23378 36482
rect 27582 36430 27634 36482
rect 28254 36430 28306 36482
rect 31950 36430 32002 36482
rect 33294 36430 33346 36482
rect 33630 36430 33682 36482
rect 37550 36430 37602 36482
rect 38334 36430 38386 36482
rect 38446 36430 38498 36482
rect 38670 36430 38722 36482
rect 38894 36430 38946 36482
rect 39902 36430 39954 36482
rect 40910 36430 40962 36482
rect 43486 36430 43538 36482
rect 45278 36430 45330 36482
rect 45390 36430 45442 36482
rect 45838 36430 45890 36482
rect 46286 36430 46338 36482
rect 2494 36318 2546 36370
rect 5070 36318 5122 36370
rect 13806 36318 13858 36370
rect 19182 36318 19234 36370
rect 21870 36318 21922 36370
rect 23886 36318 23938 36370
rect 34302 36318 34354 36370
rect 37326 36318 37378 36370
rect 40350 36318 40402 36370
rect 40686 36318 40738 36370
rect 41694 36318 41746 36370
rect 42814 36318 42866 36370
rect 43598 36318 43650 36370
rect 44046 36318 44098 36370
rect 4958 36206 5010 36258
rect 11454 36206 11506 36258
rect 12910 36206 12962 36258
rect 15598 36206 15650 36258
rect 18174 36206 18226 36258
rect 21646 36206 21698 36258
rect 24110 36206 24162 36258
rect 32622 36206 32674 36258
rect 32846 36206 32898 36258
rect 37886 36206 37938 36258
rect 41358 36206 41410 36258
rect 42142 36206 42194 36258
rect 43150 36206 43202 36258
rect 43822 36206 43874 36258
rect 44158 36206 44210 36258
rect 44382 36206 44434 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 2606 35870 2658 35922
rect 7758 35870 7810 35922
rect 22430 35870 22482 35922
rect 22654 35870 22706 35922
rect 22878 35870 22930 35922
rect 23998 35870 24050 35922
rect 24558 35870 24610 35922
rect 31726 35870 31778 35922
rect 32510 35870 32562 35922
rect 40126 35870 40178 35922
rect 40238 35870 40290 35922
rect 48750 35870 48802 35922
rect 49086 35870 49138 35922
rect 6638 35758 6690 35810
rect 6862 35758 6914 35810
rect 8878 35758 8930 35810
rect 15262 35758 15314 35810
rect 22094 35758 22146 35810
rect 23326 35758 23378 35810
rect 27918 35758 27970 35810
rect 33630 35758 33682 35810
rect 38670 35758 38722 35810
rect 40910 35758 40962 35810
rect 3390 35646 3442 35698
rect 7422 35646 7474 35698
rect 8318 35646 8370 35698
rect 8654 35646 8706 35698
rect 14814 35646 14866 35698
rect 15934 35646 15986 35698
rect 17726 35646 17778 35698
rect 21422 35646 21474 35698
rect 21534 35646 21586 35698
rect 21646 35646 21698 35698
rect 22542 35646 22594 35698
rect 23550 35646 23602 35698
rect 24110 35646 24162 35698
rect 27358 35646 27410 35698
rect 27582 35646 27634 35698
rect 28030 35646 28082 35698
rect 28590 35646 28642 35698
rect 30270 35646 30322 35698
rect 31614 35646 31666 35698
rect 32286 35646 32338 35698
rect 36990 35646 37042 35698
rect 39342 35646 39394 35698
rect 41246 35646 41298 35698
rect 45838 35646 45890 35698
rect 4062 35534 4114 35586
rect 6190 35534 6242 35586
rect 6526 35534 6578 35586
rect 7198 35534 7250 35586
rect 8990 35534 9042 35586
rect 9886 35534 9938 35586
rect 16158 35534 16210 35586
rect 16718 35534 16770 35586
rect 18398 35534 18450 35586
rect 20526 35534 20578 35586
rect 20974 35534 21026 35586
rect 26798 35534 26850 35586
rect 29262 35534 29314 35586
rect 29710 35534 29762 35586
rect 39454 35534 39506 35586
rect 41694 35534 41746 35586
rect 45278 35534 45330 35586
rect 48190 35534 48242 35586
rect 2270 35422 2322 35474
rect 2494 35422 2546 35474
rect 2606 35422 2658 35474
rect 7982 35422 8034 35474
rect 27022 35422 27074 35474
rect 29374 35422 29426 35474
rect 29822 35422 29874 35474
rect 30158 35422 30210 35474
rect 31726 35422 31778 35474
rect 40350 35422 40402 35474
rect 41246 35422 41298 35474
rect 47630 35422 47682 35474
rect 47966 35422 48018 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 2606 35086 2658 35138
rect 3502 35086 3554 35138
rect 9214 35086 9266 35138
rect 9326 35086 9378 35138
rect 27470 35086 27522 35138
rect 30382 35086 30434 35138
rect 44158 35086 44210 35138
rect 3166 34974 3218 35026
rect 3614 34974 3666 35026
rect 5070 34974 5122 35026
rect 8542 34974 8594 35026
rect 12686 34974 12738 35026
rect 14254 34974 14306 35026
rect 16382 34974 16434 35026
rect 18286 34974 18338 35026
rect 20414 34974 20466 35026
rect 32622 34974 32674 35026
rect 34750 34974 34802 35026
rect 35422 34974 35474 35026
rect 36094 34974 36146 35026
rect 37326 34974 37378 35026
rect 39454 34974 39506 35026
rect 41694 34974 41746 35026
rect 43822 34974 43874 35026
rect 44830 34974 44882 35026
rect 48190 34974 48242 35026
rect 49086 34974 49138 35026
rect 2942 34862 2994 34914
rect 4286 34862 4338 34914
rect 5630 34862 5682 34914
rect 8990 34862 9042 34914
rect 9886 34862 9938 34914
rect 13470 34862 13522 34914
rect 17838 34862 17890 34914
rect 18062 34862 18114 34914
rect 18846 34862 18898 34914
rect 20526 34862 20578 34914
rect 22990 34862 23042 34914
rect 28366 34862 28418 34914
rect 29486 34862 29538 34914
rect 30046 34862 30098 34914
rect 31950 34862 32002 34914
rect 35086 34862 35138 34914
rect 40238 34862 40290 34914
rect 41022 34862 41074 34914
rect 47630 34862 47682 34914
rect 48414 34862 48466 34914
rect 1934 34750 1986 34802
rect 4734 34750 4786 34802
rect 4846 34750 4898 34802
rect 6414 34750 6466 34802
rect 10558 34750 10610 34802
rect 18622 34750 18674 34802
rect 23550 34750 23602 34802
rect 27694 34750 27746 34802
rect 28030 34750 28082 34802
rect 29150 34750 29202 34802
rect 29822 34750 29874 34802
rect 44270 34750 44322 34802
rect 46958 34750 47010 34802
rect 2270 34638 2322 34690
rect 3726 34638 3778 34690
rect 4062 34638 4114 34690
rect 9326 34638 9378 34690
rect 27134 34638 27186 34690
rect 29262 34638 29314 34690
rect 35982 34638 36034 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 1934 34302 1986 34354
rect 4174 34302 4226 34354
rect 5630 34302 5682 34354
rect 6414 34302 6466 34354
rect 7758 34302 7810 34354
rect 10110 34302 10162 34354
rect 14254 34302 14306 34354
rect 18062 34302 18114 34354
rect 19854 34302 19906 34354
rect 24334 34302 24386 34354
rect 28590 34302 28642 34354
rect 29486 34302 29538 34354
rect 30382 34302 30434 34354
rect 33406 34302 33458 34354
rect 40238 34302 40290 34354
rect 41134 34302 41186 34354
rect 43934 34302 43986 34354
rect 44382 34302 44434 34354
rect 47182 34302 47234 34354
rect 47406 34302 47458 34354
rect 48190 34302 48242 34354
rect 48862 34302 48914 34354
rect 1710 34190 1762 34242
rect 2270 34190 2322 34242
rect 2718 34190 2770 34242
rect 2830 34190 2882 34242
rect 4062 34190 4114 34242
rect 6302 34190 6354 34242
rect 7310 34190 7362 34242
rect 7870 34190 7922 34242
rect 9662 34190 9714 34242
rect 11230 34190 11282 34242
rect 21646 34190 21698 34242
rect 28702 34190 28754 34242
rect 30606 34190 30658 34242
rect 31502 34190 31554 34242
rect 36206 34190 36258 34242
rect 37438 34190 37490 34242
rect 39566 34190 39618 34242
rect 39902 34190 39954 34242
rect 40910 34190 40962 34242
rect 48750 34190 48802 34242
rect 2046 34078 2098 34130
rect 2942 34078 2994 34130
rect 4398 34078 4450 34130
rect 4510 34078 4562 34130
rect 4622 34078 4674 34130
rect 5966 34078 6018 34130
rect 6638 34078 6690 34130
rect 9550 34078 9602 34130
rect 10558 34078 10610 34130
rect 14590 34078 14642 34130
rect 15934 34078 15986 34130
rect 16158 34078 16210 34130
rect 17390 34078 17442 34130
rect 20862 34078 20914 34130
rect 25230 34078 25282 34130
rect 28366 34078 28418 34130
rect 29262 34078 29314 34130
rect 29710 34078 29762 34130
rect 29934 34078 29986 34130
rect 30942 34078 30994 34130
rect 32174 34078 32226 34130
rect 33070 34078 33122 34130
rect 34750 34078 34802 34130
rect 36990 34078 37042 34130
rect 39230 34078 39282 34130
rect 42478 34078 42530 34130
rect 43038 34078 43090 34130
rect 43710 34078 43762 34130
rect 44718 34078 44770 34130
rect 45390 34078 45442 34130
rect 45502 34078 45554 34130
rect 45726 34078 45778 34130
rect 47070 34078 47122 34130
rect 49086 34078 49138 34130
rect 12126 33966 12178 34018
rect 18622 33966 18674 34018
rect 18846 33966 18898 34018
rect 19294 33966 19346 34018
rect 20414 33966 20466 34018
rect 23774 33966 23826 34018
rect 24446 33966 24498 34018
rect 26014 33966 26066 34018
rect 28142 33966 28194 34018
rect 29598 33966 29650 34018
rect 30494 33966 30546 34018
rect 31950 33966 32002 34018
rect 33966 33966 34018 34018
rect 34526 33966 34578 34018
rect 35646 33966 35698 34018
rect 38446 33966 38498 34018
rect 38894 33966 38946 34018
rect 42814 33966 42866 34018
rect 46174 33966 46226 34018
rect 46734 33966 46786 34018
rect 47630 33966 47682 34018
rect 3390 33854 3442 33906
rect 7198 33854 7250 33906
rect 7758 33854 7810 33906
rect 11566 33854 11618 33906
rect 11902 33854 11954 33906
rect 16494 33854 16546 33906
rect 17502 33854 17554 33906
rect 18958 33854 19010 33906
rect 19518 33854 19570 33906
rect 41246 33854 41298 33906
rect 44046 33854 44098 33906
rect 45838 33854 45890 33906
rect 46510 33854 46562 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 5854 33518 5906 33570
rect 6078 33518 6130 33570
rect 6302 33518 6354 33570
rect 17166 33518 17218 33570
rect 20750 33518 20802 33570
rect 28254 33518 28306 33570
rect 30382 33518 30434 33570
rect 30718 33518 30770 33570
rect 5070 33406 5122 33458
rect 8430 33406 8482 33458
rect 12686 33406 12738 33458
rect 16830 33406 16882 33458
rect 18622 33406 18674 33458
rect 19294 33406 19346 33458
rect 22094 33406 22146 33458
rect 23662 33406 23714 33458
rect 29486 33406 29538 33458
rect 33182 33406 33234 33458
rect 36430 33406 36482 33458
rect 40462 33406 40514 33458
rect 42590 33406 42642 33458
rect 43710 33406 43762 33458
rect 47070 33406 47122 33458
rect 49198 33406 49250 33458
rect 2158 33294 2210 33346
rect 5630 33294 5682 33346
rect 7310 33294 7362 33346
rect 7982 33294 8034 33346
rect 8878 33294 8930 33346
rect 9102 33294 9154 33346
rect 9326 33294 9378 33346
rect 9886 33294 9938 33346
rect 15150 33294 15202 33346
rect 16270 33294 16322 33346
rect 18174 33294 18226 33346
rect 20190 33294 20242 33346
rect 20414 33294 20466 33346
rect 24782 33294 24834 33346
rect 26462 33294 26514 33346
rect 27246 33294 27298 33346
rect 27358 33294 27410 33346
rect 27582 33294 27634 33346
rect 28142 33294 28194 33346
rect 28478 33294 28530 33346
rect 29374 33294 29426 33346
rect 29598 33294 29650 33346
rect 29822 33294 29874 33346
rect 30158 33294 30210 33346
rect 31838 33294 31890 33346
rect 33630 33294 33682 33346
rect 36990 33294 37042 33346
rect 43374 33294 43426 33346
rect 44830 33294 44882 33346
rect 45390 33294 45442 33346
rect 46398 33294 46450 33346
rect 2942 33182 2994 33234
rect 6414 33182 6466 33234
rect 6974 33182 7026 33234
rect 7758 33182 7810 33234
rect 9438 33182 9490 33234
rect 10558 33182 10610 33234
rect 13806 33182 13858 33234
rect 15710 33182 15762 33234
rect 16158 33182 16210 33234
rect 16382 33182 16434 33234
rect 17390 33182 17442 33234
rect 19294 33182 19346 33234
rect 19406 33182 19458 33234
rect 19630 33182 19682 33234
rect 24670 33182 24722 33234
rect 25902 33182 25954 33234
rect 32062 33182 32114 33234
rect 34302 33182 34354 33234
rect 37774 33182 37826 33234
rect 45054 33182 45106 33234
rect 45166 33182 45218 33234
rect 45838 33182 45890 33234
rect 6862 33070 6914 33122
rect 7534 33070 7586 33122
rect 13470 33070 13522 33122
rect 15374 33070 15426 33122
rect 18286 33070 18338 33122
rect 18510 33070 18562 33122
rect 18622 33070 18674 33122
rect 19070 33070 19122 33122
rect 26798 33070 26850 33122
rect 27918 33070 27970 33122
rect 29262 33070 29314 33122
rect 31166 33070 31218 33122
rect 32846 33070 32898 33122
rect 40014 33070 40066 33122
rect 43822 33070 43874 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 3166 32734 3218 32786
rect 11006 32734 11058 32786
rect 15710 32734 15762 32786
rect 19294 32734 19346 32786
rect 19406 32734 19458 32786
rect 19742 32734 19794 32786
rect 20078 32734 20130 32786
rect 20862 32734 20914 32786
rect 25790 32734 25842 32786
rect 27470 32734 27522 32786
rect 28702 32734 28754 32786
rect 33294 32734 33346 32786
rect 34302 32734 34354 32786
rect 40910 32734 40962 32786
rect 44942 32734 44994 32786
rect 45166 32734 45218 32786
rect 45278 32734 45330 32786
rect 46286 32734 46338 32786
rect 47294 32734 47346 32786
rect 5518 32622 5570 32674
rect 10110 32622 10162 32674
rect 13134 32622 13186 32674
rect 17502 32622 17554 32674
rect 17614 32622 17666 32674
rect 18062 32622 18114 32674
rect 20302 32622 20354 32674
rect 20414 32622 20466 32674
rect 26910 32622 26962 32674
rect 27022 32622 27074 32674
rect 27694 32622 27746 32674
rect 27806 32622 27858 32674
rect 28254 32622 28306 32674
rect 29374 32622 29426 32674
rect 29710 32622 29762 32674
rect 34750 32622 34802 32674
rect 42142 32622 42194 32674
rect 45502 32622 45554 32674
rect 48078 32622 48130 32674
rect 48750 32622 48802 32674
rect 1822 32510 1874 32562
rect 2270 32510 2322 32562
rect 3278 32510 3330 32562
rect 8878 32510 8930 32562
rect 9774 32510 9826 32562
rect 10222 32510 10274 32562
rect 10782 32510 10834 32562
rect 11118 32510 11170 32562
rect 12462 32510 12514 32562
rect 16494 32510 16546 32562
rect 16606 32510 16658 32562
rect 16830 32510 16882 32562
rect 17278 32510 17330 32562
rect 18286 32510 18338 32562
rect 18510 32510 18562 32562
rect 18734 32510 18786 32562
rect 19518 32510 19570 32562
rect 21198 32510 21250 32562
rect 21534 32510 21586 32562
rect 25566 32510 25618 32562
rect 27246 32510 27298 32562
rect 28478 32510 28530 32562
rect 28926 32510 28978 32562
rect 31502 32510 31554 32562
rect 32062 32510 32114 32562
rect 34190 32510 34242 32562
rect 34526 32510 34578 32562
rect 38894 32510 38946 32562
rect 41470 32510 41522 32562
rect 44718 32510 44770 32562
rect 46622 32510 46674 32562
rect 47070 32510 47122 32562
rect 47406 32510 47458 32562
rect 47630 32510 47682 32562
rect 47966 32510 48018 32562
rect 49086 32510 49138 32562
rect 3054 32398 3106 32450
rect 10446 32398 10498 32450
rect 15262 32398 15314 32450
rect 15598 32398 15650 32450
rect 18622 32398 18674 32450
rect 22318 32398 22370 32450
rect 24446 32398 24498 32450
rect 28814 32398 28866 32450
rect 29822 32398 29874 32450
rect 30718 32398 30770 32450
rect 31278 32398 31330 32450
rect 32622 32398 32674 32450
rect 33182 32398 33234 32450
rect 33742 32398 33794 32450
rect 34414 32398 34466 32450
rect 36206 32398 36258 32450
rect 41022 32398 41074 32450
rect 44270 32398 44322 32450
rect 45726 32398 45778 32450
rect 2046 32286 2098 32338
rect 2382 32286 2434 32338
rect 2830 32286 2882 32338
rect 9438 32286 9490 32338
rect 16046 32286 16098 32338
rect 26462 32286 26514 32338
rect 29262 32286 29314 32338
rect 33630 32286 33682 32338
rect 46286 32286 46338 32338
rect 46398 32286 46450 32338
rect 48078 32286 48130 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 20190 31950 20242 32002
rect 22542 31950 22594 32002
rect 2494 31838 2546 31890
rect 4622 31838 4674 31890
rect 6638 31838 6690 31890
rect 8766 31838 8818 31890
rect 9214 31838 9266 31890
rect 9774 31838 9826 31890
rect 19630 31838 19682 31890
rect 23886 31838 23938 31890
rect 27470 31838 27522 31890
rect 28030 31838 28082 31890
rect 29934 31838 29986 31890
rect 30382 31838 30434 31890
rect 33070 31838 33122 31890
rect 35198 31838 35250 31890
rect 35870 31838 35922 31890
rect 38446 31838 38498 31890
rect 39118 31838 39170 31890
rect 44830 31838 44882 31890
rect 44942 31838 44994 31890
rect 47070 31838 47122 31890
rect 49198 31838 49250 31890
rect 1822 31726 1874 31778
rect 5966 31726 6018 31778
rect 9550 31726 9602 31778
rect 9998 31726 10050 31778
rect 10446 31726 10498 31778
rect 11006 31726 11058 31778
rect 13582 31726 13634 31778
rect 19182 31726 19234 31778
rect 19854 31726 19906 31778
rect 20526 31726 20578 31778
rect 21870 31726 21922 31778
rect 22430 31726 22482 31778
rect 22990 31726 23042 31778
rect 23438 31726 23490 31778
rect 24558 31726 24610 31778
rect 30046 31726 30098 31778
rect 30718 31726 30770 31778
rect 31390 31726 31442 31778
rect 32398 31726 32450 31778
rect 35982 31726 36034 31778
rect 40014 31726 40066 31778
rect 41134 31726 41186 31778
rect 41694 31726 41746 31778
rect 42254 31726 42306 31778
rect 42926 31726 42978 31778
rect 44270 31726 44322 31778
rect 45166 31726 45218 31778
rect 45726 31726 45778 31778
rect 46286 31726 46338 31778
rect 10110 31614 10162 31666
rect 10670 31614 10722 31666
rect 17502 31614 17554 31666
rect 20750 31614 20802 31666
rect 22094 31614 22146 31666
rect 22542 31614 22594 31666
rect 25342 31614 25394 31666
rect 27918 31614 27970 31666
rect 29374 31614 29426 31666
rect 30942 31614 30994 31666
rect 31278 31614 31330 31666
rect 31614 31614 31666 31666
rect 31838 31614 31890 31666
rect 35534 31614 35586 31666
rect 37326 31614 37378 31666
rect 37774 31614 37826 31666
rect 38782 31614 38834 31666
rect 42478 31614 42530 31666
rect 43038 31614 43090 31666
rect 45614 31614 45666 31666
rect 10782 31502 10834 31554
rect 19406 31502 19458 31554
rect 19630 31502 19682 31554
rect 21534 31502 21586 31554
rect 28478 31502 28530 31554
rect 29598 31502 29650 31554
rect 29822 31502 29874 31554
rect 35758 31502 35810 31554
rect 36094 31502 36146 31554
rect 37214 31502 37266 31554
rect 37438 31502 37490 31554
rect 37550 31502 37602 31554
rect 38222 31502 38274 31554
rect 38334 31502 38386 31554
rect 38558 31502 38610 31554
rect 39678 31502 39730 31554
rect 40574 31502 40626 31554
rect 41246 31502 41298 31554
rect 41358 31502 41410 31554
rect 41470 31502 41522 31554
rect 43150 31502 43202 31554
rect 45502 31502 45554 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 2382 31166 2434 31218
rect 9550 31166 9602 31218
rect 9886 31166 9938 31218
rect 16830 31166 16882 31218
rect 17390 31166 17442 31218
rect 17614 31166 17666 31218
rect 18062 31166 18114 31218
rect 18734 31166 18786 31218
rect 19182 31166 19234 31218
rect 20750 31166 20802 31218
rect 25566 31166 25618 31218
rect 26686 31166 26738 31218
rect 27134 31166 27186 31218
rect 30942 31166 30994 31218
rect 31726 31166 31778 31218
rect 34078 31166 34130 31218
rect 34750 31166 34802 31218
rect 43486 31166 43538 31218
rect 45614 31166 45666 31218
rect 45838 31166 45890 31218
rect 48750 31166 48802 31218
rect 49086 31166 49138 31218
rect 4622 31054 4674 31106
rect 6302 31054 6354 31106
rect 6414 31054 6466 31106
rect 6638 31054 6690 31106
rect 8206 31054 8258 31106
rect 8654 31054 8706 31106
rect 16718 31054 16770 31106
rect 17838 31054 17890 31106
rect 18286 31054 18338 31106
rect 18398 31054 18450 31106
rect 20302 31054 20354 31106
rect 25902 31054 25954 31106
rect 30494 31054 30546 31106
rect 31950 31054 32002 31106
rect 34414 31054 34466 31106
rect 37998 31054 38050 31106
rect 42590 31054 42642 31106
rect 44046 31054 44098 31106
rect 46958 31054 47010 31106
rect 2606 30942 2658 30994
rect 3502 30942 3554 30994
rect 4062 30942 4114 30994
rect 4510 30942 4562 30994
rect 4846 30942 4898 30994
rect 6078 30942 6130 30994
rect 7758 30942 7810 30994
rect 7982 30942 8034 30994
rect 8318 30942 8370 30994
rect 13022 30942 13074 30994
rect 13470 30942 13522 30994
rect 20078 30942 20130 30994
rect 21422 30942 21474 30994
rect 31502 30942 31554 30994
rect 31726 30942 31778 30994
rect 33854 30942 33906 30994
rect 35310 30942 35362 30994
rect 40910 30942 40962 30994
rect 41022 30942 41074 30994
rect 41358 30942 41410 30994
rect 43598 30942 43650 30994
rect 46062 30942 46114 30994
rect 46510 30942 46562 30994
rect 47630 30942 47682 30994
rect 47742 30942 47794 30994
rect 47966 30942 48018 30994
rect 48078 30942 48130 30994
rect 2270 30830 2322 30882
rect 6862 30830 6914 30882
rect 7534 30830 7586 30882
rect 10222 30830 10274 30882
rect 12350 30830 12402 30882
rect 14254 30830 14306 30882
rect 16382 30830 16434 30882
rect 18846 30830 18898 30882
rect 19294 30830 19346 30882
rect 20638 30830 20690 30882
rect 22094 30830 22146 30882
rect 24222 30830 24274 30882
rect 24670 30830 24722 30882
rect 27694 30830 27746 30882
rect 28142 30830 28194 30882
rect 28590 30830 28642 30882
rect 29150 30830 29202 30882
rect 29710 30830 29762 30882
rect 30046 30830 30098 30882
rect 32622 30830 32674 30882
rect 33294 30830 33346 30882
rect 45838 30830 45890 30882
rect 46286 30830 46338 30882
rect 47854 30830 47906 30882
rect 2942 30718 2994 30770
rect 3054 30718 3106 30770
rect 3278 30718 3330 30770
rect 7198 30718 7250 30770
rect 17726 30718 17778 30770
rect 29934 30718 29986 30770
rect 33406 30718 33458 30770
rect 46846 30718 46898 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 28142 30382 28194 30434
rect 43486 30382 43538 30434
rect 47406 30382 47458 30434
rect 48862 30382 48914 30434
rect 2494 30270 2546 30322
rect 4622 30270 4674 30322
rect 7086 30270 7138 30322
rect 9214 30270 9266 30322
rect 11342 30270 11394 30322
rect 24110 30270 24162 30322
rect 32062 30270 32114 30322
rect 33070 30270 33122 30322
rect 36990 30270 37042 30322
rect 41582 30270 41634 30322
rect 43262 30270 43314 30322
rect 43934 30270 43986 30322
rect 45054 30270 45106 30322
rect 48302 30270 48354 30322
rect 1822 30158 1874 30210
rect 5966 30158 6018 30210
rect 6414 30158 6466 30210
rect 6974 30158 7026 30210
rect 7198 30158 7250 30210
rect 8094 30158 8146 30210
rect 12126 30158 12178 30210
rect 12686 30158 12738 30210
rect 13806 30158 13858 30210
rect 14478 30158 14530 30210
rect 14702 30158 14754 30210
rect 20638 30158 20690 30210
rect 21870 30158 21922 30210
rect 23774 30158 23826 30210
rect 25566 30158 25618 30210
rect 26238 30158 26290 30210
rect 27358 30158 27410 30210
rect 27694 30158 27746 30210
rect 27918 30158 27970 30210
rect 28366 30158 28418 30210
rect 28702 30158 28754 30210
rect 31054 30158 31106 30210
rect 35198 30158 35250 30210
rect 35982 30158 36034 30210
rect 36318 30158 36370 30210
rect 39790 30158 39842 30210
rect 40686 30158 40738 30210
rect 41134 30158 41186 30210
rect 42030 30158 42082 30210
rect 42254 30158 42306 30210
rect 42814 30158 42866 30210
rect 42926 30158 42978 30210
rect 43710 30158 43762 30210
rect 44830 30158 44882 30210
rect 45278 30158 45330 30210
rect 46062 30158 46114 30210
rect 46398 30158 46450 30210
rect 46846 30158 46898 30210
rect 47070 30158 47122 30210
rect 47406 30158 47458 30210
rect 48190 30158 48242 30210
rect 48414 30158 48466 30210
rect 48526 30158 48578 30210
rect 7422 30046 7474 30098
rect 7870 30046 7922 30098
rect 12462 30046 12514 30098
rect 14142 30046 14194 30098
rect 18398 30046 18450 30098
rect 22654 30046 22706 30098
rect 22990 30046 23042 30098
rect 23326 30046 23378 30098
rect 26798 30046 26850 30098
rect 31614 30046 31666 30098
rect 36430 30046 36482 30098
rect 39118 30046 39170 30098
rect 40350 30046 40402 30098
rect 40462 30046 40514 30098
rect 45054 30046 45106 30098
rect 45502 30046 45554 30098
rect 47742 30046 47794 30098
rect 5630 29934 5682 29986
rect 6638 29934 6690 29986
rect 15038 29934 15090 29986
rect 21422 29934 21474 29986
rect 21646 29934 21698 29986
rect 21758 29934 21810 29986
rect 22430 29934 22482 29986
rect 25006 29934 25058 29986
rect 26462 29934 26514 29986
rect 28142 29934 28194 29986
rect 29374 29934 29426 29986
rect 29710 29934 29762 29986
rect 30270 29934 30322 29986
rect 30718 29934 30770 29986
rect 32510 29934 32562 29986
rect 42702 29934 42754 29986
rect 44382 29934 44434 29986
rect 45726 29934 45778 29986
rect 45950 29934 46002 29986
rect 46622 29934 46674 29986
rect 46734 29934 46786 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 3278 29598 3330 29650
rect 5294 29598 5346 29650
rect 7646 29598 7698 29650
rect 12686 29598 12738 29650
rect 23886 29598 23938 29650
rect 24782 29598 24834 29650
rect 34750 29598 34802 29650
rect 34974 29598 35026 29650
rect 35086 29598 35138 29650
rect 36430 29598 36482 29650
rect 36542 29598 36594 29650
rect 40350 29598 40402 29650
rect 41022 29598 41074 29650
rect 41134 29598 41186 29650
rect 41358 29598 41410 29650
rect 42478 29598 42530 29650
rect 42702 29598 42754 29650
rect 48750 29598 48802 29650
rect 4846 29486 4898 29538
rect 8318 29486 8370 29538
rect 8766 29486 8818 29538
rect 10670 29486 10722 29538
rect 21422 29486 21474 29538
rect 31726 29486 31778 29538
rect 33406 29486 33458 29538
rect 34862 29486 34914 29538
rect 36654 29486 36706 29538
rect 42366 29486 42418 29538
rect 46174 29486 46226 29538
rect 48862 29486 48914 29538
rect 3166 29374 3218 29426
rect 3502 29374 3554 29426
rect 3726 29374 3778 29426
rect 3950 29374 4002 29426
rect 4286 29374 4338 29426
rect 4622 29374 4674 29426
rect 4958 29374 5010 29426
rect 5518 29374 5570 29426
rect 7310 29374 7362 29426
rect 7982 29374 8034 29426
rect 11006 29374 11058 29426
rect 13918 29374 13970 29426
rect 17502 29374 17554 29426
rect 20750 29374 20802 29426
rect 23998 29374 24050 29426
rect 25230 29374 25282 29426
rect 31390 29374 31442 29426
rect 32174 29374 32226 29426
rect 33070 29374 33122 29426
rect 33742 29374 33794 29426
rect 33966 29374 34018 29426
rect 34414 29374 34466 29426
rect 35198 29374 35250 29426
rect 35982 29374 36034 29426
rect 36766 29374 36818 29426
rect 12126 29262 12178 29314
rect 14702 29262 14754 29314
rect 16830 29262 16882 29314
rect 18174 29262 18226 29314
rect 20302 29262 20354 29314
rect 23550 29262 23602 29314
rect 27470 29262 27522 29314
rect 30830 29262 30882 29314
rect 37662 29374 37714 29426
rect 37886 29374 37938 29426
rect 38334 29374 38386 29426
rect 39342 29374 39394 29426
rect 39902 29374 39954 29426
rect 40910 29374 40962 29426
rect 42926 29374 42978 29426
rect 33854 29262 33906 29314
rect 36990 29262 37042 29314
rect 38446 29262 38498 29314
rect 41918 29262 41970 29314
rect 8654 29150 8706 29202
rect 8990 29150 9042 29202
rect 12350 29150 12402 29202
rect 31054 29150 31106 29202
rect 35646 29150 35698 29202
rect 35982 29150 36034 29202
rect 38558 29150 38610 29202
rect 41806 29150 41858 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 5966 28814 6018 28866
rect 21310 28814 21362 28866
rect 22542 28814 22594 28866
rect 35758 28814 35810 28866
rect 43150 28814 43202 28866
rect 44830 28814 44882 28866
rect 45166 28814 45218 28866
rect 47742 28814 47794 28866
rect 4286 28702 4338 28754
rect 6414 28702 6466 28754
rect 10446 28702 10498 28754
rect 12574 28702 12626 28754
rect 15150 28702 15202 28754
rect 23102 28702 23154 28754
rect 29150 28702 29202 28754
rect 35310 28702 35362 28754
rect 41582 28702 41634 28754
rect 46510 28702 46562 28754
rect 47070 28702 47122 28754
rect 48750 28702 48802 28754
rect 3278 28590 3330 28642
rect 3390 28590 3442 28642
rect 3950 28590 4002 28642
rect 4510 28590 4562 28642
rect 4734 28590 4786 28642
rect 8542 28590 8594 28642
rect 9214 28590 9266 28642
rect 9662 28590 9714 28642
rect 14702 28590 14754 28642
rect 14926 28590 14978 28642
rect 15710 28590 15762 28642
rect 17054 28590 17106 28642
rect 18734 28590 18786 28642
rect 19406 28590 19458 28642
rect 19854 28590 19906 28642
rect 20638 28590 20690 28642
rect 21758 28590 21810 28642
rect 21870 28590 21922 28642
rect 21982 28590 22034 28642
rect 23214 28590 23266 28642
rect 26350 28590 26402 28642
rect 27694 28590 27746 28642
rect 28590 28590 28642 28642
rect 31278 28590 31330 28642
rect 32062 28590 32114 28642
rect 32398 28590 32450 28642
rect 35870 28590 35922 28642
rect 36094 28590 36146 28642
rect 37326 28590 37378 28642
rect 38670 28590 38722 28642
rect 40462 28590 40514 28642
rect 42590 28590 42642 28642
rect 43038 28590 43090 28642
rect 45166 28590 45218 28642
rect 45502 28590 45554 28642
rect 46062 28590 46114 28642
rect 48078 28590 48130 28642
rect 48414 28590 48466 28642
rect 49198 28590 49250 28642
rect 3502 28478 3554 28530
rect 4174 28478 4226 28530
rect 5854 28478 5906 28530
rect 5966 28478 6018 28530
rect 15486 28478 15538 28530
rect 16718 28478 16770 28530
rect 17726 28478 17778 28530
rect 17838 28478 17890 28530
rect 18286 28478 18338 28530
rect 20190 28478 20242 28530
rect 22430 28478 22482 28530
rect 22542 28478 22594 28530
rect 24670 28478 24722 28530
rect 25790 28478 25842 28530
rect 26798 28478 26850 28530
rect 27358 28478 27410 28530
rect 28478 28478 28530 28530
rect 33182 28478 33234 28530
rect 36990 28478 37042 28530
rect 39118 28478 39170 28530
rect 40350 28478 40402 28530
rect 43150 28478 43202 28530
rect 44046 28478 44098 28530
rect 46174 28478 46226 28530
rect 46958 28478 47010 28530
rect 47182 28478 47234 28530
rect 47406 28478 47458 28530
rect 47854 28478 47906 28530
rect 16606 28366 16658 28418
rect 17166 28366 17218 28418
rect 18062 28366 18114 28418
rect 18510 28366 18562 28418
rect 26910 28366 26962 28418
rect 27582 28366 27634 28418
rect 27806 28366 27858 28418
rect 27918 28366 27970 28418
rect 44158 28366 44210 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 6414 28030 6466 28082
rect 11118 28030 11170 28082
rect 16270 28030 16322 28082
rect 16382 28030 16434 28082
rect 18398 28030 18450 28082
rect 19630 28030 19682 28082
rect 20750 28030 20802 28082
rect 21086 28030 21138 28082
rect 26014 28030 26066 28082
rect 26574 28030 26626 28082
rect 26686 28030 26738 28082
rect 26910 28030 26962 28082
rect 31726 28030 31778 28082
rect 35758 28030 35810 28082
rect 48078 28030 48130 28082
rect 4958 27918 5010 27970
rect 6526 27918 6578 27970
rect 7422 27918 7474 27970
rect 7758 27918 7810 27970
rect 8206 27918 8258 27970
rect 13806 27918 13858 27970
rect 14030 27918 14082 27970
rect 16606 27918 16658 27970
rect 17502 27918 17554 27970
rect 18622 27918 18674 27970
rect 25342 27918 25394 27970
rect 28142 27918 28194 27970
rect 32062 27918 32114 27970
rect 33518 27918 33570 27970
rect 33630 27918 33682 27970
rect 33854 27918 33906 27970
rect 34078 27918 34130 27970
rect 1822 27806 1874 27858
rect 5518 27806 5570 27858
rect 5966 27806 6018 27858
rect 7086 27806 7138 27858
rect 8654 27806 8706 27858
rect 11678 27806 11730 27858
rect 12574 27806 12626 27858
rect 15038 27806 15090 27858
rect 15262 27806 15314 27858
rect 16046 27806 16098 27858
rect 16158 27806 16210 27858
rect 17390 27806 17442 27858
rect 17950 27806 18002 27858
rect 18174 27806 18226 27858
rect 18958 27806 19010 27858
rect 19182 27806 19234 27858
rect 19406 27806 19458 27858
rect 19854 27806 19906 27858
rect 21422 27806 21474 27858
rect 24670 27806 24722 27858
rect 26350 27806 26402 27858
rect 26798 27806 26850 27858
rect 27470 27806 27522 27858
rect 31166 27806 31218 27858
rect 32286 27806 32338 27858
rect 32510 27806 32562 27858
rect 34414 27806 34466 27858
rect 34638 27806 34690 27858
rect 35086 27806 35138 27858
rect 36542 27806 36594 27858
rect 36878 27806 36930 27858
rect 38222 27806 38274 27858
rect 38446 27806 38498 27858
rect 38782 27806 38834 27858
rect 39118 27806 39170 27858
rect 44718 27806 44770 27858
rect 46846 27806 46898 27858
rect 2494 27694 2546 27746
rect 4622 27694 4674 27746
rect 7870 27694 7922 27746
rect 8318 27694 8370 27746
rect 11454 27694 11506 27746
rect 12014 27694 12066 27746
rect 12798 27694 12850 27746
rect 13694 27694 13746 27746
rect 14926 27694 14978 27746
rect 19742 27694 19794 27746
rect 21758 27694 21810 27746
rect 23886 27694 23938 27746
rect 25230 27694 25282 27746
rect 30270 27694 30322 27746
rect 30718 27694 30770 27746
rect 32174 27694 32226 27746
rect 33070 27694 33122 27746
rect 36318 27694 36370 27746
rect 44158 27694 44210 27746
rect 47070 27694 47122 27746
rect 47630 27694 47682 27746
rect 48190 27694 48242 27746
rect 48862 27694 48914 27746
rect 6862 27582 6914 27634
rect 8542 27582 8594 27634
rect 14478 27582 14530 27634
rect 17502 27582 17554 27634
rect 18398 27582 18450 27634
rect 33182 27582 33234 27634
rect 37550 27582 37602 27634
rect 46510 27582 46562 27634
rect 47518 27582 47570 27634
rect 48750 27582 48802 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 2494 27246 2546 27298
rect 4510 27246 4562 27298
rect 6078 27246 6130 27298
rect 6414 27246 6466 27298
rect 15934 27246 15986 27298
rect 17390 27246 17442 27298
rect 17614 27246 17666 27298
rect 44942 27246 44994 27298
rect 2606 27134 2658 27186
rect 5070 27134 5122 27186
rect 6638 27134 6690 27186
rect 12798 27134 12850 27186
rect 13470 27134 13522 27186
rect 14366 27134 14418 27186
rect 15374 27134 15426 27186
rect 15822 27134 15874 27186
rect 17166 27134 17218 27186
rect 18622 27134 18674 27186
rect 19406 27134 19458 27186
rect 19854 27134 19906 27186
rect 21310 27134 21362 27186
rect 24894 27134 24946 27186
rect 27022 27134 27074 27186
rect 29486 27134 29538 27186
rect 38334 27134 38386 27186
rect 40014 27134 40066 27186
rect 42142 27134 42194 27186
rect 42814 27134 42866 27186
rect 44046 27134 44098 27186
rect 45390 27134 45442 27186
rect 45838 27134 45890 27186
rect 49198 27134 49250 27186
rect 3278 27022 3330 27074
rect 3726 27022 3778 27074
rect 3950 27022 4002 27074
rect 4174 27022 4226 27074
rect 4846 27022 4898 27074
rect 12238 27022 12290 27074
rect 13918 27022 13970 27074
rect 14814 27022 14866 27074
rect 15262 27022 15314 27074
rect 16606 27022 16658 27074
rect 18286 27022 18338 27074
rect 18734 27022 18786 27074
rect 18958 27022 19010 27074
rect 19294 27022 19346 27074
rect 20750 27022 20802 27074
rect 24222 27022 24274 27074
rect 27806 27022 27858 27074
rect 29150 27022 29202 27074
rect 36206 27022 36258 27074
rect 36990 27022 37042 27074
rect 37326 27022 37378 27074
rect 39342 27022 39394 27074
rect 42478 27022 42530 27074
rect 43486 27022 43538 27074
rect 46286 27022 46338 27074
rect 2942 26910 2994 26962
rect 3614 26910 3666 26962
rect 8430 26910 8482 26962
rect 16382 26910 16434 26962
rect 16830 26910 16882 26962
rect 18510 26910 18562 26962
rect 20414 26910 20466 26962
rect 23438 26910 23490 26962
rect 29374 26910 29426 26962
rect 29598 26910 29650 26962
rect 30382 26910 30434 26962
rect 32398 26910 32450 26962
rect 37102 26910 37154 26962
rect 37662 26910 37714 26962
rect 37998 26910 38050 26962
rect 43710 26910 43762 26962
rect 43934 26910 43986 26962
rect 44830 26910 44882 26962
rect 47070 26910 47122 26962
rect 15038 26798 15090 26850
rect 15374 26798 15426 26850
rect 16718 26798 16770 26850
rect 18062 26798 18114 26850
rect 28254 26798 28306 26850
rect 29710 26798 29762 26850
rect 30718 26798 30770 26850
rect 38894 26798 38946 26850
rect 42702 26798 42754 26850
rect 42926 26798 42978 26850
rect 43038 26798 43090 26850
rect 44046 26798 44098 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 5182 26462 5234 26514
rect 14926 26462 14978 26514
rect 16494 26462 16546 26514
rect 17614 26462 17666 26514
rect 19742 26462 19794 26514
rect 20974 26462 21026 26514
rect 21422 26462 21474 26514
rect 28478 26462 28530 26514
rect 30270 26462 30322 26514
rect 31614 26462 31666 26514
rect 32062 26462 32114 26514
rect 32510 26462 32562 26514
rect 46062 26462 46114 26514
rect 46510 26462 46562 26514
rect 47630 26462 47682 26514
rect 47742 26462 47794 26514
rect 2494 26350 2546 26402
rect 13246 26350 13298 26402
rect 13582 26350 13634 26402
rect 14030 26350 14082 26402
rect 15710 26350 15762 26402
rect 17390 26350 17442 26402
rect 17838 26350 17890 26402
rect 29150 26350 29202 26402
rect 30158 26350 30210 26402
rect 30494 26350 30546 26402
rect 39790 26350 39842 26402
rect 44606 26350 44658 26402
rect 46622 26350 46674 26402
rect 46846 26350 46898 26402
rect 48078 26350 48130 26402
rect 1822 26238 1874 26290
rect 4958 26238 5010 26290
rect 6190 26238 6242 26290
rect 9550 26238 9602 26290
rect 13134 26238 13186 26290
rect 13694 26238 13746 26290
rect 14254 26238 14306 26290
rect 14590 26238 14642 26290
rect 15150 26238 15202 26290
rect 15822 26238 15874 26290
rect 16158 26238 16210 26290
rect 16382 26238 16434 26290
rect 16606 26238 16658 26290
rect 16830 26238 16882 26290
rect 18062 26238 18114 26290
rect 18398 26238 18450 26290
rect 24670 26238 24722 26290
rect 28142 26238 28194 26290
rect 28814 26238 28866 26290
rect 29486 26238 29538 26290
rect 30606 26238 30658 26290
rect 35982 26238 36034 26290
rect 39230 26238 39282 26290
rect 42142 26238 42194 26290
rect 45390 26238 45442 26290
rect 45726 26238 45778 26290
rect 47070 26238 47122 26290
rect 47518 26238 47570 26290
rect 47854 26238 47906 26290
rect 4622 26126 4674 26178
rect 6862 26126 6914 26178
rect 8990 26126 9042 26178
rect 10334 26126 10386 26178
rect 12462 26126 12514 26178
rect 14142 26126 14194 26178
rect 17726 26126 17778 26178
rect 18510 26126 18562 26178
rect 19294 26126 19346 26178
rect 21310 26126 21362 26178
rect 21758 26126 21810 26178
rect 23886 26126 23938 26178
rect 25230 26126 25282 26178
rect 27358 26126 27410 26178
rect 31054 26126 31106 26178
rect 33070 26126 33122 26178
rect 35198 26126 35250 26178
rect 36318 26126 36370 26178
rect 38446 26126 38498 26178
rect 39678 26126 39730 26178
rect 40350 26126 40402 26178
rect 41470 26126 41522 26178
rect 42478 26126 42530 26178
rect 46734 26126 46786 26178
rect 48862 26126 48914 26178
rect 5294 26014 5346 26066
rect 12686 26014 12738 26066
rect 39566 26014 39618 26066
rect 48750 26014 48802 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 4174 25678 4226 25730
rect 4846 25678 4898 25730
rect 6078 25678 6130 25730
rect 6750 25678 6802 25730
rect 7198 25678 7250 25730
rect 14478 25678 14530 25730
rect 14926 25678 14978 25730
rect 15374 25678 15426 25730
rect 23102 25678 23154 25730
rect 26798 25678 26850 25730
rect 32734 25678 32786 25730
rect 33070 25678 33122 25730
rect 5854 25566 5906 25618
rect 6862 25566 6914 25618
rect 14366 25566 14418 25618
rect 15262 25566 15314 25618
rect 17950 25566 18002 25618
rect 22094 25566 22146 25618
rect 25902 25566 25954 25618
rect 32062 25566 32114 25618
rect 33518 25566 33570 25618
rect 35534 25566 35586 25618
rect 36990 25566 37042 25618
rect 37998 25566 38050 25618
rect 46958 25566 47010 25618
rect 49086 25566 49138 25618
rect 5070 25454 5122 25506
rect 7086 25454 7138 25506
rect 7982 25454 8034 25506
rect 8430 25454 8482 25506
rect 8654 25454 8706 25506
rect 9774 25454 9826 25506
rect 10446 25454 10498 25506
rect 10782 25454 10834 25506
rect 11006 25454 11058 25506
rect 12238 25454 12290 25506
rect 12462 25454 12514 25506
rect 16270 25454 16322 25506
rect 16718 25454 16770 25506
rect 16942 25454 16994 25506
rect 17502 25454 17554 25506
rect 18734 25454 18786 25506
rect 19630 25454 19682 25506
rect 20414 25454 20466 25506
rect 20526 25454 20578 25506
rect 20750 25454 20802 25506
rect 21982 25454 22034 25506
rect 22206 25454 22258 25506
rect 22542 25454 22594 25506
rect 23438 25454 23490 25506
rect 23886 25454 23938 25506
rect 23998 25454 24050 25506
rect 24782 25454 24834 25506
rect 25454 25454 25506 25506
rect 27358 25454 27410 25506
rect 27582 25454 27634 25506
rect 27806 25454 27858 25506
rect 28030 25454 28082 25506
rect 29262 25454 29314 25506
rect 33742 25454 33794 25506
rect 33966 25454 34018 25506
rect 34302 25454 34354 25506
rect 34526 25454 34578 25506
rect 34638 25454 34690 25506
rect 35646 25454 35698 25506
rect 35870 25454 35922 25506
rect 36318 25454 36370 25506
rect 37214 25454 37266 25506
rect 37774 25454 37826 25506
rect 38334 25454 38386 25506
rect 40350 25454 40402 25506
rect 40798 25454 40850 25506
rect 42926 25454 42978 25506
rect 44270 25454 44322 25506
rect 45278 25454 45330 25506
rect 45502 25454 45554 25506
rect 46286 25454 46338 25506
rect 6414 25342 6466 25394
rect 7646 25342 7698 25394
rect 8318 25342 8370 25394
rect 10110 25342 10162 25394
rect 12126 25342 12178 25394
rect 14814 25342 14866 25394
rect 16046 25342 16098 25394
rect 18174 25342 18226 25394
rect 18286 25342 18338 25394
rect 20078 25342 20130 25394
rect 21310 25342 21362 25394
rect 22990 25342 23042 25394
rect 23774 25342 23826 25394
rect 25118 25342 25170 25394
rect 26686 25342 26738 25394
rect 27694 25342 27746 25394
rect 29934 25342 29986 25394
rect 32846 25342 32898 25394
rect 33406 25342 33458 25394
rect 35086 25342 35138 25394
rect 36430 25342 36482 25394
rect 38222 25342 38274 25394
rect 38894 25342 38946 25394
rect 41918 25342 41970 25394
rect 43598 25342 43650 25394
rect 45838 25342 45890 25394
rect 3950 25230 4002 25282
rect 4062 25230 4114 25282
rect 4510 25230 4562 25282
rect 15934 25230 15986 25282
rect 16830 25230 16882 25282
rect 19742 25230 19794 25282
rect 20302 25230 20354 25282
rect 21422 25230 21474 25282
rect 22430 25230 22482 25282
rect 23662 25230 23714 25282
rect 24446 25230 24498 25282
rect 26462 25230 26514 25282
rect 28590 25230 28642 25282
rect 35534 25230 35586 25282
rect 37550 25230 37602 25282
rect 40462 25230 40514 25282
rect 43150 25230 43202 25282
rect 43262 25230 43314 25282
rect 43374 25230 43426 25282
rect 43934 25230 43986 25282
rect 45390 25230 45442 25282
rect 45614 25230 45666 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 5854 24894 5906 24946
rect 8430 24894 8482 24946
rect 15598 24894 15650 24946
rect 22654 24894 22706 24946
rect 22766 24894 22818 24946
rect 22990 24894 23042 24946
rect 24446 24894 24498 24946
rect 31054 24894 31106 24946
rect 31614 24894 31666 24946
rect 31838 24894 31890 24946
rect 32622 24894 32674 24946
rect 41358 24894 41410 24946
rect 47182 24894 47234 24946
rect 5406 24782 5458 24834
rect 7646 24782 7698 24834
rect 9998 24782 10050 24834
rect 13806 24782 13858 24834
rect 14590 24782 14642 24834
rect 16158 24782 16210 24834
rect 16270 24782 16322 24834
rect 16830 24782 16882 24834
rect 22430 24782 22482 24834
rect 30830 24782 30882 24834
rect 36654 24782 36706 24834
rect 39230 24782 39282 24834
rect 41582 24782 41634 24834
rect 41694 24782 41746 24834
rect 41918 24782 41970 24834
rect 45838 24782 45890 24834
rect 46286 24782 46338 24834
rect 46734 24782 46786 24834
rect 1822 24670 1874 24722
rect 5182 24670 5234 24722
rect 5294 24670 5346 24722
rect 6302 24670 6354 24722
rect 6638 24670 6690 24722
rect 7982 24670 8034 24722
rect 10334 24670 10386 24722
rect 12126 24670 12178 24722
rect 12574 24670 12626 24722
rect 13134 24670 13186 24722
rect 14030 24670 14082 24722
rect 15038 24670 15090 24722
rect 15262 24670 15314 24722
rect 15486 24670 15538 24722
rect 16382 24670 16434 24722
rect 18174 24670 18226 24722
rect 19406 24670 19458 24722
rect 20750 24670 20802 24722
rect 22878 24670 22930 24722
rect 23886 24670 23938 24722
rect 25230 24670 25282 24722
rect 31390 24670 31442 24722
rect 32062 24670 32114 24722
rect 33182 24670 33234 24722
rect 36318 24670 36370 24722
rect 40014 24670 40066 24722
rect 41470 24670 41522 24722
rect 45054 24670 45106 24722
rect 45502 24670 45554 24722
rect 48078 24670 48130 24722
rect 2494 24558 2546 24610
rect 4622 24558 4674 24610
rect 6190 24558 6242 24610
rect 11902 24558 11954 24610
rect 12462 24558 12514 24610
rect 14702 24558 14754 24610
rect 15598 24558 15650 24610
rect 18622 24558 18674 24610
rect 20974 24558 21026 24610
rect 30046 24558 30098 24610
rect 33854 24558 33906 24610
rect 35982 24558 36034 24610
rect 37102 24558 37154 24610
rect 42254 24558 42306 24610
rect 44382 24558 44434 24610
rect 46174 24558 46226 24610
rect 47630 24558 47682 24610
rect 48862 24558 48914 24610
rect 6526 24446 6578 24498
rect 11790 24446 11842 24498
rect 21646 24446 21698 24498
rect 30718 24446 30770 24498
rect 31502 24446 31554 24498
rect 36318 24446 36370 24498
rect 46622 24446 46674 24498
rect 48750 24446 48802 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 12574 24110 12626 24162
rect 12910 24110 12962 24162
rect 13470 24110 13522 24162
rect 14814 24110 14866 24162
rect 15710 24110 15762 24162
rect 34862 24110 34914 24162
rect 38446 24110 38498 24162
rect 4622 23998 4674 24050
rect 6078 23998 6130 24050
rect 6638 23998 6690 24050
rect 7870 23998 7922 24050
rect 8206 23998 8258 24050
rect 9886 23998 9938 24050
rect 12014 23998 12066 24050
rect 12350 23998 12402 24050
rect 15486 23998 15538 24050
rect 16046 23998 16098 24050
rect 17054 23998 17106 24050
rect 17838 23998 17890 24050
rect 19966 23998 20018 24050
rect 21534 23998 21586 24050
rect 29262 23998 29314 24050
rect 32958 23998 33010 24050
rect 36094 23998 36146 24050
rect 36430 23998 36482 24050
rect 37550 23998 37602 24050
rect 37998 23998 38050 24050
rect 39006 23998 39058 24050
rect 39902 23998 39954 24050
rect 40686 23998 40738 24050
rect 45614 23998 45666 24050
rect 47742 23998 47794 24050
rect 48414 23998 48466 24050
rect 49198 23998 49250 24050
rect 1822 23886 1874 23938
rect 5630 23886 5682 23938
rect 7758 23886 7810 23938
rect 9102 23886 9154 23938
rect 13918 23886 13970 23938
rect 14254 23886 14306 23938
rect 16382 23886 16434 23938
rect 17502 23886 17554 23938
rect 20750 23886 20802 23938
rect 25454 23886 25506 23938
rect 27470 23886 27522 23938
rect 27694 23886 27746 23938
rect 28030 23886 28082 23938
rect 28366 23886 28418 23938
rect 29822 23886 29874 23938
rect 30158 23886 30210 23938
rect 34414 23886 34466 23938
rect 34974 23886 35026 23938
rect 35198 23886 35250 23938
rect 35422 23886 35474 23938
rect 37326 23886 37378 23938
rect 38558 23886 38610 23938
rect 43486 23886 43538 23938
rect 44158 23886 44210 23938
rect 44830 23886 44882 23938
rect 48190 23886 48242 23938
rect 48302 23886 48354 23938
rect 2494 23774 2546 23826
rect 5854 23774 5906 23826
rect 6190 23774 6242 23826
rect 14030 23774 14082 23826
rect 14590 23774 14642 23826
rect 16718 23774 16770 23826
rect 30830 23774 30882 23826
rect 33854 23774 33906 23826
rect 42814 23774 42866 23826
rect 43934 23774 43986 23826
rect 48526 23774 48578 23826
rect 48750 23774 48802 23826
rect 8766 23662 8818 23714
rect 15150 23662 15202 23714
rect 26910 23662 26962 23714
rect 27022 23662 27074 23714
rect 27134 23662 27186 23714
rect 27806 23662 27858 23714
rect 29150 23662 29202 23714
rect 29374 23662 29426 23714
rect 33518 23662 33570 23714
rect 33742 23662 33794 23714
rect 34526 23662 34578 23714
rect 38446 23662 38498 23714
rect 39454 23662 39506 23714
rect 40350 23662 40402 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 10446 23326 10498 23378
rect 11790 23326 11842 23378
rect 15822 23326 15874 23378
rect 16494 23326 16546 23378
rect 25342 23326 25394 23378
rect 29150 23326 29202 23378
rect 29822 23326 29874 23378
rect 30270 23326 30322 23378
rect 30382 23326 30434 23378
rect 31166 23326 31218 23378
rect 31502 23326 31554 23378
rect 32622 23326 32674 23378
rect 33294 23326 33346 23378
rect 35086 23326 35138 23378
rect 36542 23326 36594 23378
rect 36990 23326 37042 23378
rect 37214 23326 37266 23378
rect 38894 23326 38946 23378
rect 41022 23326 41074 23378
rect 41134 23326 41186 23378
rect 41806 23326 41858 23378
rect 42030 23326 42082 23378
rect 3390 23214 3442 23266
rect 4286 23214 4338 23266
rect 5742 23214 5794 23266
rect 6862 23214 6914 23266
rect 11678 23214 11730 23266
rect 12014 23214 12066 23266
rect 12238 23214 12290 23266
rect 13358 23214 13410 23266
rect 16606 23214 16658 23266
rect 19182 23214 19234 23266
rect 19630 23214 19682 23266
rect 23438 23214 23490 23266
rect 26462 23214 26514 23266
rect 28926 23214 28978 23266
rect 30494 23214 30546 23266
rect 31950 23214 32002 23266
rect 35422 23214 35474 23266
rect 36878 23214 36930 23266
rect 37550 23214 37602 23266
rect 38222 23214 38274 23266
rect 40910 23214 40962 23266
rect 44942 23214 44994 23266
rect 3614 23102 3666 23154
rect 4062 23102 4114 23154
rect 4398 23102 4450 23154
rect 4622 23102 4674 23154
rect 4846 23102 4898 23154
rect 5070 23102 5122 23154
rect 5294 23102 5346 23154
rect 5406 23102 5458 23154
rect 6190 23102 6242 23154
rect 10782 23102 10834 23154
rect 11006 23102 11058 23154
rect 12686 23102 12738 23154
rect 16046 23102 16098 23154
rect 18958 23102 19010 23154
rect 19406 23102 19458 23154
rect 19966 23102 20018 23154
rect 20190 23102 20242 23154
rect 20638 23102 20690 23154
rect 24222 23102 24274 23154
rect 25678 23102 25730 23154
rect 29486 23102 29538 23154
rect 30942 23102 30994 23154
rect 34190 23102 34242 23154
rect 37886 23102 37938 23154
rect 38334 23102 38386 23154
rect 43374 23102 43426 23154
rect 3502 22990 3554 23042
rect 8990 22990 9042 23042
rect 15486 22990 15538 23042
rect 18062 22990 18114 23042
rect 18510 22990 18562 23042
rect 20078 22990 20130 23042
rect 20974 22990 21026 23042
rect 21310 22990 21362 23042
rect 24670 22990 24722 23042
rect 28590 22990 28642 23042
rect 33630 22990 33682 23042
rect 33854 22990 33906 23042
rect 34750 22990 34802 23042
rect 35982 22990 36034 23042
rect 39230 22990 39282 23042
rect 39678 22990 39730 23042
rect 40126 22990 40178 23042
rect 42590 22990 42642 23042
rect 48862 22990 48914 23042
rect 19070 22878 19122 22930
rect 29262 22878 29314 22930
rect 31950 22878 32002 22930
rect 32622 22878 32674 22930
rect 34526 22878 34578 22930
rect 36206 22878 36258 22930
rect 48750 22878 48802 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 4622 22430 4674 22482
rect 9102 22430 9154 22482
rect 17054 22430 17106 22482
rect 17278 22430 17330 22482
rect 20638 22430 20690 22482
rect 21422 22430 21474 22482
rect 21758 22430 21810 22482
rect 28142 22430 28194 22482
rect 29262 22430 29314 22482
rect 30382 22430 30434 22482
rect 33294 22542 33346 22594
rect 33630 22542 33682 22594
rect 37774 22542 37826 22594
rect 38894 22542 38946 22594
rect 32062 22430 32114 22482
rect 32398 22430 32450 22482
rect 34638 22430 34690 22482
rect 41694 22430 41746 22482
rect 42590 22430 42642 22482
rect 43374 22430 43426 22482
rect 44158 22430 44210 22482
rect 44942 22430 44994 22482
rect 47070 22430 47122 22482
rect 49198 22430 49250 22482
rect 1822 22318 1874 22370
rect 6638 22318 6690 22370
rect 11342 22318 11394 22370
rect 20190 22318 20242 22370
rect 24670 22318 24722 22370
rect 25342 22318 25394 22370
rect 29934 22318 29986 22370
rect 31838 22318 31890 22370
rect 33966 22318 34018 22370
rect 34190 22318 34242 22370
rect 35198 22318 35250 22370
rect 38334 22318 38386 22370
rect 38558 22318 38610 22370
rect 39566 22318 39618 22370
rect 40686 22318 40738 22370
rect 41358 22318 41410 22370
rect 42142 22318 42194 22370
rect 43822 22318 43874 22370
rect 45166 22318 45218 22370
rect 45950 22318 46002 22370
rect 46286 22318 46338 22370
rect 2494 22206 2546 22258
rect 19406 22206 19458 22258
rect 23886 22206 23938 22258
rect 26014 22206 26066 22258
rect 29598 22206 29650 22258
rect 31390 22206 31442 22258
rect 31614 22206 31666 22258
rect 32174 22206 32226 22258
rect 32622 22206 32674 22258
rect 33070 22206 33122 22258
rect 35534 22206 35586 22258
rect 37102 22206 37154 22258
rect 37214 22206 37266 22258
rect 37326 22206 37378 22258
rect 39230 22206 39282 22258
rect 40014 22206 40066 22258
rect 43262 22206 43314 22258
rect 28590 22094 28642 22146
rect 30942 22094 30994 22146
rect 36094 22094 36146 22146
rect 36430 22094 36482 22146
rect 39902 22094 39954 22146
rect 40910 22094 40962 22146
rect 45502 22094 45554 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 2718 21758 2770 21810
rect 8766 21758 8818 21810
rect 9662 21758 9714 21810
rect 14030 21758 14082 21810
rect 20862 21758 20914 21810
rect 26350 21758 26402 21810
rect 26462 21758 26514 21810
rect 27470 21758 27522 21810
rect 27918 21758 27970 21810
rect 30606 21758 30658 21810
rect 33070 21758 33122 21810
rect 2830 21646 2882 21698
rect 10222 21646 10274 21698
rect 10558 21646 10610 21698
rect 10894 21646 10946 21698
rect 19518 21646 19570 21698
rect 21198 21646 21250 21698
rect 27694 21646 27746 21698
rect 5518 21534 5570 21586
rect 8542 21534 8594 21586
rect 8878 21534 8930 21586
rect 9774 21534 9826 21586
rect 11454 21534 11506 21586
rect 12462 21534 12514 21586
rect 13358 21534 13410 21586
rect 14254 21534 14306 21586
rect 16046 21534 16098 21586
rect 20302 21534 20354 21586
rect 21086 21534 21138 21586
rect 21310 21534 21362 21586
rect 21758 21534 21810 21586
rect 25342 21534 25394 21586
rect 25790 21534 25842 21586
rect 26014 21534 26066 21586
rect 26574 21534 26626 21586
rect 27022 21534 27074 21586
rect 27134 21534 27186 21586
rect 6190 21422 6242 21474
rect 8318 21422 8370 21474
rect 11230 21422 11282 21474
rect 11790 21422 11842 21474
rect 12126 21422 12178 21474
rect 13134 21422 13186 21474
rect 16494 21422 16546 21474
rect 16830 21422 16882 21474
rect 17390 21422 17442 21474
rect 22430 21422 22482 21474
rect 24558 21422 24610 21474
rect 25902 21422 25954 21474
rect 33294 21758 33346 21810
rect 34078 21758 34130 21810
rect 35982 21758 36034 21810
rect 36654 21758 36706 21810
rect 46846 21758 46898 21810
rect 47294 21758 47346 21810
rect 47742 21758 47794 21810
rect 29598 21646 29650 21698
rect 29710 21646 29762 21698
rect 31950 21646 32002 21698
rect 36206 21646 36258 21698
rect 46062 21646 46114 21698
rect 46958 21646 47010 21698
rect 28254 21534 28306 21586
rect 28478 21534 28530 21586
rect 28702 21534 28754 21586
rect 29822 21534 29874 21586
rect 30270 21534 30322 21586
rect 31278 21534 31330 21586
rect 31390 21534 31442 21586
rect 31502 21534 31554 21586
rect 33742 21534 33794 21586
rect 34190 21534 34242 21586
rect 35086 21534 35138 21586
rect 35534 21534 35586 21586
rect 36542 21534 36594 21586
rect 36766 21534 36818 21586
rect 37102 21534 37154 21586
rect 37550 21534 37602 21586
rect 41358 21534 41410 21586
rect 42478 21534 42530 21586
rect 45838 21534 45890 21586
rect 46398 21534 46450 21586
rect 46734 21534 46786 21586
rect 47518 21534 47570 21586
rect 48750 21534 48802 21586
rect 28366 21422 28418 21474
rect 32398 21422 32450 21474
rect 33182 21422 33234 21474
rect 34638 21422 34690 21474
rect 38222 21422 38274 21474
rect 40350 21422 40402 21474
rect 41022 21422 41074 21474
rect 41806 21422 41858 21474
rect 43262 21422 43314 21474
rect 45390 21422 45442 21474
rect 47406 21422 47458 21474
rect 9662 21310 9714 21362
rect 13694 21310 13746 21362
rect 27358 21310 27410 21362
rect 27918 21310 27970 21362
rect 29150 21310 29202 21362
rect 34078 21310 34130 21362
rect 35422 21310 35474 21362
rect 35870 21310 35922 21362
rect 40910 21310 40962 21362
rect 48750 21310 48802 21362
rect 49086 21310 49138 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 17950 20974 18002 21026
rect 34414 20974 34466 21026
rect 34862 20974 34914 21026
rect 35086 20974 35138 21026
rect 35422 20974 35474 21026
rect 38334 20974 38386 21026
rect 4622 20862 4674 20914
rect 9662 20862 9714 20914
rect 10782 20862 10834 20914
rect 12910 20862 12962 20914
rect 17054 20862 17106 20914
rect 18174 20862 18226 20914
rect 19294 20862 19346 20914
rect 21422 20862 21474 20914
rect 22318 20862 22370 20914
rect 22766 20862 22818 20914
rect 24558 20862 24610 20914
rect 26686 20862 26738 20914
rect 30718 20862 30770 20914
rect 32846 20862 32898 20914
rect 39454 20862 39506 20914
rect 40126 20862 40178 20914
rect 47070 20862 47122 20914
rect 49198 20862 49250 20914
rect 1822 20750 1874 20802
rect 6526 20750 6578 20802
rect 6750 20750 6802 20802
rect 10110 20750 10162 20802
rect 14142 20750 14194 20802
rect 17390 20750 17442 20802
rect 18398 20750 18450 20802
rect 18734 20750 18786 20802
rect 18958 20750 19010 20802
rect 19742 20750 19794 20802
rect 21534 20750 21586 20802
rect 21758 20750 21810 20802
rect 22654 20750 22706 20802
rect 22878 20750 22930 20802
rect 23886 20750 23938 20802
rect 27246 20750 27298 20802
rect 28030 20750 28082 20802
rect 29486 20750 29538 20802
rect 30046 20750 30098 20802
rect 33630 20750 33682 20802
rect 34190 20750 34242 20802
rect 35982 20750 36034 20802
rect 36318 20750 36370 20802
rect 37102 20750 37154 20802
rect 37326 20750 37378 20802
rect 38334 20750 38386 20802
rect 38670 20750 38722 20802
rect 39230 20750 39282 20802
rect 39678 20750 39730 20802
rect 39790 20750 39842 20802
rect 40350 20750 40402 20802
rect 42030 20750 42082 20802
rect 43150 20750 43202 20802
rect 45726 20750 45778 20802
rect 46286 20750 46338 20802
rect 2494 20638 2546 20690
rect 5854 20638 5906 20690
rect 6078 20638 6130 20690
rect 7534 20638 7586 20690
rect 14926 20638 14978 20690
rect 17726 20638 17778 20690
rect 20414 20638 20466 20690
rect 20750 20638 20802 20690
rect 27022 20638 27074 20690
rect 27582 20638 27634 20690
rect 35198 20638 35250 20690
rect 35758 20638 35810 20690
rect 37438 20638 37490 20690
rect 40462 20638 40514 20690
rect 41022 20638 41074 20690
rect 42366 20638 42418 20690
rect 42702 20638 42754 20690
rect 43710 20638 43762 20690
rect 44046 20638 44098 20690
rect 44942 20638 44994 20690
rect 45950 20638 46002 20690
rect 6190 20526 6242 20578
rect 17838 20526 17890 20578
rect 19630 20526 19682 20578
rect 21310 20526 21362 20578
rect 23102 20526 23154 20578
rect 27358 20526 27410 20578
rect 28254 20526 28306 20578
rect 29598 20526 29650 20578
rect 29710 20526 29762 20578
rect 33854 20526 33906 20578
rect 34078 20526 34130 20578
rect 34750 20526 34802 20578
rect 35870 20526 35922 20578
rect 37886 20526 37938 20578
rect 42254 20526 42306 20578
rect 42478 20526 42530 20578
rect 43262 20526 43314 20578
rect 43374 20526 43426 20578
rect 43486 20526 43538 20578
rect 44158 20526 44210 20578
rect 45054 20526 45106 20578
rect 45390 20526 45442 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 3054 20190 3106 20242
rect 8318 20190 8370 20242
rect 9662 20190 9714 20242
rect 23998 20190 24050 20242
rect 41246 20190 41298 20242
rect 2494 20078 2546 20130
rect 2718 20078 2770 20130
rect 7422 20078 7474 20130
rect 8878 20078 8930 20130
rect 13470 20078 13522 20130
rect 15374 20078 15426 20130
rect 16270 20078 16322 20130
rect 16382 20078 16434 20130
rect 22654 20078 22706 20130
rect 23774 20078 23826 20130
rect 24334 20078 24386 20130
rect 24670 20078 24722 20130
rect 41582 20078 41634 20130
rect 44382 20078 44434 20130
rect 46734 20078 46786 20130
rect 47406 20078 47458 20130
rect 49086 20078 49138 20130
rect 2382 19966 2434 20018
rect 2830 19966 2882 20018
rect 3166 19966 3218 20018
rect 3502 19966 3554 20018
rect 3950 19966 4002 20018
rect 7310 19966 7362 20018
rect 8430 19966 8482 20018
rect 9438 19966 9490 20018
rect 9774 19966 9826 20018
rect 14366 19966 14418 20018
rect 14478 19966 14530 20018
rect 14702 19966 14754 20018
rect 15598 19966 15650 20018
rect 15934 19966 15986 20018
rect 16046 19966 16098 20018
rect 21982 19966 22034 20018
rect 22878 19966 22930 20018
rect 23326 19966 23378 20018
rect 23438 19966 23490 20018
rect 25566 19966 25618 20018
rect 34190 19966 34242 20018
rect 34414 19966 34466 20018
rect 35086 19966 35138 20018
rect 40910 19966 40962 20018
rect 41134 19966 41186 20018
rect 41358 19966 41410 20018
rect 45166 19966 45218 20018
rect 45502 19966 45554 20018
rect 45726 19966 45778 20018
rect 46174 19966 46226 20018
rect 46622 19966 46674 20018
rect 47854 19966 47906 20018
rect 48190 19966 48242 20018
rect 48750 19966 48802 20018
rect 4622 19854 4674 19906
rect 6750 19854 6802 19906
rect 15374 19854 15426 19906
rect 16830 19854 16882 19906
rect 17502 19854 17554 19906
rect 18062 19854 18114 19906
rect 18734 19854 18786 19906
rect 19070 19854 19122 19906
rect 21198 19854 21250 19906
rect 22766 19854 22818 19906
rect 23662 19854 23714 19906
rect 27358 19854 27410 19906
rect 31166 19854 31218 19906
rect 31614 19854 31666 19906
rect 32062 19854 32114 19906
rect 32510 19854 32562 19906
rect 33182 19854 33234 19906
rect 40126 19854 40178 19906
rect 42254 19854 42306 19906
rect 45614 19854 45666 19906
rect 13582 19742 13634 19794
rect 13918 19742 13970 19794
rect 16718 19742 16770 19794
rect 17838 19742 17890 19794
rect 31054 19742 31106 19794
rect 33854 19742 33906 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 25678 19406 25730 19458
rect 4622 19294 4674 19346
rect 18398 19294 18450 19346
rect 21422 19294 21474 19346
rect 25006 19294 25058 19346
rect 28254 19294 28306 19346
rect 29710 19294 29762 19346
rect 30494 19294 30546 19346
rect 31278 19294 31330 19346
rect 34302 19294 34354 19346
rect 36430 19294 36482 19346
rect 42926 19294 42978 19346
rect 45054 19294 45106 19346
rect 47070 19294 47122 19346
rect 49198 19294 49250 19346
rect 1822 19182 1874 19234
rect 7422 19182 7474 19234
rect 8318 19182 8370 19234
rect 8542 19182 8594 19234
rect 8990 19182 9042 19234
rect 13694 19182 13746 19234
rect 14030 19182 14082 19234
rect 14702 19182 14754 19234
rect 14814 19182 14866 19234
rect 14926 19182 14978 19234
rect 20078 19182 20130 19234
rect 21310 19182 21362 19234
rect 21534 19182 21586 19234
rect 21870 19182 21922 19234
rect 22094 19182 22146 19234
rect 22430 19182 22482 19234
rect 22766 19182 22818 19234
rect 23214 19182 23266 19234
rect 23998 19182 24050 19234
rect 26126 19182 26178 19234
rect 26238 19182 26290 19234
rect 26462 19182 26514 19234
rect 26798 19182 26850 19234
rect 27246 19182 27298 19234
rect 27918 19182 27970 19234
rect 29150 19182 29202 19234
rect 29598 19182 29650 19234
rect 30158 19182 30210 19234
rect 30606 19182 30658 19234
rect 32622 19182 32674 19234
rect 33630 19182 33682 19234
rect 41918 19182 41970 19234
rect 43038 19182 43090 19234
rect 43262 19182 43314 19234
rect 44046 19182 44098 19234
rect 45502 19182 45554 19234
rect 46286 19182 46338 19234
rect 2494 19070 2546 19122
rect 5630 19070 5682 19122
rect 5854 19070 5906 19122
rect 6190 19070 6242 19122
rect 6414 19070 6466 19122
rect 6638 19070 6690 19122
rect 6750 19070 6802 19122
rect 7646 19070 7698 19122
rect 7758 19070 7810 19122
rect 9326 19070 9378 19122
rect 9438 19070 9490 19122
rect 12126 19070 12178 19122
rect 13806 19070 13858 19122
rect 22990 19070 23042 19122
rect 23662 19070 23714 19122
rect 25342 19070 25394 19122
rect 28254 19070 28306 19122
rect 30830 19070 30882 19122
rect 31166 19070 31218 19122
rect 31390 19070 31442 19122
rect 33070 19070 33122 19122
rect 39566 19070 39618 19122
rect 43486 19070 43538 19122
rect 45950 19070 46002 19122
rect 5966 18958 6018 19010
rect 8654 18958 8706 19010
rect 9102 18958 9154 19010
rect 9998 18958 10050 19010
rect 11790 18958 11842 19010
rect 12686 18958 12738 19010
rect 14254 18958 14306 19010
rect 22206 18958 22258 19010
rect 24446 18958 24498 19010
rect 29374 18958 29426 19010
rect 29710 18958 29762 19010
rect 30382 18958 30434 19010
rect 31838 18958 31890 19010
rect 32174 18958 32226 19010
rect 33182 18958 33234 19010
rect 42926 18958 42978 19010
rect 44158 18958 44210 19010
rect 44382 18958 44434 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 5070 18622 5122 18674
rect 5294 18622 5346 18674
rect 6638 18622 6690 18674
rect 14254 18622 14306 18674
rect 16606 18622 16658 18674
rect 17390 18622 17442 18674
rect 17614 18622 17666 18674
rect 19406 18622 19458 18674
rect 21086 18622 21138 18674
rect 31390 18622 31442 18674
rect 41022 18622 41074 18674
rect 48750 18622 48802 18674
rect 2494 18510 2546 18562
rect 2606 18510 2658 18562
rect 2942 18510 2994 18562
rect 3054 18510 3106 18562
rect 3278 18510 3330 18562
rect 4510 18510 4562 18562
rect 4622 18510 4674 18562
rect 4958 18510 5010 18562
rect 5518 18510 5570 18562
rect 7758 18510 7810 18562
rect 8318 18510 8370 18562
rect 8542 18510 8594 18562
rect 9662 18510 9714 18562
rect 9774 18510 9826 18562
rect 11790 18510 11842 18562
rect 17726 18510 17778 18562
rect 18510 18510 18562 18562
rect 18622 18510 18674 18562
rect 19182 18510 19234 18562
rect 31278 18510 31330 18562
rect 32062 18510 32114 18562
rect 37550 18510 37602 18562
rect 38670 18510 38722 18562
rect 42590 18510 42642 18562
rect 46510 18510 46562 18562
rect 47518 18510 47570 18562
rect 2270 18398 2322 18450
rect 3390 18398 3442 18450
rect 3726 18398 3778 18450
rect 3950 18398 4002 18450
rect 5854 18398 5906 18450
rect 6862 18398 6914 18450
rect 7422 18398 7474 18450
rect 8990 18398 9042 18450
rect 9438 18398 9490 18450
rect 11118 18398 11170 18450
rect 14590 18398 14642 18450
rect 14814 18398 14866 18450
rect 15262 18398 15314 18450
rect 15374 18398 15426 18450
rect 15598 18398 15650 18450
rect 15822 18398 15874 18450
rect 16270 18398 16322 18450
rect 16382 18398 16434 18450
rect 16494 18398 16546 18450
rect 16830 18398 16882 18450
rect 18062 18398 18114 18450
rect 19294 18398 19346 18450
rect 19742 18398 19794 18450
rect 24222 18398 24274 18450
rect 25342 18398 25394 18450
rect 25790 18398 25842 18450
rect 27358 18398 27410 18450
rect 28030 18398 28082 18450
rect 30718 18398 30770 18450
rect 31166 18398 31218 18450
rect 31502 18398 31554 18450
rect 31726 18398 31778 18450
rect 32286 18398 32338 18450
rect 33294 18398 33346 18450
rect 33966 18398 34018 18450
rect 36430 18398 36482 18450
rect 36990 18398 37042 18450
rect 40238 18398 40290 18450
rect 40910 18398 40962 18450
rect 41134 18398 41186 18450
rect 42030 18398 42082 18450
rect 46174 18398 46226 18450
rect 46734 18398 46786 18450
rect 47966 18398 48018 18450
rect 48974 18398 49026 18450
rect 3614 18286 3666 18338
rect 8766 18286 8818 18338
rect 10222 18286 10274 18338
rect 10670 18286 10722 18338
rect 13918 18286 13970 18338
rect 15710 18286 15762 18338
rect 18174 18286 18226 18338
rect 20190 18286 20242 18338
rect 21310 18286 21362 18338
rect 23438 18286 23490 18338
rect 24670 18286 24722 18338
rect 26462 18286 26514 18338
rect 26574 18286 26626 18338
rect 30158 18286 30210 18338
rect 30606 18286 30658 18338
rect 36094 18286 36146 18338
rect 42142 18286 42194 18338
rect 42478 18286 42530 18338
rect 43262 18286 43314 18338
rect 45390 18286 45442 18338
rect 4510 18174 4562 18226
rect 9998 18174 10050 18226
rect 10670 18174 10722 18226
rect 18622 18174 18674 18226
rect 20078 18174 20130 18226
rect 25230 18174 25282 18226
rect 25678 18174 25730 18226
rect 36542 18174 36594 18226
rect 37102 18174 37154 18226
rect 47070 18174 47122 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 19070 17838 19122 17890
rect 33182 17838 33234 17890
rect 44942 17838 44994 17890
rect 4622 17726 4674 17778
rect 8654 17726 8706 17778
rect 10782 17726 10834 17778
rect 13694 17726 13746 17778
rect 19406 17726 19458 17778
rect 19630 17726 19682 17778
rect 21422 17726 21474 17778
rect 22206 17726 22258 17778
rect 26910 17726 26962 17778
rect 27694 17726 27746 17778
rect 28366 17726 28418 17778
rect 29262 17726 29314 17778
rect 30718 17726 30770 17778
rect 32846 17726 32898 17778
rect 33966 17726 34018 17778
rect 37102 17726 37154 17778
rect 40350 17726 40402 17778
rect 42478 17726 42530 17778
rect 42926 17726 42978 17778
rect 43374 17726 43426 17778
rect 43822 17726 43874 17778
rect 44830 17726 44882 17778
rect 49198 17726 49250 17778
rect 1822 17614 1874 17666
rect 6302 17614 6354 17666
rect 7982 17614 8034 17666
rect 12686 17614 12738 17666
rect 18398 17614 18450 17666
rect 20190 17614 20242 17666
rect 20414 17614 20466 17666
rect 20862 17614 20914 17666
rect 22094 17614 22146 17666
rect 22318 17614 22370 17666
rect 22654 17614 22706 17666
rect 22878 17614 22930 17666
rect 23214 17614 23266 17666
rect 24110 17614 24162 17666
rect 24782 17614 24834 17666
rect 27582 17614 27634 17666
rect 28030 17614 28082 17666
rect 30046 17614 30098 17666
rect 33518 17614 33570 17666
rect 33854 17614 33906 17666
rect 34078 17614 34130 17666
rect 34526 17614 34578 17666
rect 37326 17614 37378 17666
rect 37550 17614 37602 17666
rect 38334 17614 38386 17666
rect 38446 17614 38498 17666
rect 38894 17614 38946 17666
rect 39006 17614 39058 17666
rect 39566 17614 39618 17666
rect 44158 17614 44210 17666
rect 45502 17614 45554 17666
rect 45726 17614 45778 17666
rect 46286 17614 46338 17666
rect 2494 17502 2546 17554
rect 6862 17502 6914 17554
rect 7198 17502 7250 17554
rect 7534 17502 7586 17554
rect 11118 17502 11170 17554
rect 11902 17502 11954 17554
rect 21310 17502 21362 17554
rect 23438 17502 23490 17554
rect 27358 17502 27410 17554
rect 28478 17502 28530 17554
rect 33294 17502 33346 17554
rect 34302 17502 34354 17554
rect 35422 17502 35474 17554
rect 36094 17502 36146 17554
rect 45278 17502 45330 17554
rect 47070 17502 47122 17554
rect 5966 17390 6018 17442
rect 6526 17390 6578 17442
rect 6750 17390 6802 17442
rect 11230 17390 11282 17442
rect 11454 17390 11506 17442
rect 11566 17390 11618 17442
rect 11790 17390 11842 17442
rect 12910 17390 12962 17442
rect 20302 17390 20354 17442
rect 21534 17390 21586 17442
rect 21758 17390 21810 17442
rect 22990 17390 23042 17442
rect 27806 17390 27858 17442
rect 35086 17390 35138 17442
rect 35758 17390 35810 17442
rect 39118 17390 39170 17442
rect 45614 17390 45666 17442
rect 45838 17390 45890 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 9662 17054 9714 17106
rect 16718 17054 16770 17106
rect 17838 17054 17890 17106
rect 21422 17054 21474 17106
rect 22318 17054 22370 17106
rect 23438 17054 23490 17106
rect 23886 17054 23938 17106
rect 24334 17054 24386 17106
rect 24782 17054 24834 17106
rect 25454 17054 25506 17106
rect 26238 17054 26290 17106
rect 31726 17054 31778 17106
rect 31838 17054 31890 17106
rect 33406 17054 33458 17106
rect 35534 17054 35586 17106
rect 47966 17054 48018 17106
rect 48862 17054 48914 17106
rect 1710 16942 1762 16994
rect 2270 16942 2322 16994
rect 2830 16942 2882 16994
rect 9550 16942 9602 16994
rect 14142 16942 14194 16994
rect 17726 16942 17778 16994
rect 20302 16942 20354 16994
rect 21870 16942 21922 16994
rect 27694 16942 27746 16994
rect 30270 16942 30322 16994
rect 30942 16942 30994 16994
rect 33518 16942 33570 16994
rect 33966 16942 34018 16994
rect 34078 16942 34130 16994
rect 34526 16942 34578 16994
rect 34638 16942 34690 16994
rect 35086 16942 35138 16994
rect 35758 16942 35810 16994
rect 40910 16942 40962 16994
rect 42142 16942 42194 16994
rect 45390 16942 45442 16994
rect 49086 16942 49138 16994
rect 1934 16830 1986 16882
rect 7870 16830 7922 16882
rect 8094 16830 8146 16882
rect 8542 16830 8594 16882
rect 8654 16830 8706 16882
rect 9886 16830 9938 16882
rect 12238 16830 12290 16882
rect 13022 16830 13074 16882
rect 13358 16830 13410 16882
rect 16830 16830 16882 16882
rect 21086 16830 21138 16882
rect 21646 16830 21698 16882
rect 22542 16830 22594 16882
rect 26574 16830 26626 16882
rect 27022 16830 27074 16882
rect 31502 16830 31554 16882
rect 31614 16830 31666 16882
rect 32062 16830 32114 16882
rect 36542 16830 36594 16882
rect 36654 16830 36706 16882
rect 36990 16830 37042 16882
rect 40350 16830 40402 16882
rect 41022 16830 41074 16882
rect 41470 16830 41522 16882
rect 44718 16830 44770 16882
rect 2158 16718 2210 16770
rect 8318 16718 8370 16770
rect 10110 16718 10162 16770
rect 16270 16718 16322 16770
rect 18174 16718 18226 16770
rect 21534 16718 21586 16770
rect 29822 16718 29874 16770
rect 30158 16718 30210 16770
rect 32398 16718 32450 16770
rect 37438 16718 37490 16770
rect 39566 16718 39618 16770
rect 44270 16718 44322 16770
rect 47518 16718 47570 16770
rect 47854 16718 47906 16770
rect 48750 16718 48802 16770
rect 30830 16606 30882 16658
rect 32510 16606 32562 16658
rect 33406 16606 33458 16658
rect 33966 16606 34018 16658
rect 34526 16606 34578 16658
rect 34974 16606 35026 16658
rect 48190 16606 48242 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 9550 16270 9602 16322
rect 9998 16270 10050 16322
rect 37550 16270 37602 16322
rect 48190 16270 48242 16322
rect 4622 16158 4674 16210
rect 5966 16158 6018 16210
rect 8094 16158 8146 16210
rect 11678 16158 11730 16210
rect 17166 16158 17218 16210
rect 17838 16158 17890 16210
rect 19966 16158 20018 16210
rect 21758 16158 21810 16210
rect 23550 16158 23602 16210
rect 24670 16158 24722 16210
rect 26798 16158 26850 16210
rect 27358 16158 27410 16210
rect 28366 16158 28418 16210
rect 29150 16158 29202 16210
rect 30158 16158 30210 16210
rect 30606 16158 30658 16210
rect 37214 16158 37266 16210
rect 42366 16158 42418 16210
rect 44270 16158 44322 16210
rect 45950 16158 46002 16210
rect 48414 16158 48466 16210
rect 1822 16046 1874 16098
rect 8878 16046 8930 16098
rect 9326 16046 9378 16098
rect 9774 16046 9826 16098
rect 10670 16046 10722 16098
rect 10894 16046 10946 16098
rect 11230 16046 11282 16098
rect 11566 16046 11618 16098
rect 11790 16046 11842 16098
rect 13358 16046 13410 16098
rect 13694 16046 13746 16098
rect 16830 16046 16882 16098
rect 17278 16046 17330 16098
rect 17390 16046 17442 16098
rect 20750 16046 20802 16098
rect 21310 16046 21362 16098
rect 21534 16046 21586 16098
rect 23102 16046 23154 16098
rect 23998 16046 24050 16098
rect 27470 16046 27522 16098
rect 28030 16046 28082 16098
rect 28254 16046 28306 16098
rect 35310 16046 35362 16098
rect 37326 16046 37378 16098
rect 37550 16046 37602 16098
rect 38894 16046 38946 16098
rect 39454 16046 39506 16098
rect 42702 16046 42754 16098
rect 46286 16046 46338 16098
rect 47070 16046 47122 16098
rect 47294 16046 47346 16098
rect 48862 16046 48914 16098
rect 2494 15934 2546 15986
rect 10110 15934 10162 15986
rect 10446 15934 10498 15986
rect 12126 15934 12178 15986
rect 12686 15934 12738 15986
rect 12798 15934 12850 15986
rect 13022 15934 13074 15986
rect 14030 15934 14082 15986
rect 15486 15934 15538 15986
rect 15822 15934 15874 15986
rect 16158 15934 16210 15986
rect 21758 15934 21810 15986
rect 22542 15934 22594 15986
rect 27246 15934 27298 15986
rect 27694 15934 27746 15986
rect 28478 15934 28530 15986
rect 33518 15934 33570 15986
rect 38558 15934 38610 15986
rect 39118 15934 39170 15986
rect 40238 15934 40290 15986
rect 42926 15934 42978 15986
rect 43598 15934 43650 15986
rect 46846 15934 46898 15986
rect 48638 15934 48690 15986
rect 10558 15822 10610 15874
rect 13582 15822 13634 15874
rect 14478 15822 14530 15874
rect 14814 15822 14866 15874
rect 15150 15822 15202 15874
rect 17054 15822 17106 15874
rect 22206 15822 22258 15874
rect 29262 15822 29314 15874
rect 38670 15822 38722 15874
rect 42814 15822 42866 15874
rect 45054 15822 45106 15874
rect 48750 15822 48802 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 2046 15486 2098 15538
rect 2270 15486 2322 15538
rect 3390 15486 3442 15538
rect 5630 15486 5682 15538
rect 7758 15486 7810 15538
rect 8654 15486 8706 15538
rect 16718 15486 16770 15538
rect 17614 15486 17666 15538
rect 19406 15486 19458 15538
rect 20078 15486 20130 15538
rect 20526 15486 20578 15538
rect 20862 15486 20914 15538
rect 21198 15486 21250 15538
rect 24558 15486 24610 15538
rect 25790 15486 25842 15538
rect 26126 15486 26178 15538
rect 26462 15486 26514 15538
rect 26686 15486 26738 15538
rect 37886 15486 37938 15538
rect 38670 15486 38722 15538
rect 38894 15486 38946 15538
rect 41470 15486 41522 15538
rect 2382 15374 2434 15426
rect 2830 15374 2882 15426
rect 4286 15374 4338 15426
rect 5742 15374 5794 15426
rect 6190 15374 6242 15426
rect 6974 15374 7026 15426
rect 7086 15374 7138 15426
rect 8094 15374 8146 15426
rect 8430 15374 8482 15426
rect 8766 15374 8818 15426
rect 8990 15374 9042 15426
rect 16606 15374 16658 15426
rect 28254 15374 28306 15426
rect 29598 15374 29650 15426
rect 30606 15374 30658 15426
rect 32286 15374 32338 15426
rect 32398 15374 32450 15426
rect 33182 15374 33234 15426
rect 38558 15374 38610 15426
rect 39230 15374 39282 15426
rect 39342 15374 39394 15426
rect 39678 15374 39730 15426
rect 39902 15374 39954 15426
rect 41134 15374 41186 15426
rect 41918 15374 41970 15426
rect 48862 15374 48914 15426
rect 2606 15262 2658 15314
rect 2942 15262 2994 15314
rect 3278 15262 3330 15314
rect 3614 15262 3666 15314
rect 3838 15262 3890 15314
rect 4174 15262 4226 15314
rect 5854 15262 5906 15314
rect 6526 15262 6578 15314
rect 6750 15262 6802 15314
rect 15038 15262 15090 15314
rect 15486 15262 15538 15314
rect 15710 15262 15762 15314
rect 16046 15262 16098 15314
rect 18062 15262 18114 15314
rect 18398 15262 18450 15314
rect 18846 15262 18898 15314
rect 21646 15262 21698 15314
rect 22318 15262 22370 15314
rect 27134 15262 27186 15314
rect 27582 15262 27634 15314
rect 29038 15262 29090 15314
rect 30830 15262 30882 15314
rect 32622 15262 32674 15314
rect 33518 15262 33570 15314
rect 37550 15262 37602 15314
rect 37774 15262 37826 15314
rect 42030 15262 42082 15314
rect 42142 15262 42194 15314
rect 43038 15262 43090 15314
rect 49086 15262 49138 15314
rect 10110 15150 10162 15202
rect 15822 15150 15874 15202
rect 26574 15150 26626 15202
rect 31838 15150 31890 15202
rect 33070 15150 33122 15202
rect 34302 15150 34354 15202
rect 36430 15150 36482 15202
rect 37214 15150 37266 15202
rect 40014 15150 40066 15202
rect 46062 15150 46114 15202
rect 17390 15038 17442 15090
rect 18174 15038 18226 15090
rect 31950 15038 32002 15090
rect 39230 15038 39282 15090
rect 42590 15038 42642 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 8654 14702 8706 14754
rect 4622 14590 4674 14642
rect 9214 14590 9266 14642
rect 12910 14590 12962 14642
rect 13582 14590 13634 14642
rect 14702 14590 14754 14642
rect 16830 14590 16882 14642
rect 17278 14590 17330 14642
rect 17950 14590 18002 14642
rect 26910 14590 26962 14642
rect 27918 14590 27970 14642
rect 30046 14590 30098 14642
rect 32174 14590 32226 14642
rect 35534 14590 35586 14642
rect 36094 14590 36146 14642
rect 36430 14590 36482 14642
rect 37438 14590 37490 14642
rect 38110 14590 38162 14642
rect 40798 14590 40850 14642
rect 41358 14590 41410 14642
rect 44942 14590 44994 14642
rect 45502 14590 45554 14642
rect 49198 14590 49250 14642
rect 1822 14478 1874 14530
rect 6862 14478 6914 14530
rect 8318 14478 8370 14530
rect 9438 14478 9490 14530
rect 10110 14478 10162 14530
rect 13918 14478 13970 14530
rect 19854 14478 19906 14530
rect 20078 14478 20130 14530
rect 20414 14478 20466 14530
rect 25566 14478 25618 14530
rect 28030 14478 28082 14530
rect 28366 14478 28418 14530
rect 29374 14478 29426 14530
rect 32734 14478 32786 14530
rect 37550 14478 37602 14530
rect 37998 14478 38050 14530
rect 38222 14478 38274 14530
rect 38558 14478 38610 14530
rect 39006 14478 39058 14530
rect 39118 14478 39170 14530
rect 39566 14478 39618 14530
rect 44270 14478 44322 14530
rect 45390 14478 45442 14530
rect 45726 14478 45778 14530
rect 45950 14478 46002 14530
rect 46286 14478 46338 14530
rect 2494 14366 2546 14418
rect 7086 14366 7138 14418
rect 7198 14366 7250 14418
rect 9550 14366 9602 14418
rect 10782 14366 10834 14418
rect 23662 14366 23714 14418
rect 27806 14366 27858 14418
rect 33406 14366 33458 14418
rect 37438 14366 37490 14418
rect 38894 14366 38946 14418
rect 43486 14366 43538 14418
rect 47070 14366 47122 14418
rect 5630 14254 5682 14306
rect 5966 14254 6018 14306
rect 6302 14254 6354 14306
rect 6638 14254 6690 14306
rect 8094 14254 8146 14306
rect 8542 14254 8594 14306
rect 9774 14254 9826 14306
rect 18174 14254 18226 14306
rect 18510 14254 18562 14306
rect 19294 14254 19346 14306
rect 19518 14254 19570 14306
rect 20750 14254 20802 14306
rect 27470 14254 27522 14306
rect 39790 14254 39842 14306
rect 39902 14254 39954 14306
rect 40014 14254 40066 14306
rect 40238 14254 40290 14306
rect 45054 14254 45106 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 3502 13918 3554 13970
rect 6190 13918 6242 13970
rect 6414 13918 6466 13970
rect 7310 13918 7362 13970
rect 8206 13918 8258 13970
rect 9774 13918 9826 13970
rect 9998 13918 10050 13970
rect 10782 13918 10834 13970
rect 11902 13918 11954 13970
rect 12574 13918 12626 13970
rect 12798 13918 12850 13970
rect 16830 13918 16882 13970
rect 23998 13918 24050 13970
rect 24334 13918 24386 13970
rect 26686 13918 26738 13970
rect 27246 13918 27298 13970
rect 33518 13918 33570 13970
rect 34638 13918 34690 13970
rect 34862 13918 34914 13970
rect 35534 13918 35586 13970
rect 41022 13918 41074 13970
rect 41246 13918 41298 13970
rect 41470 13918 41522 13970
rect 42814 13918 42866 13970
rect 46622 13918 46674 13970
rect 48302 13918 48354 13970
rect 3166 13806 3218 13858
rect 3278 13806 3330 13858
rect 3838 13806 3890 13858
rect 4062 13806 4114 13858
rect 4398 13806 4450 13858
rect 4846 13806 4898 13858
rect 5518 13806 5570 13858
rect 5630 13806 5682 13858
rect 6638 13806 6690 13858
rect 8318 13806 8370 13858
rect 10334 13806 10386 13858
rect 11566 13806 11618 13858
rect 12462 13806 12514 13858
rect 13918 13806 13970 13858
rect 18622 13806 18674 13858
rect 24670 13806 24722 13858
rect 33742 13806 33794 13858
rect 39342 13806 39394 13858
rect 39678 13806 39730 13858
rect 40014 13806 40066 13858
rect 46958 13806 47010 13858
rect 47742 13806 47794 13858
rect 48862 13806 48914 13858
rect 48974 13806 49026 13858
rect 3726 13694 3778 13746
rect 4174 13694 4226 13746
rect 4510 13694 4562 13746
rect 5854 13694 5906 13746
rect 6078 13694 6130 13746
rect 6974 13694 7026 13746
rect 7646 13694 7698 13746
rect 7982 13694 8034 13746
rect 8654 13694 8706 13746
rect 10558 13694 10610 13746
rect 10894 13694 10946 13746
rect 11118 13694 11170 13746
rect 13246 13694 13298 13746
rect 17278 13694 17330 13746
rect 17614 13694 17666 13746
rect 17950 13694 18002 13746
rect 19518 13694 19570 13746
rect 19742 13694 19794 13746
rect 20078 13694 20130 13746
rect 20414 13694 20466 13746
rect 23774 13694 23826 13746
rect 27022 13694 27074 13746
rect 28814 13694 28866 13746
rect 29262 13694 29314 13746
rect 32510 13694 32562 13746
rect 33070 13694 33122 13746
rect 33294 13694 33346 13746
rect 34190 13694 34242 13746
rect 34414 13694 34466 13746
rect 35758 13694 35810 13746
rect 39118 13694 39170 13746
rect 40238 13694 40290 13746
rect 41358 13694 41410 13746
rect 41694 13694 41746 13746
rect 42142 13694 42194 13746
rect 42254 13694 42306 13746
rect 43486 13694 43538 13746
rect 47518 13694 47570 13746
rect 48078 13694 48130 13746
rect 48750 13694 48802 13746
rect 8878 13582 8930 13634
rect 16046 13582 16098 13634
rect 17502 13582 17554 13634
rect 19630 13582 19682 13634
rect 21198 13582 21250 13634
rect 23326 13582 23378 13634
rect 26014 13582 26066 13634
rect 28030 13582 28082 13634
rect 28366 13582 28418 13634
rect 29934 13582 29986 13634
rect 32062 13582 32114 13634
rect 33630 13582 33682 13634
rect 34750 13582 34802 13634
rect 36542 13582 36594 13634
rect 38670 13582 38722 13634
rect 39790 13582 39842 13634
rect 41918 13582 41970 13634
rect 44158 13582 44210 13634
rect 46286 13582 46338 13634
rect 47294 13582 47346 13634
rect 8990 13470 9042 13522
rect 18510 13470 18562 13522
rect 18846 13470 18898 13522
rect 25454 13470 25506 13522
rect 25790 13470 25842 13522
rect 27918 13470 27970 13522
rect 28366 13470 28418 13522
rect 42702 13470 42754 13522
rect 43038 13470 43090 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 11342 13134 11394 13186
rect 21646 13134 21698 13186
rect 32846 13134 32898 13186
rect 45054 13134 45106 13186
rect 45838 13134 45890 13186
rect 2494 13022 2546 13074
rect 4622 13022 4674 13074
rect 7646 13022 7698 13074
rect 9774 13022 9826 13074
rect 11118 13022 11170 13074
rect 11902 13022 11954 13074
rect 14030 13022 14082 13074
rect 17278 13022 17330 13074
rect 18510 13022 18562 13074
rect 20638 13022 20690 13074
rect 24446 13022 24498 13074
rect 26574 13022 26626 13074
rect 27246 13022 27298 13074
rect 30270 13022 30322 13074
rect 33406 13022 33458 13074
rect 36094 13022 36146 13074
rect 36430 13022 36482 13074
rect 39454 13022 39506 13074
rect 41582 13022 41634 13074
rect 42030 13022 42082 13074
rect 43150 13022 43202 13074
rect 45390 13022 45442 13074
rect 1822 12910 1874 12962
rect 5630 12910 5682 12962
rect 5854 12910 5906 12962
rect 6190 12910 6242 12962
rect 6414 12910 6466 12962
rect 7086 12910 7138 12962
rect 10558 12910 10610 12962
rect 11678 12910 11730 12962
rect 12126 12910 12178 12962
rect 12462 12910 12514 12962
rect 12798 12910 12850 12962
rect 13806 12910 13858 12962
rect 14366 12910 14418 12962
rect 17726 12910 17778 12962
rect 21646 12910 21698 12962
rect 22990 12910 23042 12962
rect 23662 12910 23714 12962
rect 27694 12910 27746 12962
rect 28590 12910 28642 12962
rect 29486 12910 29538 12962
rect 29710 12910 29762 12962
rect 29934 12910 29986 12962
rect 30382 12910 30434 12962
rect 31502 12910 31554 12962
rect 32062 12910 32114 12962
rect 33070 12910 33122 12962
rect 33294 12910 33346 12962
rect 33518 12910 33570 12962
rect 34302 12910 34354 12962
rect 34862 12910 34914 12962
rect 36318 12910 36370 12962
rect 37214 12910 37266 12962
rect 37662 12910 37714 12962
rect 38670 12910 38722 12962
rect 42366 12910 42418 12962
rect 42814 12910 42866 12962
rect 43822 12910 43874 12962
rect 44046 12910 44098 12962
rect 46062 12910 46114 12962
rect 46286 12910 46338 12962
rect 47294 12910 47346 12962
rect 47518 12910 47570 12962
rect 48078 12910 48130 12962
rect 48302 12910 48354 12962
rect 49198 12910 49250 12962
rect 6750 12798 6802 12850
rect 7198 12798 7250 12850
rect 12350 12798 12402 12850
rect 12910 12798 12962 12850
rect 15150 12798 15202 12850
rect 21982 12798 22034 12850
rect 22542 12798 22594 12850
rect 22878 12798 22930 12850
rect 27918 12798 27970 12850
rect 30718 12798 30770 12850
rect 31390 12798 31442 12850
rect 34974 12798 35026 12850
rect 35310 12798 35362 12850
rect 35422 12798 35474 12850
rect 36990 12798 37042 12850
rect 46622 12798 46674 12850
rect 48190 12798 48242 12850
rect 49086 12798 49138 12850
rect 5182 12686 5234 12738
rect 5966 12686 6018 12738
rect 6638 12686 6690 12738
rect 7422 12686 7474 12738
rect 13470 12686 13522 12738
rect 22766 12686 22818 12738
rect 23214 12686 23266 12738
rect 28478 12686 28530 12738
rect 29262 12686 29314 12738
rect 29374 12686 29426 12738
rect 35646 12686 35698 12738
rect 37326 12686 37378 12738
rect 37886 12686 37938 12738
rect 38222 12686 38274 12738
rect 45166 12686 45218 12738
rect 46174 12686 46226 12738
rect 48750 12686 48802 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 3502 12350 3554 12402
rect 9550 12350 9602 12402
rect 9662 12350 9714 12402
rect 9774 12350 9826 12402
rect 15822 12350 15874 12402
rect 15934 12350 15986 12402
rect 21086 12350 21138 12402
rect 22430 12350 22482 12402
rect 22766 12350 22818 12402
rect 24446 12350 24498 12402
rect 25454 12350 25506 12402
rect 25678 12350 25730 12402
rect 31838 12350 31890 12402
rect 40014 12350 40066 12402
rect 46510 12350 46562 12402
rect 3390 12238 3442 12290
rect 3726 12238 3778 12290
rect 4510 12238 4562 12290
rect 5630 12238 5682 12290
rect 17950 12238 18002 12290
rect 18062 12238 18114 12290
rect 21422 12238 21474 12290
rect 21758 12238 21810 12290
rect 22094 12238 22146 12290
rect 30158 12238 30210 12290
rect 31054 12238 31106 12290
rect 32398 12238 32450 12290
rect 32510 12238 32562 12290
rect 35758 12238 35810 12290
rect 42814 12238 42866 12290
rect 45278 12238 45330 12290
rect 45838 12238 45890 12290
rect 46734 12238 46786 12290
rect 3838 12126 3890 12178
rect 4286 12126 4338 12178
rect 4846 12126 4898 12178
rect 5070 12126 5122 12178
rect 8766 12126 8818 12178
rect 10222 12126 10274 12178
rect 10782 12126 10834 12178
rect 14478 12126 14530 12178
rect 14814 12126 14866 12178
rect 15038 12126 15090 12178
rect 15374 12126 15426 12178
rect 15710 12126 15762 12178
rect 16382 12126 16434 12178
rect 16606 12126 16658 12178
rect 16718 12126 16770 12178
rect 17390 12126 17442 12178
rect 17838 12126 17890 12178
rect 19070 12126 19122 12178
rect 19742 12126 19794 12178
rect 23102 12126 23154 12178
rect 23326 12126 23378 12178
rect 26126 12126 26178 12178
rect 26462 12126 26514 12178
rect 29710 12126 29762 12178
rect 31166 12126 31218 12178
rect 31614 12126 31666 12178
rect 37102 12126 37154 12178
rect 38782 12126 38834 12178
rect 39230 12126 39282 12178
rect 39566 12126 39618 12178
rect 39790 12126 39842 12178
rect 41246 12126 41298 12178
rect 41470 12126 41522 12178
rect 41694 12126 41746 12178
rect 41918 12126 41970 12178
rect 42478 12126 42530 12178
rect 42702 12126 42754 12178
rect 43262 12126 43314 12178
rect 43486 12126 43538 12178
rect 44942 12126 44994 12178
rect 46062 12126 46114 12178
rect 47742 12126 47794 12178
rect 49086 12126 49138 12178
rect 4062 12014 4114 12066
rect 5966 12014 6018 12066
rect 8094 12014 8146 12066
rect 11566 12014 11618 12066
rect 13694 12014 13746 12066
rect 14142 12014 14194 12066
rect 14590 12014 14642 12066
rect 18846 12014 18898 12066
rect 20302 12014 20354 12066
rect 23998 12014 24050 12066
rect 24446 12014 24498 12066
rect 24670 12014 24722 12066
rect 25566 12014 25618 12066
rect 26798 12014 26850 12066
rect 28926 12014 28978 12066
rect 31278 12014 31330 12066
rect 39678 12014 39730 12066
rect 41022 12014 41074 12066
rect 44046 12014 44098 12066
rect 45950 12014 46002 12066
rect 47518 12014 47570 12066
rect 5294 11902 5346 11954
rect 5518 11902 5570 11954
rect 16270 11902 16322 11954
rect 19070 11902 19122 11954
rect 19406 11902 19458 11954
rect 20078 11902 20130 11954
rect 30270 11902 30322 11954
rect 42366 11902 42418 11954
rect 43150 11902 43202 11954
rect 43598 11902 43650 11954
rect 44270 11902 44322 11954
rect 44606 11902 44658 11954
rect 46398 11902 46450 11954
rect 47966 11902 48018 11954
rect 48750 11902 48802 11954
rect 49086 11902 49138 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 11342 11566 11394 11618
rect 12350 11566 12402 11618
rect 44270 11566 44322 11618
rect 49086 11566 49138 11618
rect 2494 11454 2546 11506
rect 4622 11454 4674 11506
rect 8766 11454 8818 11506
rect 11342 11454 11394 11506
rect 11790 11454 11842 11506
rect 12238 11454 12290 11506
rect 19182 11454 19234 11506
rect 19854 11454 19906 11506
rect 22430 11454 22482 11506
rect 23326 11454 23378 11506
rect 24446 11454 24498 11506
rect 26574 11454 26626 11506
rect 30942 11454 30994 11506
rect 33070 11454 33122 11506
rect 33518 11454 33570 11506
rect 35646 11454 35698 11506
rect 45614 11454 45666 11506
rect 47742 11454 47794 11506
rect 48190 11454 48242 11506
rect 1822 11342 1874 11394
rect 10782 11342 10834 11394
rect 12910 11342 12962 11394
rect 18286 11342 18338 11394
rect 19966 11342 20018 11394
rect 20414 11342 20466 11394
rect 23662 11342 23714 11394
rect 26910 11342 26962 11394
rect 28366 11342 28418 11394
rect 28590 11342 28642 11394
rect 29150 11342 29202 11394
rect 29598 11342 29650 11394
rect 30270 11342 30322 11394
rect 36430 11342 36482 11394
rect 36990 11342 37042 11394
rect 37550 11342 37602 11394
rect 42926 11342 42978 11394
rect 43486 11342 43538 11394
rect 44830 11342 44882 11394
rect 47966 11342 48018 11394
rect 48302 11342 48354 11394
rect 48638 11342 48690 11394
rect 48974 11342 49026 11394
rect 12574 11230 12626 11282
rect 13694 11230 13746 11282
rect 20862 11230 20914 11282
rect 21646 11230 21698 11282
rect 38110 11230 38162 11282
rect 43710 11230 43762 11282
rect 43822 11230 43874 11282
rect 5070 11118 5122 11170
rect 19742 11118 19794 11170
rect 21982 11118 22034 11170
rect 22990 11118 23042 11170
rect 27246 11118 27298 11170
rect 27358 11118 27410 11170
rect 27470 11118 27522 11170
rect 28030 11118 28082 11170
rect 49086 11118 49138 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 5518 10782 5570 10834
rect 5742 10782 5794 10834
rect 6638 10782 6690 10834
rect 9102 10782 9154 10834
rect 10222 10782 10274 10834
rect 16718 10782 16770 10834
rect 16830 10782 16882 10834
rect 20974 10782 21026 10834
rect 31614 10782 31666 10834
rect 31726 10782 31778 10834
rect 31838 10782 31890 10834
rect 32398 10782 32450 10834
rect 37102 10782 37154 10834
rect 42366 10782 42418 10834
rect 45838 10782 45890 10834
rect 5854 10670 5906 10722
rect 6862 10670 6914 10722
rect 7422 10670 7474 10722
rect 10894 10670 10946 10722
rect 11790 10670 11842 10722
rect 13806 10670 13858 10722
rect 18398 10670 18450 10722
rect 28814 10670 28866 10722
rect 32510 10670 32562 10722
rect 34078 10670 34130 10722
rect 34974 10670 35026 10722
rect 35198 10670 35250 10722
rect 36654 10670 36706 10722
rect 41246 10670 41298 10722
rect 44718 10670 44770 10722
rect 46734 10670 46786 10722
rect 47294 10670 47346 10722
rect 48750 10670 48802 10722
rect 48974 10670 49026 10722
rect 6526 10558 6578 10610
rect 6974 10558 7026 10610
rect 7646 10558 7698 10610
rect 10558 10558 10610 10610
rect 11230 10558 11282 10610
rect 13022 10558 13074 10610
rect 16158 10558 16210 10610
rect 16606 10558 16658 10610
rect 17726 10558 17778 10610
rect 21310 10558 21362 10610
rect 25342 10558 25394 10610
rect 29374 10558 29426 10610
rect 30046 10558 30098 10610
rect 31166 10558 31218 10610
rect 31390 10558 31442 10610
rect 32174 10558 32226 10610
rect 33070 10558 33122 10610
rect 33518 10558 33570 10610
rect 34414 10558 34466 10610
rect 34526 10558 34578 10610
rect 35422 10558 35474 10610
rect 35646 10558 35698 10610
rect 36094 10558 36146 10610
rect 36318 10558 36370 10610
rect 37550 10558 37602 10610
rect 41918 10558 41970 10610
rect 45502 10558 45554 10610
rect 46062 10558 46114 10610
rect 48078 10558 48130 10610
rect 5294 10446 5346 10498
rect 7198 10446 7250 10498
rect 7982 10446 8034 10498
rect 9886 10446 9938 10498
rect 12798 10446 12850 10498
rect 15934 10446 15986 10498
rect 20526 10446 20578 10498
rect 22094 10446 22146 10498
rect 24222 10446 24274 10498
rect 24670 10446 24722 10498
rect 26014 10446 26066 10498
rect 28142 10446 28194 10498
rect 30718 10446 30770 10498
rect 34190 10446 34242 10498
rect 35758 10446 35810 10498
rect 36542 10446 36594 10498
rect 38222 10446 38274 10498
rect 40350 10446 40402 10498
rect 42590 10446 42642 10498
rect 47630 10446 47682 10498
rect 48862 10446 48914 10498
rect 8206 10334 8258 10386
rect 8542 10334 8594 10386
rect 11566 10334 11618 10386
rect 11902 10334 11954 10386
rect 41470 10334 41522 10386
rect 41694 10334 41746 10386
rect 46510 10334 46562 10386
rect 46846 10334 46898 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 11902 9998 11954 10050
rect 20302 9998 20354 10050
rect 25790 9998 25842 10050
rect 26462 9998 26514 10050
rect 45390 9998 45442 10050
rect 5854 9886 5906 9938
rect 9438 9886 9490 9938
rect 11566 9886 11618 9938
rect 12462 9886 12514 9938
rect 15262 9886 15314 9938
rect 19742 9886 19794 9938
rect 20078 9886 20130 9938
rect 21758 9886 21810 9938
rect 25678 9886 25730 9938
rect 26686 9886 26738 9938
rect 35646 9886 35698 9938
rect 37550 9886 37602 9938
rect 41134 9886 41186 9938
rect 44830 9886 44882 9938
rect 47070 9886 47122 9938
rect 49198 9886 49250 9938
rect 4734 9774 4786 9826
rect 7310 9774 7362 9826
rect 7758 9774 7810 9826
rect 7870 9774 7922 9826
rect 8318 9774 8370 9826
rect 8766 9774 8818 9826
rect 12238 9774 12290 9826
rect 12910 9774 12962 9826
rect 13694 9774 13746 9826
rect 15598 9774 15650 9826
rect 15710 9774 15762 9826
rect 15822 9774 15874 9826
rect 16830 9774 16882 9826
rect 21646 9774 21698 9826
rect 21982 9774 22034 9826
rect 22878 9774 22930 9826
rect 23550 9774 23602 9826
rect 23774 9774 23826 9826
rect 27134 9774 27186 9826
rect 27806 9774 27858 9826
rect 28142 9774 28194 9826
rect 29374 9774 29426 9826
rect 30942 9774 30994 9826
rect 31278 9774 31330 9826
rect 32846 9774 32898 9826
rect 36430 9774 36482 9826
rect 37102 9774 37154 9826
rect 38222 9774 38274 9826
rect 41470 9774 41522 9826
rect 45054 9774 45106 9826
rect 46286 9774 46338 9826
rect 5182 9662 5234 9714
rect 17614 9662 17666 9714
rect 22766 9662 22818 9714
rect 23214 9662 23266 9714
rect 24446 9662 24498 9714
rect 25566 9662 25618 9714
rect 26126 9662 26178 9714
rect 27470 9662 27522 9714
rect 28590 9662 28642 9714
rect 29598 9662 29650 9714
rect 33518 9662 33570 9714
rect 36094 9662 36146 9714
rect 39006 9662 39058 9714
rect 6302 9550 6354 9602
rect 6638 9550 6690 9602
rect 7086 9550 7138 9602
rect 7198 9550 7250 9602
rect 7646 9550 7698 9602
rect 13918 9550 13970 9602
rect 14814 9550 14866 9602
rect 16270 9550 16322 9602
rect 20638 9550 20690 9602
rect 22430 9550 22482 9602
rect 22654 9550 22706 9602
rect 24222 9550 24274 9602
rect 24334 9550 24386 9602
rect 24782 9550 24834 9602
rect 30270 9550 30322 9602
rect 42478 9550 42530 9602
rect 45838 9550 45890 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 8542 9214 8594 9266
rect 8990 9214 9042 9266
rect 9998 9214 10050 9266
rect 10782 9214 10834 9266
rect 11566 9214 11618 9266
rect 11678 9214 11730 9266
rect 12238 9214 12290 9266
rect 14478 9214 14530 9266
rect 16046 9214 16098 9266
rect 18286 9214 18338 9266
rect 18846 9214 18898 9266
rect 19070 9214 19122 9266
rect 22318 9214 22370 9266
rect 23326 9214 23378 9266
rect 25342 9214 25394 9266
rect 25566 9214 25618 9266
rect 27134 9214 27186 9266
rect 28366 9214 28418 9266
rect 31502 9214 31554 9266
rect 39342 9214 39394 9266
rect 40462 9214 40514 9266
rect 41246 9214 41298 9266
rect 41806 9214 41858 9266
rect 42030 9214 42082 9266
rect 46734 9214 46786 9266
rect 47742 9214 47794 9266
rect 5966 9102 6018 9154
rect 12910 9102 12962 9154
rect 13694 9102 13746 9154
rect 15262 9102 15314 9154
rect 16382 9102 16434 9154
rect 16718 9102 16770 9154
rect 20638 9102 20690 9154
rect 21422 9102 21474 9154
rect 25902 9102 25954 9154
rect 30158 9102 30210 9154
rect 31054 9102 31106 9154
rect 32510 9102 32562 9154
rect 33854 9102 33906 9154
rect 33966 9102 34018 9154
rect 36654 9102 36706 9154
rect 39566 9102 39618 9154
rect 45054 9102 45106 9154
rect 48750 9102 48802 9154
rect 5294 8990 5346 9042
rect 11006 8990 11058 9042
rect 11454 8990 11506 9042
rect 13134 8990 13186 9042
rect 13582 8990 13634 9042
rect 13918 8990 13970 9042
rect 15598 8990 15650 9042
rect 19518 8990 19570 9042
rect 20526 8990 20578 9042
rect 21646 8990 21698 9042
rect 22878 8990 22930 9042
rect 23550 8990 23602 9042
rect 23774 8990 23826 9042
rect 24110 8990 24162 9042
rect 24446 8990 24498 9042
rect 24558 8990 24610 9042
rect 24670 8990 24722 9042
rect 25230 8990 25282 9042
rect 25790 8990 25842 9042
rect 28926 8990 28978 9042
rect 29822 8990 29874 9042
rect 30046 8990 30098 9042
rect 30718 8990 30770 9042
rect 31614 8990 31666 9042
rect 32174 8990 32226 9042
rect 34190 8990 34242 9042
rect 37438 8990 37490 9042
rect 37886 8990 37938 9042
rect 38334 8990 38386 9042
rect 38782 8990 38834 9042
rect 39230 8990 39282 9042
rect 39678 8990 39730 9042
rect 41358 8990 41410 9042
rect 45838 8990 45890 9042
rect 46398 8990 46450 9042
rect 46622 8990 46674 9042
rect 46846 8990 46898 9042
rect 47070 8990 47122 9042
rect 47406 8990 47458 9042
rect 47630 8990 47682 9042
rect 47854 8990 47906 9042
rect 48078 8990 48130 9042
rect 49086 8990 49138 9042
rect 8094 8878 8146 8930
rect 10446 8878 10498 8930
rect 11006 8878 11058 8930
rect 12574 8878 12626 8930
rect 10222 8766 10274 8818
rect 15038 8878 15090 8930
rect 17502 8878 17554 8930
rect 18174 8878 18226 8930
rect 18958 8878 19010 8930
rect 20078 8878 20130 8930
rect 23662 8878 23714 8930
rect 26462 8878 26514 8930
rect 27918 8878 27970 8930
rect 28702 8878 28754 8930
rect 34526 8878 34578 8930
rect 41918 8878 41970 8930
rect 42590 8878 42642 8930
rect 42926 8878 42978 8930
rect 11902 8766 11954 8818
rect 12574 8766 12626 8818
rect 17390 8766 17442 8818
rect 18510 8766 18562 8818
rect 20190 8766 20242 8818
rect 20638 8766 20690 8818
rect 25902 8766 25954 8818
rect 26350 8766 26402 8818
rect 29150 8766 29202 8818
rect 29598 8766 29650 8818
rect 31502 8766 31554 8818
rect 32062 8766 32114 8818
rect 32398 8766 32450 8818
rect 33406 8766 33458 8818
rect 42366 8766 42418 8818
rect 42702 8766 42754 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 36990 8430 37042 8482
rect 8654 8318 8706 8370
rect 9550 8318 9602 8370
rect 11342 8318 11394 8370
rect 11678 8318 11730 8370
rect 13918 8318 13970 8370
rect 15486 8318 15538 8370
rect 16942 8318 16994 8370
rect 19070 8318 19122 8370
rect 20750 8318 20802 8370
rect 24110 8318 24162 8370
rect 26238 8318 26290 8370
rect 44270 8318 44322 8370
rect 47070 8318 47122 8370
rect 49198 8318 49250 8370
rect 7198 8206 7250 8258
rect 7646 8206 7698 8258
rect 7758 8206 7810 8258
rect 8206 8206 8258 8258
rect 8430 8206 8482 8258
rect 10222 8206 10274 8258
rect 10782 8206 10834 8258
rect 11118 8206 11170 8258
rect 12014 8206 12066 8258
rect 12350 8206 12402 8258
rect 12686 8206 12738 8258
rect 14142 8206 14194 8258
rect 16158 8206 16210 8258
rect 19406 8206 19458 8258
rect 19854 8206 19906 8258
rect 21422 8206 21474 8258
rect 21758 8206 21810 8258
rect 23102 8206 23154 8258
rect 23438 8206 23490 8258
rect 26798 8206 26850 8258
rect 28366 8206 28418 8258
rect 28590 8206 28642 8258
rect 29150 8206 29202 8258
rect 30942 8206 30994 8258
rect 32398 8206 32450 8258
rect 33742 8206 33794 8258
rect 34526 8206 34578 8258
rect 35870 8206 35922 8258
rect 37102 8206 37154 8258
rect 37550 8206 37602 8258
rect 37774 8206 37826 8258
rect 38782 8206 38834 8258
rect 41358 8206 41410 8258
rect 45502 8206 45554 8258
rect 45950 8206 46002 8258
rect 46286 8206 46338 8258
rect 6974 8094 7026 8146
rect 9886 8094 9938 8146
rect 10670 8094 10722 8146
rect 12238 8094 12290 8146
rect 13022 8094 13074 8146
rect 14814 8094 14866 8146
rect 15150 8094 15202 8146
rect 20526 8094 20578 8146
rect 21310 8094 21362 8146
rect 22766 8094 22818 8146
rect 26574 8094 26626 8146
rect 27694 8094 27746 8146
rect 28142 8094 28194 8146
rect 30158 8094 30210 8146
rect 33070 8094 33122 8146
rect 33182 8094 33234 8146
rect 34078 8094 34130 8146
rect 35086 8094 35138 8146
rect 36318 8094 36370 8146
rect 42142 8094 42194 8146
rect 45278 8094 45330 8146
rect 5070 7982 5122 8034
rect 6078 7982 6130 8034
rect 6638 7982 6690 8034
rect 7086 7982 7138 8034
rect 7534 7982 7586 8034
rect 8990 7982 9042 8034
rect 9662 7982 9714 8034
rect 10558 7982 10610 8034
rect 15374 7982 15426 8034
rect 20638 7982 20690 8034
rect 22878 7982 22930 8034
rect 27582 7982 27634 8034
rect 28478 7982 28530 8034
rect 29262 7982 29314 8034
rect 32622 7982 32674 8034
rect 32846 7982 32898 8034
rect 33966 7982 34018 8034
rect 34750 7982 34802 8034
rect 35422 7982 35474 8034
rect 35982 7982 36034 8034
rect 36094 7982 36146 8034
rect 36206 7982 36258 8034
rect 37886 7982 37938 8034
rect 39454 7982 39506 8034
rect 44942 7982 44994 8034
rect 45614 7982 45666 8034
rect 45726 7982 45778 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 13022 7646 13074 7698
rect 13246 7646 13298 7698
rect 24334 7646 24386 7698
rect 24446 7646 24498 7698
rect 30270 7646 30322 7698
rect 32286 7646 32338 7698
rect 38894 7646 38946 7698
rect 39566 7646 39618 7698
rect 42366 7646 42418 7698
rect 42478 7646 42530 7698
rect 48862 7646 48914 7698
rect 5294 7534 5346 7586
rect 7758 7534 7810 7586
rect 13470 7534 13522 7586
rect 16046 7534 16098 7586
rect 23214 7534 23266 7586
rect 23326 7534 23378 7586
rect 25230 7534 25282 7586
rect 30046 7534 30098 7586
rect 30494 7534 30546 7586
rect 32510 7534 32562 7586
rect 33182 7534 33234 7586
rect 33630 7534 33682 7586
rect 34078 7534 34130 7586
rect 34974 7534 35026 7586
rect 38558 7534 38610 7586
rect 40014 7534 40066 7586
rect 40910 7534 40962 7586
rect 48974 7534 49026 7586
rect 4622 7422 4674 7474
rect 7982 7422 8034 7474
rect 8318 7422 8370 7474
rect 8990 7422 9042 7474
rect 9774 7422 9826 7474
rect 16830 7422 16882 7474
rect 22654 7422 22706 7474
rect 22990 7422 23042 7474
rect 23774 7422 23826 7474
rect 25342 7422 25394 7474
rect 25566 7422 25618 7474
rect 27582 7422 27634 7474
rect 27806 7422 27858 7474
rect 28030 7422 28082 7474
rect 28478 7422 28530 7474
rect 30606 7422 30658 7474
rect 31054 7422 31106 7474
rect 31614 7422 31666 7474
rect 32958 7422 33010 7474
rect 33294 7422 33346 7474
rect 34750 7422 34802 7474
rect 38222 7422 38274 7474
rect 39230 7422 39282 7474
rect 39790 7422 39842 7474
rect 41246 7422 41298 7474
rect 41582 7422 41634 7474
rect 42030 7422 42082 7474
rect 42590 7422 42642 7474
rect 43038 7422 43090 7474
rect 7422 7310 7474 7362
rect 7870 7310 7922 7362
rect 10558 7310 10610 7362
rect 12686 7310 12738 7362
rect 13134 7310 13186 7362
rect 13918 7310 13970 7362
rect 17726 7310 17778 7362
rect 25678 7310 25730 7362
rect 30494 7310 30546 7362
rect 33966 7310 34018 7362
rect 35310 7310 35362 7362
rect 37438 7310 37490 7362
rect 39566 7310 39618 7362
rect 41134 7310 41186 7362
rect 41694 7310 41746 7362
rect 45726 7310 45778 7362
rect 23998 7198 24050 7250
rect 24558 7198 24610 7250
rect 26462 7198 26514 7250
rect 32174 7198 32226 7250
rect 34302 7198 34354 7250
rect 48750 7198 48802 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 7086 6862 7138 6914
rect 7422 6862 7474 6914
rect 8094 6862 8146 6914
rect 30606 6862 30658 6914
rect 30830 6862 30882 6914
rect 34750 6862 34802 6914
rect 5966 6750 6018 6802
rect 8318 6750 8370 6802
rect 9550 6750 9602 6802
rect 11678 6750 11730 6802
rect 12014 6750 12066 6802
rect 17390 6750 17442 6802
rect 20638 6750 20690 6802
rect 22654 6750 22706 6802
rect 23326 6750 23378 6802
rect 25454 6750 25506 6802
rect 30046 6750 30098 6802
rect 32062 6750 32114 6802
rect 34190 6750 34242 6802
rect 35758 6750 35810 6802
rect 37662 6750 37714 6802
rect 39454 6750 39506 6802
rect 41582 6750 41634 6802
rect 42478 6750 42530 6802
rect 43262 6750 43314 6802
rect 45390 6750 45442 6802
rect 49198 6750 49250 6802
rect 5182 6638 5234 6690
rect 6302 6638 6354 6690
rect 6750 6638 6802 6690
rect 8878 6638 8930 6690
rect 12238 6638 12290 6690
rect 12350 6638 12402 6690
rect 12686 6638 12738 6690
rect 13022 6638 13074 6690
rect 13358 6638 13410 6690
rect 13582 6638 13634 6690
rect 13694 6638 13746 6690
rect 13918 6638 13970 6690
rect 14590 6638 14642 6690
rect 15262 6638 15314 6690
rect 17726 6638 17778 6690
rect 21422 6638 21474 6690
rect 21870 6638 21922 6690
rect 22430 6638 22482 6690
rect 23326 6638 23378 6690
rect 29486 6638 29538 6690
rect 29710 6638 29762 6690
rect 30382 6638 30434 6690
rect 31278 6638 31330 6690
rect 34526 6638 34578 6690
rect 35086 6638 35138 6690
rect 36094 6638 36146 6690
rect 36990 6638 37042 6690
rect 37774 6638 37826 6690
rect 38782 6638 38834 6690
rect 41918 6638 41970 6690
rect 42590 6638 42642 6690
rect 43038 6638 43090 6690
rect 46286 6638 46338 6690
rect 47070 6638 47122 6690
rect 18510 6526 18562 6578
rect 21758 6526 21810 6578
rect 29038 6526 29090 6578
rect 29934 6526 29986 6578
rect 36430 6526 36482 6578
rect 37102 6526 37154 6578
rect 38334 6526 38386 6578
rect 42142 6526 42194 6578
rect 42702 6526 42754 6578
rect 42926 6526 42978 6578
rect 43710 6526 43762 6578
rect 44158 6526 44210 6578
rect 45502 6526 45554 6578
rect 45950 6526 46002 6578
rect 4734 6414 4786 6466
rect 7198 6414 7250 6466
rect 7758 6414 7810 6466
rect 30494 6414 30546 6466
rect 42366 6414 42418 6466
rect 43262 6414 43314 6466
rect 43486 6414 43538 6466
rect 44046 6414 44098 6466
rect 44942 6414 44994 6466
rect 45390 6414 45442 6466
rect 45726 6414 45778 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4734 6078 4786 6130
rect 17726 6078 17778 6130
rect 17838 6078 17890 6130
rect 39118 6078 39170 6130
rect 39902 6078 39954 6130
rect 40014 6078 40066 6130
rect 46734 6078 46786 6130
rect 46846 6078 46898 6130
rect 46958 6078 47010 6130
rect 47518 6078 47570 6130
rect 48750 6078 48802 6130
rect 6190 5966 6242 6018
rect 8990 5966 9042 6018
rect 17950 5966 18002 6018
rect 19630 5966 19682 6018
rect 20750 5966 20802 6018
rect 23550 5966 23602 6018
rect 24222 5966 24274 6018
rect 25454 5966 25506 6018
rect 25790 5966 25842 6018
rect 27134 5966 27186 6018
rect 28590 5966 28642 6018
rect 39230 5966 39282 6018
rect 39454 5966 39506 6018
rect 40126 5966 40178 6018
rect 46510 5966 46562 6018
rect 5518 5854 5570 5906
rect 8654 5854 8706 5906
rect 14366 5854 14418 5906
rect 16158 5854 16210 5906
rect 16942 5854 16994 5906
rect 18622 5854 18674 5906
rect 18958 5854 19010 5906
rect 20078 5854 20130 5906
rect 23662 5854 23714 5906
rect 24446 5854 24498 5906
rect 25902 5854 25954 5906
rect 26910 5854 26962 5906
rect 27806 5854 27858 5906
rect 31838 5854 31890 5906
rect 38334 5854 38386 5906
rect 38670 5854 38722 5906
rect 39006 5854 39058 5906
rect 41246 5854 41298 5906
rect 47182 5854 47234 5906
rect 47742 5854 47794 5906
rect 48974 5854 49026 5906
rect 4286 5742 4338 5794
rect 5182 5742 5234 5794
rect 8318 5742 8370 5794
rect 9998 5742 10050 5794
rect 16270 5742 16322 5794
rect 19070 5742 19122 5794
rect 22878 5742 22930 5794
rect 23214 5742 23266 5794
rect 25566 5742 25618 5794
rect 30718 5742 30770 5794
rect 31950 5742 32002 5794
rect 33742 5742 33794 5794
rect 42926 5742 42978 5794
rect 4286 5630 4338 5682
rect 5070 5630 5122 5682
rect 16718 5630 16770 5682
rect 26574 5630 26626 5682
rect 32398 5630 32450 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 7198 5294 7250 5346
rect 19070 5294 19122 5346
rect 27470 5294 27522 5346
rect 30382 5294 30434 5346
rect 34078 5294 34130 5346
rect 36430 5294 36482 5346
rect 5182 5182 5234 5234
rect 6078 5182 6130 5234
rect 6526 5182 6578 5234
rect 12910 5182 12962 5234
rect 15262 5182 15314 5234
rect 15598 5182 15650 5234
rect 18958 5182 19010 5234
rect 20414 5182 20466 5234
rect 22318 5182 22370 5234
rect 25006 5182 25058 5234
rect 27134 5182 27186 5234
rect 30830 5182 30882 5234
rect 35758 5182 35810 5234
rect 36990 5182 37042 5234
rect 39118 5182 39170 5234
rect 43150 5182 43202 5234
rect 46062 5182 46114 5234
rect 48190 5182 48242 5234
rect 48750 5182 48802 5234
rect 7422 5070 7474 5122
rect 7982 5070 8034 5122
rect 8430 5070 8482 5122
rect 8766 5070 8818 5122
rect 8990 5070 9042 5122
rect 9998 5070 10050 5122
rect 13694 5070 13746 5122
rect 13918 5070 13970 5122
rect 14590 5070 14642 5122
rect 14926 5070 14978 5122
rect 18510 5070 18562 5122
rect 19742 5070 19794 5122
rect 20190 5070 20242 5122
rect 21310 5070 21362 5122
rect 24334 5070 24386 5122
rect 27582 5070 27634 5122
rect 29262 5070 29314 5122
rect 30494 5070 30546 5122
rect 32958 5070 33010 5122
rect 33742 5070 33794 5122
rect 34190 5070 34242 5122
rect 34414 5070 34466 5122
rect 34750 5070 34802 5122
rect 35086 5070 35138 5122
rect 35422 5070 35474 5122
rect 36430 5070 36482 5122
rect 39902 5070 39954 5122
rect 40350 5070 40402 5122
rect 43598 5070 43650 5122
rect 43710 5070 43762 5122
rect 43822 5070 43874 5122
rect 44046 5070 44098 5122
rect 45278 5070 45330 5122
rect 49198 5070 49250 5122
rect 10782 4958 10834 5010
rect 15150 4958 15202 5010
rect 17726 4958 17778 5010
rect 20750 4958 20802 5010
rect 27694 4958 27746 5010
rect 29598 4958 29650 5010
rect 35646 4958 35698 5010
rect 36094 4958 36146 5010
rect 41022 4958 41074 5010
rect 6862 4846 6914 4898
rect 7758 4846 7810 4898
rect 7870 4846 7922 4898
rect 9438 4846 9490 4898
rect 9550 4846 9602 4898
rect 9662 4846 9714 4898
rect 28142 4846 28194 4898
rect 29710 4846 29762 4898
rect 29822 4846 29874 4898
rect 34862 4846 34914 4898
rect 43934 4846 43986 4898
rect 44830 4846 44882 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 4846 4510 4898 4562
rect 8542 4510 8594 4562
rect 12910 4510 12962 4562
rect 13134 4510 13186 4562
rect 20414 4510 20466 4562
rect 24558 4510 24610 4562
rect 32286 4510 32338 4562
rect 33966 4510 34018 4562
rect 48750 4510 48802 4562
rect 49086 4510 49138 4562
rect 16046 4398 16098 4450
rect 24670 4398 24722 4450
rect 25230 4398 25282 4450
rect 25790 4398 25842 4450
rect 26686 4398 26738 4450
rect 26910 4398 26962 4450
rect 27022 4398 27074 4450
rect 30718 4398 30770 4450
rect 31278 4398 31330 4450
rect 31614 4398 31666 4450
rect 32510 4398 32562 4450
rect 33070 4398 33122 4450
rect 35086 4398 35138 4450
rect 41694 4398 41746 4450
rect 44158 4398 44210 4450
rect 44382 4398 44434 4450
rect 48078 4398 48130 4450
rect 5070 4286 5122 4338
rect 9662 4286 9714 4338
rect 13470 4286 13522 4338
rect 16830 4286 16882 4338
rect 17502 4286 17554 4338
rect 24110 4286 24162 4338
rect 25454 4286 25506 4338
rect 26462 4286 26514 4338
rect 27582 4286 27634 4338
rect 31054 4286 31106 4338
rect 33742 4286 33794 4338
rect 34414 4286 34466 4338
rect 37550 4286 37602 4338
rect 40910 4286 40962 4338
rect 44830 4286 44882 4338
rect 5854 4174 5906 4226
rect 7982 4174 8034 4226
rect 8430 4174 8482 4226
rect 10334 4174 10386 4226
rect 12462 4174 12514 4226
rect 13022 4174 13074 4226
rect 13918 4174 13970 4226
rect 20526 4174 20578 4226
rect 21198 4174 21250 4226
rect 23326 4174 23378 4226
rect 25342 4174 25394 4226
rect 26238 4174 26290 4226
rect 28254 4174 28306 4226
rect 30382 4174 30434 4226
rect 31166 4174 31218 4226
rect 37214 4174 37266 4226
rect 43822 4174 43874 4226
rect 44270 4174 44322 4226
rect 45614 4174 45666 4226
rect 47742 4174 47794 4226
rect 8318 4062 8370 4114
rect 18510 4062 18562 4114
rect 24558 4062 24610 4114
rect 26126 4062 26178 4114
rect 32174 4062 32226 4114
rect 38558 4062 38610 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 9550 3726 9602 3778
rect 9886 3726 9938 3778
rect 10446 3726 10498 3778
rect 10782 3726 10834 3778
rect 11342 3726 11394 3778
rect 13246 3726 13298 3778
rect 47406 3726 47458 3778
rect 5070 3614 5122 3666
rect 6526 3614 6578 3666
rect 10222 3614 10274 3666
rect 11230 3614 11282 3666
rect 11790 3614 11842 3666
rect 20862 3614 20914 3666
rect 22990 3614 23042 3666
rect 25342 3614 25394 3666
rect 27470 3614 27522 3666
rect 30494 3614 30546 3666
rect 32958 3614 33010 3666
rect 35086 3614 35138 3666
rect 36766 3614 36818 3666
rect 38894 3614 38946 3666
rect 40798 3614 40850 3666
rect 44718 3614 44770 3666
rect 46846 3614 46898 3666
rect 47518 3614 47570 3666
rect 48750 3614 48802 3666
rect 11678 3502 11730 3554
rect 12014 3502 12066 3554
rect 12238 3502 12290 3554
rect 16382 3502 16434 3554
rect 17054 3502 17106 3554
rect 19742 3502 19794 3554
rect 23774 3502 23826 3554
rect 24558 3502 24610 3554
rect 31390 3502 31442 3554
rect 32286 3502 32338 3554
rect 35982 3502 36034 3554
rect 39790 3502 39842 3554
rect 42814 3502 42866 3554
rect 44046 3502 44098 3554
rect 49198 3502 49250 3554
rect 9774 3390 9826 3442
rect 1710 3278 1762 3330
rect 3166 3278 3218 3330
rect 5518 3278 5570 3330
rect 6750 3278 6802 3330
rect 7422 3278 7474 3330
rect 7870 3278 7922 3330
rect 8318 3278 8370 3330
rect 8766 3278 8818 3330
rect 13134 3334 13186 3386
rect 13246 3390 13298 3442
rect 17278 3390 17330 3442
rect 43038 3390 43090 3442
rect 47630 3390 47682 3442
rect 15374 3278 15426 3330
rect 19182 3278 19234 3330
rect 28366 3278 28418 3330
rect 48078 3278 48130 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 7422 1710 7474 1762
rect 8318 1710 8370 1762
<< metal2 >>
rect 6272 50200 6384 51000
rect 19040 50200 19152 51000
rect 31808 50200 31920 51000
rect 44576 50200 44688 51000
rect 5516 48018 5572 48030
rect 5516 47966 5518 48018
rect 5570 47966 5572 48018
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 5516 46786 5572 47966
rect 6300 46900 6356 50200
rect 6524 48018 6580 48030
rect 6524 47966 6526 48018
rect 6578 47966 6580 48018
rect 6524 47682 6580 47966
rect 6524 47630 6526 47682
rect 6578 47630 6580 47682
rect 6524 47618 6580 47630
rect 19068 47572 19124 50200
rect 31836 48244 31892 50200
rect 31612 48188 31892 48244
rect 44604 48244 44660 50200
rect 48188 48916 48244 48926
rect 44604 48188 44884 48244
rect 30828 48018 30884 48030
rect 30828 47966 30830 48018
rect 30882 47966 30884 48018
rect 19068 47570 19348 47572
rect 19068 47518 19070 47570
rect 19122 47518 19348 47570
rect 19068 47516 19348 47518
rect 19068 47506 19124 47516
rect 19292 47458 19348 47516
rect 30828 47570 30884 47966
rect 30828 47518 30830 47570
rect 30882 47518 30884 47570
rect 30828 47506 30884 47518
rect 31612 48018 31668 48188
rect 31612 47966 31614 48018
rect 31666 47966 31668 48018
rect 19292 47406 19294 47458
rect 19346 47406 19348 47458
rect 19292 47394 19348 47406
rect 31612 47458 31668 47966
rect 33740 48020 33796 48030
rect 31612 47406 31614 47458
rect 31666 47406 31668 47458
rect 31612 47394 31668 47406
rect 32172 47458 32228 47470
rect 32172 47406 32174 47458
rect 32226 47406 32228 47458
rect 6860 47346 6916 47358
rect 6860 47294 6862 47346
rect 6914 47294 6916 47346
rect 6300 46834 6356 46844
rect 6636 47234 6692 47246
rect 6636 47182 6638 47234
rect 6690 47182 6692 47234
rect 5516 46734 5518 46786
rect 5570 46734 5572 46786
rect 5516 46722 5572 46734
rect 6636 46788 6692 47182
rect 6860 46788 6916 47294
rect 15820 47348 15876 47358
rect 11900 46900 11956 46910
rect 6636 46722 6692 46732
rect 6748 46732 6916 46788
rect 8428 46788 8484 46798
rect 6300 46674 6356 46686
rect 6300 46622 6302 46674
rect 6354 46622 6356 46674
rect 3388 46564 3444 46574
rect 3388 46470 3444 46508
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4508 45890 4564 45902
rect 4508 45838 4510 45890
rect 4562 45838 4564 45890
rect 3052 45780 3108 45790
rect 3052 45218 3108 45724
rect 4396 45780 4452 45790
rect 4396 45686 4452 45724
rect 3052 45166 3054 45218
rect 3106 45166 3108 45218
rect 3052 45154 3108 45166
rect 2268 45108 2324 45118
rect 1820 45106 2324 45108
rect 1820 45054 2270 45106
rect 2322 45054 2324 45106
rect 1820 45052 2324 45054
rect 1820 44322 1876 45052
rect 2268 45042 2324 45052
rect 4508 44884 4564 45838
rect 4732 45892 4788 45902
rect 4732 45890 4900 45892
rect 4732 45838 4734 45890
rect 4786 45838 4900 45890
rect 4732 45836 4900 45838
rect 4732 45826 4788 45836
rect 1820 44270 1822 44322
rect 1874 44270 1876 44322
rect 1820 42754 1876 44270
rect 4060 44828 4564 44884
rect 2492 44210 2548 44222
rect 2492 44158 2494 44210
rect 2546 44158 2548 44210
rect 2492 43708 2548 44158
rect 2492 43652 2996 43708
rect 2940 43650 2996 43652
rect 2940 43598 2942 43650
rect 2994 43598 2996 43650
rect 2940 43586 2996 43598
rect 3500 43652 3556 43662
rect 3052 43540 3108 43550
rect 3052 43446 3108 43484
rect 3500 43538 3556 43596
rect 3500 43486 3502 43538
rect 3554 43486 3556 43538
rect 3500 43474 3556 43486
rect 3948 43540 4004 43550
rect 3276 43428 3332 43438
rect 3276 43334 3332 43372
rect 2492 43316 2548 43326
rect 2492 42866 2548 43260
rect 3836 43316 3892 43326
rect 3836 43222 3892 43260
rect 3948 43316 4004 43484
rect 4060 43316 4116 44828
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4620 44434 4676 44446
rect 4620 44382 4622 44434
rect 4674 44382 4676 44434
rect 4620 44324 4676 44382
rect 4620 44258 4676 44268
rect 4844 43652 4900 45836
rect 4956 45890 5012 45902
rect 4956 45838 4958 45890
rect 5010 45838 5012 45890
rect 4956 45780 5012 45838
rect 5852 45892 5908 45902
rect 6300 45892 6356 46622
rect 6748 46562 6804 46732
rect 8428 46694 8484 46732
rect 9548 46788 9604 46798
rect 9604 46732 9716 46788
rect 9548 46722 9604 46732
rect 6748 46510 6750 46562
rect 6802 46510 6804 46562
rect 6748 46498 6804 46510
rect 7084 46674 7140 46686
rect 7084 46622 7086 46674
rect 7138 46622 7140 46674
rect 7084 46564 7140 46622
rect 8092 46674 8148 46686
rect 8092 46622 8094 46674
rect 8146 46622 8148 46674
rect 5852 45890 6020 45892
rect 5852 45838 5854 45890
rect 5906 45838 6020 45890
rect 5852 45836 6020 45838
rect 5852 45826 5908 45836
rect 4956 45714 5012 45724
rect 5180 44996 5236 45006
rect 5180 44902 5236 44940
rect 5852 44996 5908 45006
rect 5964 44996 6020 45836
rect 6300 45826 6356 45836
rect 7084 45890 7140 46508
rect 7084 45838 7086 45890
rect 7138 45838 7140 45890
rect 6748 45778 6804 45790
rect 6748 45726 6750 45778
rect 6802 45726 6804 45778
rect 6076 45668 6132 45678
rect 6076 45574 6132 45612
rect 6076 44996 6132 45006
rect 6748 44996 6804 45726
rect 5964 44994 6244 44996
rect 5964 44942 6078 44994
rect 6130 44942 6244 44994
rect 5964 44940 6244 44942
rect 5740 44324 5796 44334
rect 5740 43764 5796 44268
rect 5852 44322 5908 44940
rect 6076 44930 6132 44940
rect 5852 44270 5854 44322
rect 5906 44270 5908 44322
rect 5852 43988 5908 44270
rect 6188 44322 6244 44940
rect 6748 44930 6804 44940
rect 6188 44270 6190 44322
rect 6242 44270 6244 44322
rect 6188 44258 6244 44270
rect 6076 44212 6132 44222
rect 5852 43922 5908 43932
rect 5964 44210 6132 44212
rect 5964 44158 6078 44210
rect 6130 44158 6132 44210
rect 5964 44156 6132 44158
rect 5740 43698 5796 43708
rect 4844 43586 4900 43596
rect 5628 43652 5684 43662
rect 5628 43558 5684 43596
rect 5292 43426 5348 43438
rect 5292 43374 5294 43426
rect 5346 43374 5348 43426
rect 3948 43314 4116 43316
rect 3948 43262 3950 43314
rect 4002 43262 4116 43314
rect 3948 43260 4116 43262
rect 3948 43250 4004 43260
rect 2492 42814 2494 42866
rect 2546 42814 2548 42866
rect 2492 42802 2548 42814
rect 1820 42702 1822 42754
rect 1874 42702 1876 42754
rect 1820 41860 1876 42702
rect 2268 41860 2324 41870
rect 1820 41858 2324 41860
rect 1820 41806 2270 41858
rect 2322 41806 2324 41858
rect 1820 41804 2324 41806
rect 1820 41186 1876 41804
rect 1820 41134 1822 41186
rect 1874 41134 1876 41186
rect 1820 41122 1876 41134
rect 2156 39620 2212 41804
rect 2268 41794 2324 41804
rect 2492 41076 2548 41086
rect 2492 41074 2660 41076
rect 2492 41022 2494 41074
rect 2546 41022 2660 41074
rect 2492 41020 2660 41022
rect 2492 41010 2548 41020
rect 2604 40290 2660 41020
rect 2604 40238 2606 40290
rect 2658 40238 2660 40290
rect 2604 40226 2660 40238
rect 2716 40514 2772 40526
rect 2716 40462 2718 40514
rect 2770 40462 2772 40514
rect 1820 39618 2212 39620
rect 1820 39566 2158 39618
rect 2210 39566 2212 39618
rect 1820 39564 2212 39566
rect 1820 38834 1876 39564
rect 2156 39554 2212 39564
rect 1820 38782 1822 38834
rect 1874 38782 1876 38834
rect 1820 36482 1876 38782
rect 2492 38722 2548 38734
rect 2492 38670 2494 38722
rect 2546 38670 2548 38722
rect 2492 38276 2548 38670
rect 2604 38276 2660 38286
rect 2492 38274 2660 38276
rect 2492 38222 2606 38274
rect 2658 38222 2660 38274
rect 2492 38220 2660 38222
rect 2604 38210 2660 38220
rect 2716 38052 2772 40462
rect 2940 40404 2996 40414
rect 2940 40290 2996 40348
rect 3724 40404 3780 40414
rect 3724 40310 3780 40348
rect 2940 40238 2942 40290
rect 2994 40238 2996 40290
rect 2940 40226 2996 40238
rect 2940 39506 2996 39518
rect 2940 39454 2942 39506
rect 2994 39454 2996 39506
rect 2940 39396 2996 39454
rect 2940 39330 2996 39340
rect 2940 38724 2996 38734
rect 2940 38274 2996 38668
rect 4060 38668 4116 43260
rect 4172 43316 4228 43326
rect 4172 43222 4228 43260
rect 4284 43316 4340 43326
rect 4732 43316 4788 43326
rect 4284 43314 4788 43316
rect 4284 43262 4286 43314
rect 4338 43262 4734 43314
rect 4786 43262 4788 43314
rect 4284 43260 4788 43262
rect 4284 40516 4340 43260
rect 4732 43250 4788 43260
rect 5068 43314 5124 43326
rect 5068 43262 5070 43314
rect 5122 43262 5124 43314
rect 4956 43204 5012 43214
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4844 43148 4956 43204
rect 4844 42980 4900 43148
rect 4956 43138 5012 43148
rect 4620 42924 4900 42980
rect 4620 42866 4676 42924
rect 4620 42814 4622 42866
rect 4674 42814 4676 42866
rect 4620 42802 4676 42814
rect 5068 42868 5124 43262
rect 5292 43204 5348 43374
rect 5964 43428 6020 44156
rect 6076 44146 6132 44156
rect 6636 44098 6692 44110
rect 6636 44046 6638 44098
rect 6690 44046 6692 44098
rect 6188 43988 6244 43998
rect 6076 43876 6132 43886
rect 6188 43876 6244 43932
rect 6412 43988 6468 43998
rect 6188 43820 6356 43876
rect 6076 43650 6132 43820
rect 6076 43598 6078 43650
rect 6130 43598 6132 43650
rect 6076 43586 6132 43598
rect 6188 43650 6244 43662
rect 6188 43598 6190 43650
rect 6242 43598 6244 43650
rect 6188 43428 6244 43598
rect 6300 43650 6356 43820
rect 6300 43598 6302 43650
rect 6354 43598 6356 43650
rect 6300 43586 6356 43598
rect 6412 43428 6468 43932
rect 6636 43540 6692 44046
rect 7084 43988 7140 45838
rect 7308 46564 7364 46574
rect 7196 45780 7252 45790
rect 7196 45686 7252 45724
rect 7308 45778 7364 46508
rect 8092 46564 8148 46622
rect 8092 46498 8148 46508
rect 8204 46562 8260 46574
rect 8204 46510 8206 46562
rect 8258 46510 8260 46562
rect 7308 45726 7310 45778
rect 7362 45726 7364 45778
rect 7308 45668 7364 45726
rect 7308 45602 7364 45612
rect 7756 45892 7812 45902
rect 7084 43922 7140 43932
rect 7196 45108 7252 45118
rect 7084 43650 7140 43662
rect 7084 43598 7086 43650
rect 7138 43598 7140 43650
rect 6748 43540 6804 43550
rect 6636 43538 6804 43540
rect 6636 43486 6750 43538
rect 6802 43486 6804 43538
rect 6636 43484 6804 43486
rect 5964 43372 6468 43428
rect 5292 43138 5348 43148
rect 6300 43092 6356 43102
rect 5068 42802 5124 42812
rect 6076 42868 6132 42878
rect 6076 42774 6132 42812
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4620 41298 4676 41310
rect 4620 41246 4622 41298
rect 4674 41246 4676 41298
rect 4508 40516 4564 40526
rect 4284 40460 4508 40516
rect 4508 40290 4564 40460
rect 4620 40404 4676 41246
rect 6300 41300 6356 43036
rect 6412 42980 6468 42990
rect 6412 42886 6468 42924
rect 6636 42756 6692 42766
rect 6748 42756 6804 43484
rect 7084 43540 7140 43598
rect 7084 43474 7140 43484
rect 6524 42754 6804 42756
rect 6524 42702 6638 42754
rect 6690 42702 6804 42754
rect 6524 42700 6804 42702
rect 6860 42980 6916 42990
rect 6412 41300 6468 41310
rect 6300 41298 6468 41300
rect 6300 41246 6414 41298
rect 6466 41246 6468 41298
rect 6300 41244 6468 41246
rect 6412 41234 6468 41244
rect 6524 41074 6580 42700
rect 6636 42690 6692 42700
rect 6860 42084 6916 42924
rect 7084 42756 7140 42766
rect 7196 42756 7252 45052
rect 7756 45108 7812 45836
rect 8204 45218 8260 46510
rect 8428 45780 8484 45790
rect 8428 45778 9604 45780
rect 8428 45726 8430 45778
rect 8482 45726 9604 45778
rect 8428 45724 9604 45726
rect 8428 45714 8484 45724
rect 8204 45166 8206 45218
rect 8258 45166 8260 45218
rect 8204 45154 8260 45166
rect 7756 45042 7812 45052
rect 8988 45108 9044 45118
rect 8988 44434 9044 45052
rect 9548 44994 9604 45724
rect 9548 44942 9550 44994
rect 9602 44942 9604 44994
rect 9548 44930 9604 44942
rect 9660 45330 9716 46732
rect 10556 46004 10612 46014
rect 9660 45278 9662 45330
rect 9714 45278 9716 45330
rect 8988 44382 8990 44434
rect 9042 44382 9044 44434
rect 8988 44370 9044 44382
rect 7644 43764 7700 43774
rect 7644 43670 7700 43708
rect 7420 43652 7476 43662
rect 7420 43558 7476 43596
rect 8204 43650 8260 43662
rect 8204 43598 8206 43650
rect 8258 43598 8260 43650
rect 7532 43428 7588 43438
rect 7532 43334 7588 43372
rect 8092 43316 8148 43326
rect 8092 43222 8148 43260
rect 8204 43204 8260 43598
rect 8876 43650 8932 43662
rect 8876 43598 8878 43650
rect 8930 43598 8932 43650
rect 8540 43540 8596 43550
rect 8764 43540 8820 43550
rect 8596 43538 8820 43540
rect 8596 43486 8766 43538
rect 8818 43486 8820 43538
rect 8596 43484 8820 43486
rect 8540 43474 8596 43484
rect 8764 43474 8820 43484
rect 8876 43540 8932 43598
rect 8876 43474 8932 43484
rect 8204 43138 8260 43148
rect 8428 43316 8484 43326
rect 8428 42868 8484 43260
rect 8428 42802 8484 42812
rect 8876 43314 8932 43326
rect 8876 43262 8878 43314
rect 8930 43262 8932 43314
rect 7084 42754 7252 42756
rect 7084 42702 7086 42754
rect 7138 42702 7252 42754
rect 7084 42700 7252 42702
rect 8876 42756 8932 43262
rect 7084 42690 7140 42700
rect 8876 42690 8932 42700
rect 7756 42644 7812 42654
rect 8204 42644 8260 42654
rect 7756 42642 7924 42644
rect 7756 42590 7758 42642
rect 7810 42590 7924 42642
rect 7756 42588 7924 42590
rect 7756 42578 7812 42588
rect 6748 42028 6916 42084
rect 6636 41972 6692 41982
rect 6636 41878 6692 41916
rect 6748 41186 6804 42028
rect 7868 41858 7924 42588
rect 7980 42196 8036 42206
rect 7980 42102 8036 42140
rect 8204 41970 8260 42588
rect 8204 41918 8206 41970
rect 8258 41918 8260 41970
rect 8204 41906 8260 41918
rect 8316 42196 8372 42206
rect 7868 41806 7870 41858
rect 7922 41806 7924 41858
rect 7868 41794 7924 41806
rect 6972 41188 7028 41198
rect 6748 41134 6750 41186
rect 6802 41134 6804 41186
rect 6748 41122 6804 41134
rect 6860 41186 7028 41188
rect 6860 41134 6974 41186
rect 7026 41134 7028 41186
rect 6860 41132 7028 41134
rect 6524 41022 6526 41074
rect 6578 41022 6580 41074
rect 6524 41010 6580 41022
rect 5740 40962 5796 40974
rect 5740 40910 5742 40962
rect 5794 40910 5796 40962
rect 5740 40852 5796 40910
rect 6076 40964 6132 40974
rect 6076 40962 6244 40964
rect 6076 40910 6078 40962
rect 6130 40910 6244 40962
rect 6076 40908 6244 40910
rect 6076 40898 6132 40908
rect 5292 40796 5796 40852
rect 5292 40740 5348 40796
rect 4620 40310 4676 40348
rect 4956 40684 5348 40740
rect 4508 40238 4510 40290
rect 4562 40238 4564 40290
rect 4508 40226 4564 40238
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4956 39620 5012 40684
rect 6188 40628 6244 40908
rect 6860 40740 6916 41132
rect 6972 41122 7028 41132
rect 8316 41074 8372 42140
rect 9660 42196 9716 45278
rect 10444 46002 10612 46004
rect 10444 45950 10558 46002
rect 10610 45950 10612 46002
rect 10444 45948 10612 45950
rect 9884 44882 9940 44894
rect 9884 44830 9886 44882
rect 9938 44830 9940 44882
rect 9772 43428 9828 43438
rect 9772 43334 9828 43372
rect 9884 43314 9940 44830
rect 10444 43540 10500 45948
rect 10556 45938 10612 45948
rect 11452 43650 11508 43662
rect 11452 43598 11454 43650
rect 11506 43598 11508 43650
rect 10444 43446 10500 43484
rect 10892 43538 10948 43550
rect 10892 43486 10894 43538
rect 10946 43486 10948 43538
rect 10780 43428 10836 43438
rect 10892 43428 10948 43486
rect 11228 43540 11284 43550
rect 11228 43446 11284 43484
rect 10836 43372 10948 43428
rect 10780 43362 10836 43372
rect 9884 43262 9886 43314
rect 9938 43262 9940 43314
rect 9884 43250 9940 43262
rect 10444 43316 10500 43326
rect 11116 43316 11172 43326
rect 9884 42868 9940 42878
rect 9884 42774 9940 42812
rect 10332 42756 10388 42766
rect 10332 42662 10388 42700
rect 10220 42644 10276 42654
rect 10220 42550 10276 42588
rect 9660 42130 9716 42140
rect 8652 41972 8708 41982
rect 8652 41878 8708 41916
rect 9996 41970 10052 41982
rect 9996 41918 9998 41970
rect 10050 41918 10052 41970
rect 8316 41022 8318 41074
rect 8370 41022 8372 41074
rect 8316 41010 8372 41022
rect 9548 41298 9604 41310
rect 9548 41246 9550 41298
rect 9602 41246 9604 41298
rect 5068 40516 5124 40526
rect 5068 40402 5124 40460
rect 5068 40350 5070 40402
rect 5122 40350 5124 40402
rect 5068 40338 5124 40350
rect 5404 40516 5460 40526
rect 5404 40402 5460 40460
rect 5404 40350 5406 40402
rect 5458 40350 5460 40402
rect 5404 40338 5460 40350
rect 5740 40402 5796 40414
rect 5740 40350 5742 40402
rect 5794 40350 5796 40402
rect 5292 40290 5348 40302
rect 5292 40238 5294 40290
rect 5346 40238 5348 40290
rect 5068 40068 5124 40078
rect 5068 39730 5124 40012
rect 5292 39956 5348 40238
rect 5740 40292 5796 40350
rect 6076 40292 6132 40302
rect 5740 40290 6132 40292
rect 5740 40238 6078 40290
rect 6130 40238 6132 40290
rect 5740 40236 6132 40238
rect 6076 40068 6132 40236
rect 6076 40002 6132 40012
rect 5292 39900 5684 39956
rect 5068 39678 5070 39730
rect 5122 39678 5124 39730
rect 5068 39666 5124 39678
rect 4620 38724 4676 38734
rect 4956 38724 5012 39564
rect 5628 39618 5684 39900
rect 6188 39844 6244 40572
rect 6636 40684 6916 40740
rect 7420 40964 7476 40974
rect 7644 40964 7700 40974
rect 7420 40962 7700 40964
rect 7420 40910 7422 40962
rect 7474 40910 7646 40962
rect 7698 40910 7700 40962
rect 7420 40908 7700 40910
rect 6636 40626 6692 40684
rect 6636 40574 6638 40626
rect 6690 40574 6692 40626
rect 6636 40562 6692 40574
rect 6300 40404 6356 40414
rect 6300 40310 6356 40348
rect 5964 39788 6244 39844
rect 6748 40068 6804 40078
rect 5628 39566 5630 39618
rect 5682 39566 5684 39618
rect 5628 39554 5684 39566
rect 5852 39618 5908 39630
rect 5852 39566 5854 39618
rect 5906 39566 5908 39618
rect 5852 39508 5908 39566
rect 5740 39396 5796 39406
rect 5740 39302 5796 39340
rect 4620 38722 5012 38724
rect 4620 38670 4622 38722
rect 4674 38670 5012 38722
rect 4620 38668 5012 38670
rect 5292 38724 5348 38762
rect 4060 38612 4340 38668
rect 4620 38658 4676 38668
rect 5292 38658 5348 38668
rect 5852 38722 5908 39452
rect 5964 38948 6020 39788
rect 6076 39620 6132 39630
rect 6076 39618 6468 39620
rect 6076 39566 6078 39618
rect 6130 39566 6468 39618
rect 6076 39564 6468 39566
rect 6076 39554 6132 39564
rect 5964 38834 6020 38892
rect 5964 38782 5966 38834
rect 6018 38782 6020 38834
rect 5964 38770 6020 38782
rect 5852 38670 5854 38722
rect 5906 38670 5908 38722
rect 5852 38658 5908 38670
rect 2940 38222 2942 38274
rect 2994 38222 2996 38274
rect 2940 38210 2996 38222
rect 2716 37938 2772 37996
rect 2716 37886 2718 37938
rect 2770 37886 2772 37938
rect 2716 37874 2772 37886
rect 1932 37492 1988 37502
rect 3276 37492 3332 37502
rect 1932 37490 3332 37492
rect 1932 37438 1934 37490
rect 1986 37438 3278 37490
rect 3330 37438 3332 37490
rect 1932 37436 3332 37438
rect 1932 37426 1988 37436
rect 2268 37266 2324 37278
rect 2268 37214 2270 37266
rect 2322 37214 2324 37266
rect 2268 36708 2324 37214
rect 3052 37266 3108 37278
rect 3052 37214 3054 37266
rect 3106 37214 3108 37266
rect 2268 36642 2324 36652
rect 2828 36708 2884 36718
rect 1820 36430 1822 36482
rect 1874 36430 1876 36482
rect 1820 36418 1876 36430
rect 2492 36370 2548 36382
rect 2492 36318 2494 36370
rect 2546 36318 2548 36370
rect 2492 35924 2548 36318
rect 2604 35924 2660 35934
rect 2492 35922 2660 35924
rect 2492 35870 2606 35922
rect 2658 35870 2660 35922
rect 2492 35868 2660 35870
rect 2604 35858 2660 35868
rect 2268 35476 2324 35486
rect 2268 35474 2436 35476
rect 2268 35422 2270 35474
rect 2322 35422 2436 35474
rect 2268 35420 2436 35422
rect 2268 35410 2324 35420
rect 1932 35252 1988 35262
rect 1932 34804 1988 35196
rect 1708 34802 1988 34804
rect 1708 34750 1934 34802
rect 1986 34750 1988 34802
rect 1708 34748 1988 34750
rect 1708 34244 1764 34748
rect 1932 34738 1988 34748
rect 2268 34692 2324 34702
rect 2268 34598 2324 34636
rect 1932 34354 1988 34366
rect 1932 34302 1934 34354
rect 1986 34302 1988 34354
rect 1708 34242 1876 34244
rect 1708 34190 1710 34242
rect 1762 34190 1876 34242
rect 1708 34188 1876 34190
rect 1708 34178 1764 34188
rect 1820 32562 1876 34188
rect 1820 32510 1822 32562
rect 1874 32510 1876 32562
rect 1820 32498 1876 32510
rect 1932 32452 1988 34302
rect 2268 34356 2324 34366
rect 2268 34242 2324 34300
rect 2268 34190 2270 34242
rect 2322 34190 2324 34242
rect 2268 34178 2324 34190
rect 2044 34132 2100 34142
rect 2044 34038 2100 34076
rect 1932 32386 1988 32396
rect 2156 33346 2212 33358
rect 2156 33294 2158 33346
rect 2210 33294 2212 33346
rect 2044 32338 2100 32350
rect 2044 32286 2046 32338
rect 2098 32286 2100 32338
rect 1820 32004 1876 32014
rect 1820 31778 1876 31948
rect 1820 31726 1822 31778
rect 1874 31726 1876 31778
rect 1820 30210 1876 31726
rect 2044 30884 2100 32286
rect 2156 32004 2212 33294
rect 2268 32564 2324 32574
rect 2380 32564 2436 35420
rect 2492 35474 2548 35486
rect 2492 35422 2494 35474
rect 2546 35422 2548 35474
rect 2492 35140 2548 35422
rect 2492 35074 2548 35084
rect 2604 35474 2660 35486
rect 2604 35422 2606 35474
rect 2658 35422 2660 35474
rect 2604 35138 2660 35422
rect 2604 35086 2606 35138
rect 2658 35086 2660 35138
rect 2604 35074 2660 35086
rect 2716 34804 2772 34814
rect 2716 34356 2772 34748
rect 2716 34242 2772 34300
rect 2716 34190 2718 34242
rect 2770 34190 2772 34242
rect 2716 34178 2772 34190
rect 2828 34242 2884 36652
rect 3052 35252 3108 37214
rect 3052 35186 3108 35196
rect 3164 35028 3220 37436
rect 3276 37426 3332 37436
rect 3500 37378 3556 37390
rect 3500 37326 3502 37378
rect 3554 37326 3556 37378
rect 2828 34190 2830 34242
rect 2882 34190 2884 34242
rect 2828 34178 2884 34190
rect 2940 34914 2996 34926
rect 2940 34862 2942 34914
rect 2994 34862 2996 34914
rect 2940 34692 2996 34862
rect 2940 34130 2996 34636
rect 2940 34078 2942 34130
rect 2994 34078 2996 34130
rect 2940 33908 2996 34078
rect 3164 34132 3220 34972
rect 3388 35698 3444 35710
rect 3388 35646 3390 35698
rect 3442 35646 3444 35698
rect 3388 34916 3444 35646
rect 3500 35476 3556 37326
rect 3612 37044 3668 37054
rect 4284 37044 4340 38612
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 5628 38052 5684 38062
rect 5628 37938 5684 37996
rect 5628 37886 5630 37938
rect 5682 37886 5684 37938
rect 5628 37874 5684 37886
rect 5964 37826 6020 37838
rect 5964 37774 5966 37826
rect 6018 37774 6020 37826
rect 4620 37378 4676 37390
rect 4620 37326 4622 37378
rect 4674 37326 4676 37378
rect 4620 37044 4676 37326
rect 3612 37042 4004 37044
rect 3612 36990 3614 37042
rect 3666 36990 4004 37042
rect 3612 36988 4004 36990
rect 3612 36978 3668 36988
rect 3500 35420 3892 35476
rect 3500 35252 3556 35262
rect 3500 35138 3556 35196
rect 3500 35086 3502 35138
rect 3554 35086 3556 35138
rect 3500 35074 3556 35086
rect 3612 35028 3668 35038
rect 3612 34934 3668 34972
rect 3388 34850 3444 34860
rect 3836 34804 3892 35420
rect 3836 34738 3892 34748
rect 3724 34692 3780 34702
rect 3724 34598 3780 34636
rect 3948 34244 4004 36988
rect 4284 36988 4676 37044
rect 4956 37268 5012 37278
rect 5964 37268 6020 37774
rect 6412 37380 6468 39564
rect 6748 38836 6804 40012
rect 7308 39620 7364 39630
rect 7420 39620 7476 40908
rect 7644 40898 7700 40908
rect 7980 40964 8036 40974
rect 8652 40964 8708 40974
rect 9100 40964 9156 40974
rect 7980 40962 8148 40964
rect 7980 40910 7982 40962
rect 8034 40910 8148 40962
rect 7980 40908 8148 40910
rect 7980 40898 8036 40908
rect 7756 40628 7812 40638
rect 7644 40516 7700 40526
rect 7644 40402 7700 40460
rect 7756 40514 7812 40572
rect 7756 40462 7758 40514
rect 7810 40462 7812 40514
rect 7756 40450 7812 40462
rect 7644 40350 7646 40402
rect 7698 40350 7700 40402
rect 7308 39618 7476 39620
rect 7308 39566 7310 39618
rect 7362 39566 7476 39618
rect 7308 39564 7476 39566
rect 7532 39620 7588 39630
rect 7308 39554 7364 39564
rect 7532 39526 7588 39564
rect 7644 39618 7700 40350
rect 8092 40402 8148 40908
rect 8652 40962 9268 40964
rect 8652 40910 8654 40962
rect 8706 40910 9102 40962
rect 9154 40910 9268 40962
rect 8652 40908 9268 40910
rect 8652 40898 8708 40908
rect 9100 40898 9156 40908
rect 8316 40628 8372 40638
rect 8092 40350 8094 40402
rect 8146 40350 8148 40402
rect 7980 40290 8036 40302
rect 7980 40238 7982 40290
rect 8034 40238 8036 40290
rect 7644 39566 7646 39618
rect 7698 39566 7700 39618
rect 6860 39396 6916 39406
rect 6860 39394 7028 39396
rect 6860 39342 6862 39394
rect 6914 39342 7028 39394
rect 6860 39340 7028 39342
rect 6860 39330 6916 39340
rect 6860 38836 6916 38846
rect 6748 38834 6916 38836
rect 6748 38782 6862 38834
rect 6914 38782 6916 38834
rect 6748 38780 6916 38782
rect 6860 38770 6916 38780
rect 6972 38836 7028 39340
rect 7644 39284 7700 39566
rect 7532 39228 7700 39284
rect 7756 39620 7812 39630
rect 6972 38668 7028 38780
rect 7084 38948 7140 38958
rect 7084 38834 7140 38892
rect 7084 38782 7086 38834
rect 7138 38782 7140 38834
rect 7084 38770 7140 38782
rect 7532 38834 7588 39228
rect 7644 38948 7700 38958
rect 7756 38948 7812 39564
rect 7980 39284 8036 40238
rect 8092 39508 8148 40350
rect 8204 40516 8260 40526
rect 8204 39618 8260 40460
rect 8204 39566 8206 39618
rect 8258 39566 8260 39618
rect 8204 39554 8260 39566
rect 8316 39508 8372 40572
rect 8764 40514 8820 40526
rect 8764 40462 8766 40514
rect 8818 40462 8820 40514
rect 8764 40404 8820 40462
rect 8428 40348 8820 40404
rect 8428 39732 8484 40348
rect 8540 40180 8596 40190
rect 8876 40180 8932 40190
rect 8540 40178 8820 40180
rect 8540 40126 8542 40178
rect 8594 40126 8820 40178
rect 8540 40124 8820 40126
rect 8540 40114 8596 40124
rect 8540 39732 8596 39742
rect 8428 39676 8540 39732
rect 8540 39666 8596 39676
rect 8428 39508 8484 39518
rect 8316 39506 8484 39508
rect 8316 39454 8430 39506
rect 8482 39454 8484 39506
rect 8316 39452 8484 39454
rect 8092 39442 8148 39452
rect 8428 39442 8484 39452
rect 8540 39508 8596 39518
rect 8540 39414 8596 39452
rect 7980 39228 8596 39284
rect 7644 38946 7812 38948
rect 7644 38894 7646 38946
rect 7698 38894 7812 38946
rect 7644 38892 7812 38894
rect 7644 38882 7700 38892
rect 7532 38782 7534 38834
rect 7586 38782 7588 38834
rect 7532 38770 7588 38782
rect 8540 38834 8596 39228
rect 8540 38782 8542 38834
rect 8594 38782 8596 38834
rect 8540 38770 8596 38782
rect 6412 37286 6468 37324
rect 6860 38612 7028 38668
rect 8428 38722 8484 38734
rect 8428 38670 8430 38722
rect 8482 38670 8484 38722
rect 8428 38668 8484 38670
rect 8652 38668 8708 40124
rect 8764 39844 8820 40124
rect 8876 40086 8932 40124
rect 8988 39844 9044 39854
rect 8764 39842 9044 39844
rect 8764 39790 8990 39842
rect 9042 39790 9044 39842
rect 8764 39788 9044 39790
rect 8988 39778 9044 39788
rect 8988 39060 9044 39070
rect 8876 39004 8988 39060
rect 8876 38946 8932 39004
rect 8988 38994 9044 39004
rect 8876 38894 8878 38946
rect 8930 38894 8932 38946
rect 8876 38882 8932 38894
rect 9212 38668 9268 40908
rect 9548 40516 9604 41246
rect 9996 41188 10052 41918
rect 9996 41122 10052 41132
rect 9548 40450 9604 40460
rect 9884 41076 9940 41086
rect 9436 40180 9492 40190
rect 9492 40124 9828 40180
rect 9436 40114 9492 40124
rect 9324 39730 9380 39742
rect 9324 39678 9326 39730
rect 9378 39678 9380 39730
rect 9324 39620 9380 39678
rect 9324 39554 9380 39564
rect 9548 38836 9604 38846
rect 9548 38742 9604 38780
rect 9772 38834 9828 40124
rect 9884 39060 9940 41020
rect 10332 40402 10388 40414
rect 10332 40350 10334 40402
rect 10386 40350 10388 40402
rect 10220 39508 10276 39518
rect 9884 38994 9940 39004
rect 10108 39452 10220 39508
rect 10108 38946 10164 39452
rect 10220 39442 10276 39452
rect 10108 38894 10110 38946
rect 10162 38894 10164 38946
rect 10108 38882 10164 38894
rect 9772 38782 9774 38834
rect 9826 38782 9828 38834
rect 9772 38770 9828 38782
rect 6076 37268 6132 37278
rect 5964 37212 6076 37268
rect 4956 37044 5012 37212
rect 6076 37174 6132 37212
rect 6524 37044 6580 37054
rect 4956 36988 5236 37044
rect 4060 35588 4116 35598
rect 4060 35586 4228 35588
rect 4060 35534 4062 35586
rect 4114 35534 4228 35586
rect 4060 35532 4228 35534
rect 4060 35522 4116 35532
rect 4060 34690 4116 34702
rect 4060 34638 4062 34690
rect 4114 34638 4116 34690
rect 4060 34468 4116 34638
rect 4060 34402 4116 34412
rect 4172 34354 4228 35532
rect 4284 35140 4340 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4620 36596 4676 36606
rect 4620 35476 4676 36540
rect 5068 36370 5124 36382
rect 5068 36318 5070 36370
rect 5122 36318 5124 36370
rect 4956 36258 5012 36270
rect 4956 36206 4958 36258
rect 5010 36206 5012 36258
rect 4620 35420 4900 35476
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4844 35140 4900 35420
rect 4284 35084 4452 35140
rect 4172 34302 4174 34354
rect 4226 34302 4228 34354
rect 4172 34290 4228 34302
rect 4284 34914 4340 34926
rect 4284 34862 4286 34914
rect 4338 34862 4340 34914
rect 4060 34244 4116 34254
rect 3948 34242 4116 34244
rect 3948 34190 4062 34242
rect 4114 34190 4116 34242
rect 3948 34188 4116 34190
rect 4060 34178 4116 34188
rect 3164 34066 3220 34076
rect 3388 33908 3444 33918
rect 2940 33842 2996 33852
rect 3276 33906 3444 33908
rect 3276 33854 3390 33906
rect 3442 33854 3444 33906
rect 3276 33852 3444 33854
rect 2940 33236 2996 33246
rect 2940 33234 3220 33236
rect 2940 33182 2942 33234
rect 2994 33182 3220 33234
rect 2940 33180 3220 33182
rect 2940 33170 2996 33180
rect 3164 32786 3220 33180
rect 3164 32734 3166 32786
rect 3218 32734 3220 32786
rect 3164 32722 3220 32734
rect 2268 32562 2772 32564
rect 2268 32510 2270 32562
rect 2322 32510 2772 32562
rect 2268 32508 2772 32510
rect 2268 32498 2324 32508
rect 2156 31938 2212 31948
rect 2380 32338 2436 32350
rect 2380 32286 2382 32338
rect 2434 32286 2436 32338
rect 2380 31948 2436 32286
rect 2716 32340 2772 32508
rect 3276 32562 3332 33852
rect 3388 33842 3444 33852
rect 4284 33908 4340 34862
rect 4396 34580 4452 35084
rect 4732 35084 4900 35140
rect 4732 34802 4788 35084
rect 4732 34750 4734 34802
rect 4786 34750 4788 34802
rect 4732 34692 4788 34750
rect 4732 34626 4788 34636
rect 4844 34802 4900 34814
rect 4844 34750 4846 34802
rect 4898 34750 4900 34802
rect 4844 34580 4900 34750
rect 4396 34524 4676 34580
rect 4508 34356 4564 34366
rect 4396 34130 4452 34142
rect 4396 34078 4398 34130
rect 4450 34078 4452 34130
rect 4396 33908 4452 34078
rect 4508 34130 4564 34300
rect 4508 34078 4510 34130
rect 4562 34078 4564 34130
rect 4508 34066 4564 34078
rect 4620 34130 4676 34524
rect 4844 34514 4900 34524
rect 4620 34078 4622 34130
rect 4674 34078 4676 34130
rect 4620 34066 4676 34078
rect 4956 33908 5012 36206
rect 5068 35028 5124 36318
rect 5068 34934 5124 34972
rect 4396 33852 5012 33908
rect 4284 32676 4340 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 5068 33460 5124 33470
rect 5068 33366 5124 33404
rect 3276 32510 3278 32562
rect 3330 32510 3332 32562
rect 3276 32498 3332 32510
rect 3948 32620 4340 32676
rect 3052 32452 3108 32462
rect 3052 32358 3108 32396
rect 2828 32340 2884 32350
rect 2716 32338 2884 32340
rect 2716 32286 2830 32338
rect 2882 32286 2884 32338
rect 2716 32284 2884 32286
rect 2828 31948 2884 32284
rect 2268 31892 2324 31902
rect 2380 31892 2548 31948
rect 2828 31892 3108 31948
rect 2268 31220 2324 31836
rect 2492 31890 2548 31892
rect 2492 31838 2494 31890
rect 2546 31838 2548 31890
rect 2492 31826 2548 31838
rect 2380 31220 2436 31230
rect 2268 31218 2436 31220
rect 2268 31166 2382 31218
rect 2434 31166 2436 31218
rect 2268 31164 2436 31166
rect 2380 31154 2436 31164
rect 2604 30996 2660 31006
rect 2604 30902 2660 30940
rect 2268 30884 2324 30894
rect 2044 30882 2324 30884
rect 2044 30830 2270 30882
rect 2322 30830 2324 30882
rect 2044 30828 2324 30830
rect 2268 30818 2324 30828
rect 2940 30772 2996 30782
rect 2716 30770 2996 30772
rect 2716 30718 2942 30770
rect 2994 30718 2996 30770
rect 2716 30716 2996 30718
rect 2716 30436 2772 30716
rect 2940 30706 2996 30716
rect 3052 30770 3108 31892
rect 3500 30996 3556 31006
rect 3500 30902 3556 30940
rect 3052 30718 3054 30770
rect 3106 30718 3108 30770
rect 2492 30380 2772 30436
rect 3052 30436 3108 30718
rect 2492 30322 2548 30380
rect 3052 30370 3108 30380
rect 3276 30770 3332 30782
rect 3276 30718 3278 30770
rect 3330 30718 3332 30770
rect 2492 30270 2494 30322
rect 2546 30270 2548 30322
rect 2492 30258 2548 30270
rect 1820 30158 1822 30210
rect 1874 30158 1876 30210
rect 1820 30146 1876 30158
rect 3276 29650 3332 30718
rect 3276 29598 3278 29650
rect 3330 29598 3332 29650
rect 3276 29586 3332 29598
rect 3164 29428 3220 29438
rect 3164 29426 3332 29428
rect 3164 29374 3166 29426
rect 3218 29374 3332 29426
rect 3164 29372 3332 29374
rect 3164 29362 3220 29372
rect 3276 28756 3332 29372
rect 2604 28644 2660 28654
rect 3276 28644 3332 28700
rect 3500 29426 3556 29438
rect 3500 29374 3502 29426
rect 3554 29374 3556 29426
rect 1820 27858 1876 27870
rect 1820 27806 1822 27858
rect 1874 27806 1876 27858
rect 1820 26292 1876 27806
rect 2492 27746 2548 27758
rect 2492 27694 2494 27746
rect 2546 27694 2548 27746
rect 2492 27298 2548 27694
rect 2492 27246 2494 27298
rect 2546 27246 2548 27298
rect 2492 27234 2548 27246
rect 2604 27186 2660 28588
rect 2604 27134 2606 27186
rect 2658 27134 2660 27186
rect 2604 27122 2660 27134
rect 2940 28642 3332 28644
rect 2940 28590 3278 28642
rect 3330 28590 3332 28642
rect 2940 28588 3332 28590
rect 2492 26964 2548 26974
rect 2492 26402 2548 26908
rect 2940 26962 2996 28588
rect 3276 28578 3332 28588
rect 3388 28644 3444 28654
rect 3388 28550 3444 28588
rect 3500 28532 3556 29374
rect 3724 29426 3780 29438
rect 3724 29374 3726 29426
rect 3778 29374 3780 29426
rect 3612 28644 3668 28654
rect 3612 28532 3668 28588
rect 3500 28530 3668 28532
rect 3500 28478 3502 28530
rect 3554 28478 3668 28530
rect 3500 28476 3668 28478
rect 3724 28532 3780 29374
rect 3948 29426 4004 32620
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4620 31892 4676 31902
rect 4620 31798 4676 31836
rect 4956 31892 5012 31902
rect 5012 31836 5124 31892
rect 4956 31826 5012 31836
rect 4732 31164 5012 31220
rect 4620 31108 4676 31118
rect 4732 31108 4788 31164
rect 4620 31106 4788 31108
rect 4620 31054 4622 31106
rect 4674 31054 4788 31106
rect 4620 31052 4788 31054
rect 4620 31042 4676 31052
rect 4060 30996 4116 31006
rect 4508 30996 4564 31006
rect 4060 30902 4116 30940
rect 4284 30994 4564 30996
rect 4284 30942 4510 30994
rect 4562 30942 4564 30994
rect 4284 30940 4564 30942
rect 4284 29428 4340 30940
rect 4508 30930 4564 30940
rect 4844 30994 4900 31006
rect 4844 30942 4846 30994
rect 4898 30942 4900 30994
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4620 30324 4676 30334
rect 4844 30324 4900 30942
rect 4620 30322 4900 30324
rect 4620 30270 4622 30322
rect 4674 30270 4900 30322
rect 4620 30268 4900 30270
rect 4620 30258 4676 30268
rect 4732 29540 4788 30268
rect 4956 30100 5012 31164
rect 4956 30034 5012 30044
rect 5068 29876 5124 31836
rect 5180 31668 5236 36988
rect 6300 36594 6356 36606
rect 6300 36542 6302 36594
rect 6354 36542 6356 36594
rect 6188 35586 6244 35598
rect 6188 35534 6190 35586
rect 6242 35534 6244 35586
rect 6188 35028 6244 35534
rect 6300 35588 6356 36542
rect 6300 35522 6356 35532
rect 6524 35586 6580 36988
rect 6524 35534 6526 35586
rect 6578 35534 6580 35586
rect 6524 35522 6580 35534
rect 6636 35810 6692 35822
rect 6636 35758 6638 35810
rect 6690 35758 6692 35810
rect 6636 35588 6692 35758
rect 6860 35812 6916 38612
rect 7532 38610 7588 38622
rect 8428 38612 8708 38668
rect 8764 38612 8820 38622
rect 7532 38558 7534 38610
rect 7586 38558 7588 38610
rect 6860 35810 7476 35812
rect 6860 35758 6862 35810
rect 6914 35758 7476 35810
rect 6860 35756 7476 35758
rect 6860 35746 6916 35756
rect 7420 35700 7476 35756
rect 7420 35606 7476 35644
rect 6636 35522 6692 35532
rect 7196 35588 7252 35598
rect 7196 35494 7252 35532
rect 5628 34916 5684 34926
rect 5516 34860 5628 34916
rect 5516 32674 5572 34860
rect 5628 34822 5684 34860
rect 5740 34804 5796 34814
rect 5628 34356 5684 34366
rect 5740 34356 5796 34748
rect 5628 34354 5796 34356
rect 5628 34302 5630 34354
rect 5682 34302 5796 34354
rect 5628 34300 5796 34302
rect 5852 34692 5908 34702
rect 5628 34290 5684 34300
rect 5852 33570 5908 34636
rect 5852 33518 5854 33570
rect 5906 33518 5908 33570
rect 5852 33506 5908 33518
rect 5964 34130 6020 34142
rect 5964 34078 5966 34130
rect 6018 34078 6020 34130
rect 5964 33572 6020 34078
rect 6076 33572 6132 33582
rect 5964 33570 6132 33572
rect 5964 33518 6078 33570
rect 6130 33518 6132 33570
rect 5964 33516 6132 33518
rect 6188 33572 6244 34972
rect 7308 35028 7364 35038
rect 6412 34802 6468 34814
rect 6412 34750 6414 34802
rect 6466 34750 6468 34802
rect 6300 34356 6356 34366
rect 6300 34242 6356 34300
rect 6412 34354 6468 34750
rect 6412 34302 6414 34354
rect 6466 34302 6468 34354
rect 6412 34290 6468 34302
rect 6300 34190 6302 34242
rect 6354 34190 6356 34242
rect 6300 34178 6356 34190
rect 7308 34242 7364 34972
rect 7532 34356 7588 38558
rect 8540 37380 8596 37390
rect 8092 37266 8148 37278
rect 8092 37214 8094 37266
rect 8146 37214 8148 37266
rect 8092 36596 8148 37214
rect 8540 37268 8596 37324
rect 8764 37268 8820 38556
rect 8540 37266 8820 37268
rect 8540 37214 8542 37266
rect 8594 37214 8820 37266
rect 8540 37212 8820 37214
rect 8876 38612 9268 38668
rect 10332 38668 10388 40350
rect 10444 40402 10500 43260
rect 10892 43314 11172 43316
rect 10892 43262 11118 43314
rect 11170 43262 11172 43314
rect 10892 43260 11172 43262
rect 10780 42756 10836 42766
rect 10780 42662 10836 42700
rect 10668 41858 10724 41870
rect 10668 41806 10670 41858
rect 10722 41806 10724 41858
rect 10444 40350 10446 40402
rect 10498 40350 10500 40402
rect 10444 40338 10500 40350
rect 10556 40964 10612 40974
rect 10556 40402 10612 40908
rect 10668 40626 10724 41806
rect 10668 40574 10670 40626
rect 10722 40574 10724 40626
rect 10668 40562 10724 40574
rect 10892 40514 10948 43260
rect 11116 43250 11172 43260
rect 11452 42756 11508 43598
rect 11564 42980 11620 42990
rect 11564 42886 11620 42924
rect 11452 42690 11508 42700
rect 11676 41076 11732 41086
rect 11676 40982 11732 41020
rect 10892 40462 10894 40514
rect 10946 40462 10948 40514
rect 10892 40450 10948 40462
rect 10556 40350 10558 40402
rect 10610 40350 10612 40402
rect 10556 40338 10612 40350
rect 11452 39508 11508 39518
rect 11452 39414 11508 39452
rect 11900 38668 11956 46844
rect 12236 44322 12292 44334
rect 12236 44270 12238 44322
rect 12290 44270 12292 44322
rect 12236 44100 12292 44270
rect 12684 44100 12740 44110
rect 12236 44098 12740 44100
rect 12236 44046 12686 44098
rect 12738 44046 12740 44098
rect 12236 44044 12740 44046
rect 12012 43540 12068 43550
rect 12012 42754 12068 43484
rect 12012 42702 12014 42754
rect 12066 42702 12068 42754
rect 12012 42690 12068 42702
rect 12124 42756 12180 42766
rect 12124 42662 12180 42700
rect 12348 42756 12404 42766
rect 12348 42754 12628 42756
rect 12348 42702 12350 42754
rect 12402 42702 12628 42754
rect 12348 42700 12628 42702
rect 12348 42690 12404 42700
rect 12572 41748 12628 42700
rect 12684 41972 12740 44044
rect 13916 43540 13972 43550
rect 13580 43538 13972 43540
rect 13580 43486 13918 43538
rect 13970 43486 13972 43538
rect 13580 43484 13972 43486
rect 12684 41906 12740 41916
rect 13468 41970 13524 41982
rect 13468 41918 13470 41970
rect 13522 41918 13524 41970
rect 12796 41858 12852 41870
rect 12796 41806 12798 41858
rect 12850 41806 12852 41858
rect 12796 41748 12852 41806
rect 12572 41692 12964 41748
rect 12908 41298 12964 41692
rect 12908 41246 12910 41298
rect 12962 41246 12964 41298
rect 12908 41234 12964 41246
rect 12460 41188 12516 41198
rect 12236 41132 12460 41188
rect 12236 39620 12292 41132
rect 12460 41094 12516 41132
rect 12796 40964 12852 40974
rect 12796 40870 12852 40908
rect 13468 39844 13524 41918
rect 13580 41188 13636 43484
rect 13916 43474 13972 43484
rect 14700 43428 14756 43438
rect 14700 43426 14868 43428
rect 14700 43374 14702 43426
rect 14754 43374 14868 43426
rect 14700 43372 14868 43374
rect 14700 43362 14756 43372
rect 14812 42642 14868 43372
rect 14812 42590 14814 42642
rect 14866 42590 14868 42642
rect 14812 42578 14868 42590
rect 15148 42644 15204 42654
rect 15148 42550 15204 42588
rect 13804 42082 13860 42094
rect 13804 42030 13806 42082
rect 13858 42030 13860 42082
rect 13804 41300 13860 42030
rect 14252 41300 14308 41310
rect 13804 41298 14308 41300
rect 13804 41246 14254 41298
rect 14306 41246 14308 41298
rect 13804 41244 14308 41246
rect 14252 41234 14308 41244
rect 13580 40514 13636 41132
rect 13580 40462 13582 40514
rect 13634 40462 13636 40514
rect 13580 40450 13636 40462
rect 13692 39844 13748 39854
rect 13468 39842 13748 39844
rect 13468 39790 13694 39842
rect 13746 39790 13748 39842
rect 13468 39788 13748 39790
rect 13692 39778 13748 39788
rect 12236 39618 12516 39620
rect 12236 39566 12238 39618
rect 12290 39566 12516 39618
rect 12236 39564 12516 39566
rect 12236 39554 12292 39564
rect 12460 38834 12516 39564
rect 12460 38782 12462 38834
rect 12514 38782 12516 38834
rect 9996 38612 10052 38622
rect 10332 38612 10612 38668
rect 11900 38612 12068 38668
rect 8540 37202 8596 37212
rect 8316 37044 8372 37054
rect 8316 36950 8372 36988
rect 8652 37042 8708 37054
rect 8652 36990 8654 37042
rect 8706 36990 8708 37042
rect 8652 36708 8708 36990
rect 7756 35924 7812 35934
rect 8092 35924 8148 36540
rect 8428 36652 8708 36708
rect 8428 36594 8484 36652
rect 8876 36596 8932 38612
rect 9996 38518 10052 38556
rect 10556 38052 10612 38612
rect 10556 37958 10612 37996
rect 10892 37938 10948 37950
rect 10892 37886 10894 37938
rect 10946 37886 10948 37938
rect 10780 37828 10836 37838
rect 10780 37734 10836 37772
rect 8428 36542 8430 36594
rect 8482 36542 8484 36594
rect 8428 36530 8484 36542
rect 8764 36540 8932 36596
rect 9660 37154 9716 37166
rect 9660 37102 9662 37154
rect 9714 37102 9716 37154
rect 7756 35922 8148 35924
rect 7756 35870 7758 35922
rect 7810 35870 8148 35922
rect 7756 35868 8148 35870
rect 7756 35858 7812 35868
rect 8316 35700 8372 35710
rect 8316 35606 8372 35644
rect 8652 35700 8708 35710
rect 8652 35606 8708 35644
rect 7980 35474 8036 35486
rect 7980 35422 7982 35474
rect 8034 35422 8036 35474
rect 7980 35140 8036 35422
rect 7980 35074 8036 35084
rect 8540 35028 8596 35038
rect 8540 34934 8596 34972
rect 7756 34356 7812 34366
rect 7532 34354 7812 34356
rect 7532 34302 7758 34354
rect 7810 34302 7812 34354
rect 7532 34300 7812 34302
rect 7756 34290 7812 34300
rect 7868 34356 7924 34366
rect 7308 34190 7310 34242
rect 7362 34190 7364 34242
rect 7308 34178 7364 34190
rect 7868 34242 7924 34300
rect 7868 34190 7870 34242
rect 7922 34190 7924 34242
rect 7868 34178 7924 34190
rect 6636 34130 6692 34142
rect 6636 34078 6638 34130
rect 6690 34078 6692 34130
rect 6636 33908 6692 34078
rect 7196 33908 7252 33918
rect 6636 33906 7252 33908
rect 6636 33854 7198 33906
rect 7250 33854 7252 33906
rect 6636 33852 7252 33854
rect 6300 33572 6356 33582
rect 6188 33570 6356 33572
rect 6188 33518 6302 33570
rect 6354 33518 6356 33570
rect 6188 33516 6356 33518
rect 7196 33572 7252 33852
rect 7756 33908 7812 33918
rect 7756 33906 7924 33908
rect 7756 33854 7758 33906
rect 7810 33854 7924 33906
rect 7756 33852 7924 33854
rect 7756 33842 7812 33852
rect 7196 33516 7476 33572
rect 5964 33460 6020 33516
rect 6076 33506 6132 33516
rect 6300 33506 6356 33516
rect 7420 33460 7476 33516
rect 7420 33404 7700 33460
rect 5964 33394 6020 33404
rect 5516 32622 5518 32674
rect 5570 32622 5572 32674
rect 5516 32004 5572 32622
rect 5516 31938 5572 31948
rect 5628 33346 5684 33358
rect 5628 33294 5630 33346
rect 5682 33294 5684 33346
rect 5628 31892 5684 33294
rect 7308 33346 7364 33358
rect 7308 33294 7310 33346
rect 7362 33294 7364 33346
rect 6412 33236 6468 33246
rect 6972 33236 7028 33246
rect 7308 33236 7364 33294
rect 6412 33234 6580 33236
rect 6412 33182 6414 33234
rect 6466 33182 6580 33234
rect 6412 33180 6580 33182
rect 6412 33170 6468 33180
rect 5628 31826 5684 31836
rect 5964 32004 6020 32014
rect 5964 31778 6020 31948
rect 5964 31726 5966 31778
rect 6018 31726 6020 31778
rect 5964 31714 6020 31726
rect 5180 31612 5684 31668
rect 4956 29820 5124 29876
rect 5292 30100 5348 30110
rect 4844 29540 4900 29550
rect 4732 29538 4900 29540
rect 4732 29486 4846 29538
rect 4898 29486 4900 29538
rect 4732 29484 4900 29486
rect 3948 29374 3950 29426
rect 4002 29374 4004 29426
rect 3948 29362 4004 29374
rect 4060 29426 4340 29428
rect 4060 29374 4286 29426
rect 4338 29374 4340 29426
rect 4060 29372 4340 29374
rect 4060 28868 4116 29372
rect 4284 29362 4340 29372
rect 4620 29428 4676 29438
rect 4620 29334 4676 29372
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 3500 28466 3556 28476
rect 3724 28466 3780 28476
rect 3836 28812 4116 28868
rect 4732 28868 4788 28878
rect 3276 27300 3332 27310
rect 3276 27074 3332 27244
rect 3836 27300 3892 28812
rect 4284 28756 4340 28766
rect 3948 28754 4340 28756
rect 3948 28702 4286 28754
rect 4338 28702 4340 28754
rect 3948 28700 4340 28702
rect 3948 28642 4004 28700
rect 4284 28690 4340 28700
rect 4396 28756 4452 28766
rect 3948 28590 3950 28642
rect 4002 28590 4004 28642
rect 3948 28578 4004 28590
rect 3836 27234 3892 27244
rect 4172 28532 4228 28542
rect 4396 28532 4452 28700
rect 4508 28644 4564 28654
rect 4508 28550 4564 28588
rect 4732 28642 4788 28812
rect 4732 28590 4734 28642
rect 4786 28590 4788 28642
rect 4732 28578 4788 28590
rect 4172 28530 4452 28532
rect 4172 28478 4174 28530
rect 4226 28478 4452 28530
rect 4172 28476 4452 28478
rect 4844 28532 4900 29484
rect 4956 29426 5012 29820
rect 4956 29374 4958 29426
rect 5010 29374 5012 29426
rect 4956 29362 5012 29374
rect 5292 29650 5348 30044
rect 5292 29598 5294 29650
rect 5346 29598 5348 29650
rect 5292 28644 5348 29598
rect 5628 29986 5684 31612
rect 6300 31108 6356 31118
rect 6300 31014 6356 31052
rect 6412 31106 6468 31118
rect 6412 31054 6414 31106
rect 6466 31054 6468 31106
rect 6076 30994 6132 31006
rect 6076 30942 6078 30994
rect 6130 30942 6132 30994
rect 5964 30772 6020 30782
rect 5964 30210 6020 30716
rect 5964 30158 5966 30210
rect 6018 30158 6020 30210
rect 5964 30146 6020 30158
rect 5628 29934 5630 29986
rect 5682 29934 5684 29986
rect 5292 28578 5348 28588
rect 5516 29428 5572 29438
rect 3276 27022 3278 27074
rect 3330 27022 3332 27074
rect 3276 27010 3332 27022
rect 3724 27074 3780 27086
rect 3724 27022 3726 27074
rect 3778 27022 3780 27074
rect 2940 26910 2942 26962
rect 2994 26910 2996 26962
rect 2940 26898 2996 26910
rect 3612 26964 3668 27002
rect 3612 26898 3668 26908
rect 2492 26350 2494 26402
rect 2546 26350 2548 26402
rect 2492 26338 2548 26350
rect 1820 26198 1876 26236
rect 3724 25620 3780 27022
rect 3948 27074 4004 27086
rect 3948 27022 3950 27074
rect 4002 27022 4004 27074
rect 3948 26852 4004 27022
rect 4172 27074 4228 28476
rect 4844 27972 4900 28476
rect 4956 27972 5012 27982
rect 4844 27970 5012 27972
rect 4844 27918 4958 27970
rect 5010 27918 5012 27970
rect 4844 27916 5012 27918
rect 4956 27906 5012 27916
rect 4620 27860 4676 27870
rect 4620 27746 4676 27804
rect 5516 27860 5572 29372
rect 5628 28868 5684 29934
rect 5628 28802 5684 28812
rect 5964 28868 6020 28878
rect 6076 28868 6132 30942
rect 6412 30996 6468 31054
rect 6524 31108 6580 33180
rect 6972 33234 7140 33236
rect 6972 33182 6974 33234
rect 7026 33182 7140 33234
rect 6972 33180 7140 33182
rect 6972 33170 7028 33180
rect 6860 33124 6916 33134
rect 6636 33122 6916 33124
rect 6636 33070 6862 33122
rect 6914 33070 6916 33122
rect 6636 33068 6916 33070
rect 6636 31890 6692 33068
rect 6860 33058 6916 33068
rect 6636 31838 6638 31890
rect 6690 31838 6692 31890
rect 6636 31826 6692 31838
rect 6972 33012 7028 33022
rect 6636 31108 6692 31118
rect 6524 31106 6692 31108
rect 6524 31054 6638 31106
rect 6690 31054 6692 31106
rect 6524 31052 6692 31054
rect 6636 31042 6692 31052
rect 6412 30940 6580 30996
rect 6412 30772 6468 30782
rect 6412 30210 6468 30716
rect 6412 30158 6414 30210
rect 6466 30158 6468 30210
rect 6412 30146 6468 30158
rect 5964 28866 6132 28868
rect 5964 28814 5966 28866
rect 6018 28814 6132 28866
rect 5964 28812 6132 28814
rect 5964 28802 6020 28812
rect 6412 28756 6468 28766
rect 6412 28662 6468 28700
rect 5964 28644 6020 28654
rect 5516 27766 5572 27804
rect 5852 28530 5908 28542
rect 5852 28478 5854 28530
rect 5906 28478 5908 28530
rect 5852 27860 5908 28478
rect 5964 28530 6020 28588
rect 6524 28532 6580 30940
rect 6860 30884 6916 30894
rect 6860 30790 6916 30828
rect 6972 30210 7028 32956
rect 7084 30322 7140 33180
rect 7308 33170 7364 33180
rect 7532 33122 7588 33134
rect 7532 33070 7534 33122
rect 7586 33070 7588 33122
rect 7532 33012 7588 33070
rect 7196 32956 7588 33012
rect 7196 31556 7252 32956
rect 7196 31500 7476 31556
rect 7196 30772 7252 30782
rect 7196 30678 7252 30716
rect 7084 30270 7086 30322
rect 7138 30270 7140 30322
rect 7084 30258 7140 30270
rect 7196 30548 7252 30558
rect 6972 30158 6974 30210
rect 7026 30158 7028 30210
rect 6972 30146 7028 30158
rect 7196 30210 7252 30492
rect 7196 30158 7198 30210
rect 7250 30158 7252 30210
rect 7196 30146 7252 30158
rect 7420 30098 7476 31500
rect 7644 30996 7700 33404
rect 7756 33236 7812 33246
rect 7756 33142 7812 33180
rect 7756 30996 7812 31006
rect 7644 30994 7812 30996
rect 7644 30942 7758 30994
rect 7810 30942 7812 30994
rect 7644 30940 7812 30942
rect 7868 30996 7924 33852
rect 8764 33572 8820 36540
rect 9212 36484 9268 36494
rect 9212 36390 9268 36428
rect 8876 36372 8932 36382
rect 9660 36372 9716 37102
rect 10892 36706 10948 37886
rect 11788 37828 11844 37838
rect 11788 37378 11844 37772
rect 11788 37326 11790 37378
rect 11842 37326 11844 37378
rect 11788 37314 11844 37326
rect 10892 36654 10894 36706
rect 10946 36654 10948 36706
rect 10892 36642 10948 36654
rect 10220 36596 10276 36606
rect 10220 36502 10276 36540
rect 11228 36596 11284 36606
rect 8876 35810 8932 36316
rect 9548 36316 9660 36372
rect 8876 35758 8878 35810
rect 8930 35758 8932 35810
rect 8876 35746 8932 35758
rect 9212 36260 9268 36270
rect 8988 35586 9044 35598
rect 8988 35534 8990 35586
rect 9042 35534 9044 35586
rect 8988 35252 9044 35534
rect 8988 35186 9044 35196
rect 9212 35138 9268 36204
rect 9212 35086 9214 35138
rect 9266 35086 9268 35138
rect 9212 35074 9268 35086
rect 9324 35140 9380 35150
rect 9324 35046 9380 35084
rect 8428 33516 8820 33572
rect 8988 34914 9044 34926
rect 8988 34862 8990 34914
rect 9042 34862 9044 34914
rect 8988 33572 9044 34862
rect 9324 34692 9380 34702
rect 9324 34598 9380 34636
rect 9548 34130 9604 36316
rect 9660 36306 9716 36316
rect 9884 36484 9940 36494
rect 9660 35700 9716 35710
rect 9660 34242 9716 35644
rect 9884 35586 9940 36428
rect 10556 36484 10612 36494
rect 10556 36390 10612 36428
rect 11228 36482 11284 36540
rect 11228 36430 11230 36482
rect 11282 36430 11284 36482
rect 11228 36418 11284 36430
rect 11564 36484 11620 36494
rect 11564 36390 11620 36428
rect 11788 36482 11844 36494
rect 11788 36430 11790 36482
rect 11842 36430 11844 36482
rect 11452 36260 11508 36270
rect 11452 36166 11508 36204
rect 9884 35534 9886 35586
rect 9938 35534 9940 35586
rect 9660 34190 9662 34242
rect 9714 34190 9716 34242
rect 9660 34178 9716 34190
rect 9772 35140 9828 35150
rect 9548 34078 9550 34130
rect 9602 34078 9604 34130
rect 9548 34066 9604 34078
rect 8988 33516 9268 33572
rect 8428 33460 8484 33516
rect 7980 33458 8484 33460
rect 7980 33406 8430 33458
rect 8482 33406 8484 33458
rect 7980 33404 8484 33406
rect 7980 33346 8036 33404
rect 7980 33294 7982 33346
rect 8034 33294 8036 33346
rect 7980 33282 8036 33294
rect 7980 30996 8036 31006
rect 7868 30994 8036 30996
rect 7868 30942 7982 30994
rect 8034 30942 8036 30994
rect 7868 30940 8036 30942
rect 7756 30930 7812 30940
rect 7980 30930 8036 30940
rect 7532 30884 7588 30894
rect 7532 30790 7588 30828
rect 8092 30660 8148 33404
rect 8428 33394 8484 33404
rect 8876 33346 8932 33358
rect 8876 33294 8878 33346
rect 8930 33294 8932 33346
rect 8316 33236 8372 33246
rect 8316 31220 8372 33180
rect 8876 33124 8932 33294
rect 9100 33348 9156 33358
rect 9212 33348 9268 33516
rect 9324 33348 9380 33358
rect 9212 33346 9380 33348
rect 9212 33294 9326 33346
rect 9378 33294 9380 33346
rect 9212 33292 9380 33294
rect 9100 33254 9156 33292
rect 8876 33058 8932 33068
rect 8876 32564 8932 32574
rect 8876 32562 9268 32564
rect 8876 32510 8878 32562
rect 8930 32510 9268 32562
rect 8876 32508 9268 32510
rect 8876 32498 8932 32508
rect 8764 32004 8820 32014
rect 8764 31890 8820 31948
rect 8764 31838 8766 31890
rect 8818 31838 8820 31890
rect 8764 31826 8820 31838
rect 9212 31890 9268 32508
rect 9212 31838 9214 31890
rect 9266 31838 9268 31890
rect 9212 31780 9268 31838
rect 9212 31714 9268 31724
rect 9324 31668 9380 33292
rect 9436 33236 9492 33246
rect 9436 33142 9492 33180
rect 9772 32564 9828 35084
rect 9884 34914 9940 35534
rect 9884 34862 9886 34914
rect 9938 34862 9940 34914
rect 9884 33346 9940 34862
rect 10444 35252 10500 35262
rect 10108 34356 10164 34366
rect 10108 34262 10164 34300
rect 10444 34132 10500 35196
rect 11788 35252 11844 36430
rect 12012 35476 12068 38612
rect 12460 37268 12516 38782
rect 12684 39618 12740 39630
rect 12684 39566 12686 39618
rect 12738 39566 12740 39618
rect 12684 38276 12740 39566
rect 14028 39620 14084 39630
rect 14028 39526 14084 39564
rect 14252 39618 14308 39630
rect 14252 39566 14254 39618
rect 14306 39566 14308 39618
rect 12908 39396 12964 39406
rect 12908 39394 13300 39396
rect 12908 39342 12910 39394
rect 12962 39342 13300 39394
rect 12908 39340 13300 39342
rect 12908 39330 12964 39340
rect 13244 38946 13300 39340
rect 13244 38894 13246 38946
rect 13298 38894 13300 38946
rect 13244 38882 13300 38894
rect 13916 38724 13972 38734
rect 12684 38210 12740 38220
rect 13580 38276 13636 38286
rect 13580 38182 13636 38220
rect 13916 38274 13972 38668
rect 13916 38222 13918 38274
rect 13970 38222 13972 38274
rect 13916 38210 13972 38222
rect 14140 38052 14196 38062
rect 14252 38052 14308 39566
rect 15036 39620 15092 39630
rect 15036 39526 15092 39564
rect 14924 39508 14980 39518
rect 14140 38050 14308 38052
rect 14140 37998 14142 38050
rect 14194 37998 14308 38050
rect 14140 37996 14308 37998
rect 14140 37986 14196 37996
rect 12908 37268 12964 37278
rect 12460 37266 12964 37268
rect 12460 37214 12462 37266
rect 12514 37214 12910 37266
rect 12962 37214 12964 37266
rect 12460 37212 12964 37214
rect 12460 37202 12516 37212
rect 12908 37202 12964 37212
rect 13692 37154 13748 37166
rect 13692 37102 13694 37154
rect 13746 37102 13748 37154
rect 12684 36482 12740 36494
rect 12684 36430 12686 36482
rect 12738 36430 12740 36482
rect 12684 36372 12740 36430
rect 12684 36306 12740 36316
rect 12908 36260 12964 36270
rect 13692 36260 13748 37102
rect 14140 36482 14196 36494
rect 14140 36430 14142 36482
rect 14194 36430 14196 36482
rect 13804 36372 13860 36382
rect 13804 36278 13860 36316
rect 12908 36258 13076 36260
rect 12908 36206 12910 36258
rect 12962 36206 13076 36258
rect 12908 36204 13076 36206
rect 12908 36194 12964 36204
rect 12012 35420 12964 35476
rect 11788 35186 11844 35196
rect 12684 35252 12740 35262
rect 12684 35026 12740 35196
rect 12684 34974 12686 35026
rect 12738 34974 12740 35026
rect 12684 34962 12740 34974
rect 10556 34802 10612 34814
rect 10556 34750 10558 34802
rect 10610 34750 10612 34802
rect 10556 34692 10612 34750
rect 10556 34626 10612 34636
rect 11228 34242 11284 34254
rect 11228 34190 11230 34242
rect 11282 34190 11284 34242
rect 10556 34132 10612 34142
rect 10444 34130 10612 34132
rect 10444 34078 10558 34130
rect 10610 34078 10612 34130
rect 10444 34076 10612 34078
rect 10556 34066 10612 34076
rect 11228 34020 11284 34190
rect 9884 33294 9886 33346
rect 9938 33294 9940 33346
rect 9884 33282 9940 33294
rect 11004 33348 11060 33358
rect 10556 33236 10612 33246
rect 10556 33142 10612 33180
rect 10892 33124 10948 33134
rect 10108 32676 10164 32686
rect 10108 32582 10164 32620
rect 10780 32676 10836 32686
rect 9772 32470 9828 32508
rect 10220 32562 10276 32574
rect 10220 32510 10222 32562
rect 10274 32510 10276 32562
rect 9324 31602 9380 31612
rect 9436 32338 9492 32350
rect 9436 32286 9438 32338
rect 9490 32286 9492 32338
rect 9436 31780 9492 32286
rect 9884 32004 9940 32014
rect 10220 32004 10276 32510
rect 10780 32562 10836 32620
rect 10780 32510 10782 32562
rect 10834 32510 10836 32562
rect 10780 32498 10836 32510
rect 9940 31948 10276 32004
rect 10444 32450 10500 32462
rect 10444 32398 10446 32450
rect 10498 32398 10500 32450
rect 9772 31892 9828 31902
rect 9772 31798 9828 31836
rect 9548 31780 9604 31790
rect 9436 31778 9604 31780
rect 9436 31726 9550 31778
rect 9602 31726 9604 31778
rect 9436 31724 9604 31726
rect 8204 31108 8260 31118
rect 8204 31014 8260 31052
rect 7420 30046 7422 30098
rect 7474 30046 7476 30098
rect 7420 30034 7476 30046
rect 7756 30604 8148 30660
rect 8316 30994 8372 31164
rect 8652 31108 8708 31118
rect 8652 31014 8708 31052
rect 9212 31108 9268 31118
rect 8316 30942 8318 30994
rect 8370 30942 8372 30994
rect 6636 29986 6692 29998
rect 6636 29934 6638 29986
rect 6690 29934 6692 29986
rect 6636 29428 6692 29934
rect 7644 29652 7700 29662
rect 7756 29652 7812 30604
rect 8316 30548 8372 30942
rect 8316 30482 8372 30492
rect 7868 30436 7924 30446
rect 7868 30098 7924 30380
rect 8316 30324 8372 30334
rect 8092 30212 8148 30222
rect 7868 30046 7870 30098
rect 7922 30046 7924 30098
rect 7868 30034 7924 30046
rect 7980 30210 8148 30212
rect 7980 30158 8094 30210
rect 8146 30158 8148 30210
rect 7980 30156 8148 30158
rect 7644 29650 7812 29652
rect 7644 29598 7646 29650
rect 7698 29598 7812 29650
rect 7644 29596 7812 29598
rect 6636 29362 6692 29372
rect 7308 29428 7364 29438
rect 7308 29334 7364 29372
rect 5964 28478 5966 28530
rect 6018 28478 6020 28530
rect 5964 28466 6020 28478
rect 6412 28476 6580 28532
rect 6636 28644 6692 28654
rect 6412 28082 6468 28476
rect 6412 28030 6414 28082
rect 6466 28030 6468 28082
rect 6412 28018 6468 28030
rect 6524 27970 6580 27982
rect 6524 27918 6526 27970
rect 6578 27918 6580 27970
rect 4620 27694 4622 27746
rect 4674 27694 4676 27746
rect 4620 27682 4676 27694
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4508 27300 4564 27310
rect 4508 27206 4564 27244
rect 5068 27300 5124 27310
rect 5068 27188 5124 27244
rect 4956 27186 5124 27188
rect 4956 27134 5070 27186
rect 5122 27134 5124 27186
rect 4956 27132 5124 27134
rect 4172 27022 4174 27074
rect 4226 27022 4228 27074
rect 4172 27010 4228 27022
rect 4844 27076 4900 27086
rect 4844 26982 4900 27020
rect 3948 26786 4004 26796
rect 4956 26292 5012 27132
rect 5068 27122 5124 27132
rect 5292 27076 5348 27086
rect 5068 26852 5124 26862
rect 5124 26796 5236 26852
rect 5068 26786 5124 26796
rect 5180 26514 5236 26796
rect 5180 26462 5182 26514
rect 5234 26462 5236 26514
rect 5180 26450 5236 26462
rect 4620 26290 5012 26292
rect 4620 26238 4958 26290
rect 5010 26238 5012 26290
rect 4620 26236 5012 26238
rect 4620 26178 4676 26236
rect 4956 26226 5012 26236
rect 4620 26126 4622 26178
rect 4674 26126 4676 26178
rect 4620 26114 4676 26126
rect 5292 26066 5348 27020
rect 5292 26014 5294 26066
rect 5346 26014 5348 26066
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4844 25844 4900 25854
rect 4172 25732 4228 25742
rect 4172 25638 4228 25676
rect 4844 25730 4900 25788
rect 4844 25678 4846 25730
rect 4898 25678 4900 25730
rect 4844 25666 4900 25678
rect 5292 25732 5348 26014
rect 5292 25666 5348 25676
rect 3780 25564 3892 25620
rect 3724 25554 3780 25564
rect 1820 24722 1876 24734
rect 1820 24670 1822 24722
rect 1874 24670 1876 24722
rect 1820 23938 1876 24670
rect 2492 24612 2548 24622
rect 2492 24518 2548 24556
rect 3836 24052 3892 25564
rect 5852 25618 5908 27804
rect 5964 27858 6020 27870
rect 5964 27806 5966 27858
rect 6018 27806 6020 27858
rect 5964 27300 6020 27806
rect 6524 27748 6580 27918
rect 6524 27682 6580 27692
rect 5964 27234 6020 27244
rect 6076 27636 6132 27646
rect 6076 27298 6132 27580
rect 6076 27246 6078 27298
rect 6130 27246 6132 27298
rect 6076 25844 6132 27246
rect 6412 27300 6468 27310
rect 6412 27206 6468 27244
rect 6636 27186 6692 28588
rect 7084 28420 7140 28430
rect 7084 27858 7140 28364
rect 7084 27806 7086 27858
rect 7138 27806 7140 27858
rect 6636 27134 6638 27186
rect 6690 27134 6692 27186
rect 6636 27122 6692 27134
rect 6860 27634 6916 27646
rect 6860 27582 6862 27634
rect 6914 27582 6916 27634
rect 6860 26908 6916 27582
rect 7084 27300 7140 27806
rect 7420 27970 7476 27982
rect 7420 27918 7422 27970
rect 7474 27918 7476 27970
rect 7420 27860 7476 27918
rect 7420 27794 7476 27804
rect 7084 27234 7140 27244
rect 6860 26852 7028 26908
rect 6188 26292 6244 26302
rect 6188 26198 6244 26236
rect 6860 26180 6916 26190
rect 6076 25730 6132 25788
rect 6076 25678 6078 25730
rect 6130 25678 6132 25730
rect 6076 25666 6132 25678
rect 6748 26178 6916 26180
rect 6748 26126 6862 26178
rect 6914 26126 6916 26178
rect 6748 26124 6916 26126
rect 6748 25730 6804 26124
rect 6860 26114 6916 26124
rect 6748 25678 6750 25730
rect 6802 25678 6804 25730
rect 6748 25666 6804 25678
rect 6972 25732 7028 26852
rect 7644 26068 7700 29596
rect 7980 29428 8036 30156
rect 8092 30146 8148 30156
rect 8316 29538 8372 30268
rect 9212 30322 9268 31052
rect 9212 30270 9214 30322
rect 9266 30270 9268 30322
rect 9212 30258 9268 30270
rect 8316 29486 8318 29538
rect 8370 29486 8372 29538
rect 8316 29428 8372 29486
rect 7756 28532 7812 28542
rect 7756 27970 7812 28476
rect 7756 27918 7758 27970
rect 7810 27918 7812 27970
rect 7756 27906 7812 27918
rect 7868 27748 7924 27758
rect 7868 27654 7924 27692
rect 7644 26012 7924 26068
rect 7196 25732 7252 25742
rect 6972 25676 7196 25732
rect 7196 25638 7252 25676
rect 5852 25566 5854 25618
rect 5906 25566 5908 25618
rect 5068 25506 5124 25518
rect 5068 25454 5070 25506
rect 5122 25454 5124 25506
rect 3948 25282 4004 25294
rect 3948 25230 3950 25282
rect 4002 25230 4004 25282
rect 3948 25172 4004 25230
rect 3948 25106 4004 25116
rect 4060 25282 4116 25294
rect 4060 25230 4062 25282
rect 4114 25230 4116 25282
rect 4060 24164 4116 25230
rect 4508 25284 4564 25294
rect 4508 25282 4788 25284
rect 4508 25230 4510 25282
rect 4562 25230 4788 25282
rect 4508 25228 4788 25230
rect 4508 25218 4564 25228
rect 4620 24610 4676 24622
rect 4620 24558 4622 24610
rect 4674 24558 4676 24610
rect 4620 24500 4676 24558
rect 4732 24500 4788 25228
rect 5068 25172 5124 25454
rect 5124 25116 5460 25172
rect 5068 25106 5124 25116
rect 5404 24834 5460 25116
rect 5852 24946 5908 25566
rect 5852 24894 5854 24946
rect 5906 24894 5908 24946
rect 5852 24882 5908 24894
rect 6300 25620 6356 25630
rect 5404 24782 5406 24834
rect 5458 24782 5460 24834
rect 5180 24722 5236 24734
rect 5180 24670 5182 24722
rect 5234 24670 5236 24722
rect 5180 24500 5236 24670
rect 4732 24444 4900 24500
rect 4620 24434 4676 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4620 24164 4676 24174
rect 4060 24108 4564 24164
rect 3836 23996 4452 24052
rect 1820 23886 1822 23938
rect 1874 23886 1876 23938
rect 1820 22370 1876 23886
rect 2492 23826 2548 23838
rect 2492 23774 2494 23826
rect 2546 23774 2548 23826
rect 2492 23380 2548 23774
rect 2492 23314 2548 23324
rect 4284 23380 4340 23390
rect 3388 23268 3444 23278
rect 3388 23174 3444 23212
rect 4284 23266 4340 23324
rect 4284 23214 4286 23266
rect 4338 23214 4340 23266
rect 4284 23202 4340 23214
rect 3612 23154 3668 23166
rect 3612 23102 3614 23154
rect 3666 23102 3668 23154
rect 1820 22318 1822 22370
rect 1874 22318 1876 22370
rect 1820 20804 1876 22318
rect 2828 23044 2884 23054
rect 2492 22260 2548 22270
rect 2492 22258 2772 22260
rect 2492 22206 2494 22258
rect 2546 22206 2772 22258
rect 2492 22204 2772 22206
rect 2492 22194 2548 22204
rect 2716 21810 2772 22204
rect 2716 21758 2718 21810
rect 2770 21758 2772 21810
rect 2716 21746 2772 21758
rect 2828 21698 2884 22988
rect 3500 23044 3556 23054
rect 3500 22950 3556 22988
rect 3612 22596 3668 23102
rect 4060 23156 4116 23166
rect 4060 23062 4116 23100
rect 4396 23154 4452 23996
rect 4396 23102 4398 23154
rect 4450 23102 4452 23154
rect 4396 23090 4452 23102
rect 4508 23156 4564 24108
rect 4620 24050 4676 24108
rect 4620 23998 4622 24050
rect 4674 23998 4676 24050
rect 4620 23986 4676 23998
rect 4844 23828 4900 24444
rect 5180 23940 5236 24444
rect 5180 23874 5236 23884
rect 5292 24722 5348 24734
rect 5292 24670 5294 24722
rect 5346 24670 5348 24722
rect 4844 23268 4900 23772
rect 5292 23492 5348 24670
rect 5404 24164 5460 24782
rect 6300 24722 6356 25564
rect 6860 25620 6916 25630
rect 6860 25526 6916 25564
rect 7644 25620 7700 25630
rect 7084 25508 7140 25518
rect 7084 25414 7140 25452
rect 6412 25396 6468 25406
rect 6468 25340 6692 25396
rect 6412 25302 6468 25340
rect 6300 24670 6302 24722
rect 6354 24670 6356 24722
rect 6300 24658 6356 24670
rect 6636 24722 6692 25340
rect 7644 25394 7700 25564
rect 7644 25342 7646 25394
rect 7698 25342 7700 25394
rect 7644 25330 7700 25342
rect 7868 25284 7924 26012
rect 7980 25506 8036 29372
rect 8092 29372 8372 29428
rect 8764 29538 8820 29550
rect 8764 29486 8766 29538
rect 8818 29486 8820 29538
rect 8092 27748 8148 29372
rect 8652 29202 8708 29214
rect 8652 29150 8654 29202
rect 8706 29150 8708 29202
rect 8540 28644 8596 28654
rect 8204 28642 8596 28644
rect 8204 28590 8542 28642
rect 8594 28590 8596 28642
rect 8204 28588 8596 28590
rect 8204 27970 8260 28588
rect 8540 28578 8596 28588
rect 8204 27918 8206 27970
rect 8258 27918 8260 27970
rect 8204 27906 8260 27918
rect 8652 27858 8708 29150
rect 8764 28644 8820 29486
rect 8764 28578 8820 28588
rect 8988 29204 9044 29214
rect 9436 29204 9492 31724
rect 9548 31714 9604 31724
rect 9548 31220 9604 31230
rect 9548 31126 9604 31164
rect 9884 31218 9940 31948
rect 9884 31166 9886 31218
rect 9938 31166 9940 31218
rect 9884 31154 9940 31166
rect 9996 31778 10052 31790
rect 9996 31726 9998 31778
rect 10050 31726 10052 31778
rect 9996 31668 10052 31726
rect 10444 31778 10500 32398
rect 10444 31726 10446 31778
rect 10498 31726 10500 31778
rect 9996 30324 10052 31612
rect 10108 31666 10164 31678
rect 10108 31614 10110 31666
rect 10162 31614 10164 31666
rect 10108 30324 10164 31614
rect 10444 31108 10500 31726
rect 10780 31892 10836 31902
rect 10668 31666 10724 31678
rect 10668 31614 10670 31666
rect 10722 31614 10724 31666
rect 10668 31220 10724 31614
rect 10780 31554 10836 31836
rect 10892 31780 10948 33068
rect 11004 32786 11060 33292
rect 11004 32734 11006 32786
rect 11058 32734 11060 32786
rect 11004 32722 11060 32734
rect 11228 32676 11284 33964
rect 12124 34020 12180 34030
rect 12124 33926 12180 33964
rect 12684 34020 12740 34030
rect 11564 33906 11620 33918
rect 11564 33854 11566 33906
rect 11618 33854 11620 33906
rect 11564 33124 11620 33854
rect 11900 33906 11956 33918
rect 11900 33854 11902 33906
rect 11954 33854 11956 33906
rect 11900 33684 11956 33854
rect 11564 33058 11620 33068
rect 11676 33628 11956 33684
rect 11228 32610 11284 32620
rect 11116 32564 11172 32574
rect 11116 32470 11172 32508
rect 11676 32564 11732 33628
rect 12684 33458 12740 33964
rect 12684 33406 12686 33458
rect 12738 33406 12740 33458
rect 12684 33394 12740 33406
rect 12572 33348 12628 33358
rect 11676 32498 11732 32508
rect 12460 33292 12572 33348
rect 12460 32562 12516 33292
rect 12572 33282 12628 33292
rect 12460 32510 12462 32562
rect 12514 32510 12516 32562
rect 12460 32498 12516 32510
rect 11004 31780 11060 31790
rect 10892 31778 11060 31780
rect 10892 31726 11006 31778
rect 11058 31726 11060 31778
rect 10892 31724 11060 31726
rect 11004 31714 11060 31724
rect 12572 31780 12628 31790
rect 10780 31502 10782 31554
rect 10834 31502 10836 31554
rect 10780 31490 10836 31502
rect 10668 31154 10724 31164
rect 10444 31042 10500 31052
rect 12124 30996 12180 31006
rect 10220 30882 10276 30894
rect 10220 30830 10222 30882
rect 10274 30830 10276 30882
rect 10220 30548 10276 30830
rect 10220 30482 10276 30492
rect 11340 30324 11396 30334
rect 10108 30322 11396 30324
rect 10108 30270 11342 30322
rect 11394 30270 11396 30322
rect 10108 30268 11396 30270
rect 9996 30258 10052 30268
rect 11340 30258 11396 30268
rect 12124 30210 12180 30940
rect 12348 30884 12404 30894
rect 12348 30882 12516 30884
rect 12348 30830 12350 30882
rect 12402 30830 12516 30882
rect 12348 30828 12516 30830
rect 12348 30818 12404 30828
rect 12124 30158 12126 30210
rect 12178 30158 12180 30210
rect 12124 30146 12180 30158
rect 12460 30098 12516 30828
rect 12460 30046 12462 30098
rect 12514 30046 12516 30098
rect 12460 30034 12516 30046
rect 10668 29540 10724 29550
rect 8988 29202 9492 29204
rect 8988 29150 8990 29202
rect 9042 29150 9492 29202
rect 8988 29148 9492 29150
rect 10444 29538 10724 29540
rect 10444 29486 10670 29538
rect 10722 29486 10724 29538
rect 10444 29484 10724 29486
rect 8988 28420 9044 29148
rect 10444 28754 10500 29484
rect 10668 29474 10724 29484
rect 11004 29428 11060 29438
rect 11004 29426 11172 29428
rect 11004 29374 11006 29426
rect 11058 29374 11172 29426
rect 11004 29372 11172 29374
rect 11004 29362 11060 29372
rect 10444 28702 10446 28754
rect 10498 28702 10500 28754
rect 10444 28690 10500 28702
rect 8988 28354 9044 28364
rect 9212 28644 9268 28654
rect 9660 28644 9716 28654
rect 9212 28642 9716 28644
rect 9212 28590 9214 28642
rect 9266 28590 9662 28642
rect 9714 28590 9716 28642
rect 9212 28588 9716 28590
rect 8652 27806 8654 27858
rect 8706 27806 8708 27858
rect 8652 27794 8708 27806
rect 8316 27748 8372 27758
rect 8092 27746 8372 27748
rect 8092 27694 8318 27746
rect 8370 27694 8372 27746
rect 8092 27692 8372 27694
rect 8316 27682 8372 27692
rect 8988 27748 9044 27758
rect 8540 27636 8596 27646
rect 8540 27542 8596 27580
rect 8428 26962 8484 26974
rect 8428 26910 8430 26962
rect 8482 26910 8484 26962
rect 8428 26292 8484 26910
rect 8428 26226 8484 26236
rect 8988 26180 9044 27692
rect 9212 26292 9268 28588
rect 9660 28578 9716 28588
rect 11116 28082 11172 29372
rect 12124 29316 12180 29326
rect 12124 29092 12180 29260
rect 11116 28030 11118 28082
rect 11170 28030 11172 28082
rect 11116 28018 11172 28030
rect 11676 29036 12180 29092
rect 12348 29202 12404 29214
rect 12348 29150 12350 29202
rect 12402 29150 12404 29202
rect 11676 27858 11732 29036
rect 12348 28084 12404 29150
rect 12572 28980 12628 31724
rect 12684 30210 12740 30222
rect 12684 30158 12686 30210
rect 12738 30158 12740 30210
rect 12684 29650 12740 30158
rect 12684 29598 12686 29650
rect 12738 29598 12740 29650
rect 12684 29586 12740 29598
rect 12572 28924 12740 28980
rect 12348 28018 12404 28028
rect 12572 28754 12628 28766
rect 12572 28702 12574 28754
rect 12626 28702 12628 28754
rect 11676 27806 11678 27858
rect 11730 27806 11732 27858
rect 11676 27794 11732 27806
rect 12572 27858 12628 28702
rect 12572 27806 12574 27858
rect 12626 27806 12628 27858
rect 11452 27748 11508 27758
rect 11452 27654 11508 27692
rect 12012 27748 12068 27758
rect 12012 27654 12068 27692
rect 12572 27412 12628 27806
rect 12572 27346 12628 27356
rect 12684 27188 12740 28924
rect 12796 27748 12852 27758
rect 12796 27654 12852 27692
rect 12796 27188 12852 27198
rect 12236 27186 12852 27188
rect 12236 27134 12798 27186
rect 12850 27134 12852 27186
rect 12236 27132 12852 27134
rect 12236 27074 12292 27132
rect 12796 27122 12852 27132
rect 12236 27022 12238 27074
rect 12290 27022 12292 27074
rect 12236 27010 12292 27022
rect 12908 26908 12964 35420
rect 13020 35028 13076 36204
rect 13692 36194 13748 36204
rect 14140 35812 14196 36430
rect 14252 36484 14308 37996
rect 14812 38052 14868 38062
rect 14924 38052 14980 39452
rect 15148 39396 15204 39406
rect 15484 39396 15540 39406
rect 15148 39394 15484 39396
rect 15148 39342 15150 39394
rect 15202 39342 15484 39394
rect 15148 39340 15484 39342
rect 15148 39330 15204 39340
rect 15484 39330 15540 39340
rect 15596 39394 15652 39406
rect 15596 39342 15598 39394
rect 15650 39342 15652 39394
rect 15372 38724 15428 38734
rect 15372 38722 15540 38724
rect 15372 38670 15374 38722
rect 15426 38670 15540 38722
rect 15372 38668 15540 38670
rect 15372 38658 15428 38668
rect 15484 38612 15540 38668
rect 14812 38050 14980 38052
rect 14812 37998 14814 38050
rect 14866 37998 14980 38050
rect 14812 37996 14980 37998
rect 15148 38052 15204 38062
rect 14812 37986 14868 37996
rect 15148 37958 15204 37996
rect 15372 37938 15428 37950
rect 15372 37886 15374 37938
rect 15426 37886 15428 37938
rect 15036 37828 15092 37838
rect 15036 37734 15092 37772
rect 15372 37716 15428 37886
rect 15372 37650 15428 37660
rect 15484 37380 15540 38556
rect 15596 38052 15652 39342
rect 15708 38724 15764 38762
rect 15708 38658 15764 38668
rect 15820 38164 15876 47292
rect 19852 47348 19908 47358
rect 19852 47254 19908 47292
rect 26572 47348 26628 47358
rect 26572 47346 27076 47348
rect 26572 47294 26574 47346
rect 26626 47294 27076 47346
rect 26572 47292 27076 47294
rect 26572 47282 26628 47292
rect 26236 47236 26292 47246
rect 26012 47234 26292 47236
rect 26012 47182 26238 47234
rect 26290 47182 26292 47234
rect 26012 47180 26292 47182
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 26012 46786 26068 47180
rect 26236 47170 26292 47180
rect 26012 46734 26014 46786
rect 26066 46734 26068 46786
rect 26012 46722 26068 46734
rect 21644 46674 21700 46686
rect 21644 46622 21646 46674
rect 21698 46622 21700 46674
rect 18844 46562 18900 46574
rect 20972 46564 21028 46574
rect 18844 46510 18846 46562
rect 18898 46510 18900 46562
rect 18396 45220 18452 45230
rect 18844 45220 18900 46510
rect 20412 46562 21028 46564
rect 20412 46510 20974 46562
rect 21026 46510 21028 46562
rect 20412 46508 21028 46510
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 16492 44324 16548 44334
rect 16492 44230 16548 44268
rect 18396 44324 18452 45164
rect 17164 44212 17220 44222
rect 17164 44210 17444 44212
rect 17164 44158 17166 44210
rect 17218 44158 17444 44210
rect 17164 44156 17444 44158
rect 17164 44146 17220 44156
rect 17388 43762 17444 44156
rect 17388 43710 17390 43762
rect 17442 43710 17444 43762
rect 17388 43698 17444 43710
rect 17724 43540 17780 43550
rect 17724 43538 18004 43540
rect 17724 43486 17726 43538
rect 17778 43486 18004 43538
rect 17724 43484 18004 43486
rect 17724 43474 17780 43484
rect 16828 43428 16884 43438
rect 16828 43426 16996 43428
rect 16828 43374 16830 43426
rect 16882 43374 16996 43426
rect 16828 43372 16996 43374
rect 16828 43362 16884 43372
rect 16828 42754 16884 42766
rect 16828 42702 16830 42754
rect 16882 42702 16884 42754
rect 16492 42644 16548 42654
rect 16492 42550 16548 42588
rect 16828 42082 16884 42702
rect 16828 42030 16830 42082
rect 16882 42030 16884 42082
rect 16828 42018 16884 42030
rect 16380 41970 16436 41982
rect 16380 41918 16382 41970
rect 16434 41918 16436 41970
rect 16380 41860 16436 41918
rect 16380 41794 16436 41804
rect 16716 41970 16772 41982
rect 16716 41918 16718 41970
rect 16770 41918 16772 41970
rect 16380 41300 16436 41310
rect 16156 40292 16212 40302
rect 16156 39508 16212 40236
rect 16380 39618 16436 41244
rect 16716 41188 16772 41918
rect 16940 41860 16996 43372
rect 17052 42754 17108 42766
rect 17052 42702 17054 42754
rect 17106 42702 17108 42754
rect 17052 41860 17108 42702
rect 17948 42194 18004 43484
rect 18396 43538 18452 44268
rect 18396 43486 18398 43538
rect 18450 43486 18452 43538
rect 18396 43474 18452 43486
rect 18508 45164 18900 45220
rect 18508 44436 18564 45164
rect 18508 43316 18564 44380
rect 18396 43260 18564 43316
rect 18732 44994 18788 45006
rect 18732 44942 18734 44994
rect 18786 44942 18788 44994
rect 18396 42866 18452 43260
rect 18396 42814 18398 42866
rect 18450 42814 18452 42866
rect 18396 42802 18452 42814
rect 18284 42532 18340 42542
rect 18620 42532 18676 42542
rect 18284 42438 18340 42476
rect 18508 42476 18620 42532
rect 17948 42142 17950 42194
rect 18002 42142 18004 42194
rect 17948 42130 18004 42142
rect 18508 42084 18564 42476
rect 18620 42466 18676 42476
rect 18732 42196 18788 44942
rect 20412 44546 20468 46508
rect 20972 46498 21028 46508
rect 21644 45220 21700 46622
rect 21644 45126 21700 45164
rect 23884 46676 23940 46686
rect 20412 44494 20414 44546
rect 20466 44494 20468 44546
rect 20412 44482 20468 44494
rect 23548 45106 23604 45118
rect 23548 45054 23550 45106
rect 23602 45054 23604 45106
rect 19292 44436 19348 44446
rect 18956 44434 19348 44436
rect 18956 44382 19294 44434
rect 19346 44382 19348 44434
rect 18956 44380 19348 44382
rect 18956 42308 19012 44380
rect 19292 44370 19348 44380
rect 21980 44436 22036 44446
rect 21980 44322 22036 44380
rect 21980 44270 21982 44322
rect 22034 44270 22036 44322
rect 21980 44258 22036 44270
rect 20300 44212 20356 44222
rect 20300 44118 20356 44156
rect 22316 44212 22372 44222
rect 22316 44118 22372 44156
rect 22988 44210 23044 44222
rect 22988 44158 22990 44210
rect 23042 44158 23044 44210
rect 21644 44100 21700 44110
rect 22204 44100 22260 44110
rect 21644 44006 21700 44044
rect 22092 44098 22260 44100
rect 22092 44046 22206 44098
rect 22258 44046 22260 44098
rect 22092 44044 22260 44046
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19068 43428 19124 43438
rect 19068 43426 20020 43428
rect 19068 43374 19070 43426
rect 19122 43374 20020 43426
rect 19068 43372 20020 43374
rect 19068 43362 19124 43372
rect 19964 42978 20020 43372
rect 21196 43426 21252 43438
rect 21196 43374 21198 43426
rect 21250 43374 21252 43426
rect 19964 42926 19966 42978
rect 20018 42926 20020 42978
rect 19964 42914 20020 42926
rect 20188 42980 20244 42990
rect 19180 42868 19236 42878
rect 19180 42774 19236 42812
rect 20076 42644 20132 42654
rect 20076 42550 20132 42588
rect 19068 42532 19124 42542
rect 19068 42438 19124 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 18956 42252 19236 42308
rect 19836 42298 20100 42308
rect 18732 42130 18788 42140
rect 18396 42028 18564 42084
rect 18956 42082 19012 42094
rect 18956 42030 18958 42082
rect 19010 42030 19012 42082
rect 18284 41972 18340 41982
rect 17388 41860 17444 41870
rect 17052 41858 17444 41860
rect 17052 41806 17390 41858
rect 17442 41806 17444 41858
rect 17052 41804 17444 41806
rect 16940 41794 16996 41804
rect 16716 41122 16772 41132
rect 17052 41186 17108 41198
rect 17052 41134 17054 41186
rect 17106 41134 17108 41186
rect 17052 41076 17108 41134
rect 17052 40964 17108 41020
rect 16380 39566 16382 39618
rect 16434 39566 16436 39618
rect 16380 39554 16436 39566
rect 16492 40908 17108 40964
rect 16492 39618 16548 40908
rect 16492 39566 16494 39618
rect 16546 39566 16548 39618
rect 16492 39554 16548 39566
rect 16604 40740 16660 40750
rect 16604 40402 16660 40684
rect 16604 40350 16606 40402
rect 16658 40350 16660 40402
rect 15932 39394 15988 39406
rect 15932 39342 15934 39394
rect 15986 39342 15988 39394
rect 15932 38612 15988 39342
rect 16156 38722 16212 39452
rect 16156 38670 16158 38722
rect 16210 38670 16212 38722
rect 16156 38668 16212 38670
rect 15932 38546 15988 38556
rect 16044 38612 16212 38668
rect 16380 38834 16436 38846
rect 16380 38782 16382 38834
rect 16434 38782 16436 38834
rect 15596 37986 15652 37996
rect 15708 38108 15876 38164
rect 15596 37380 15652 37390
rect 15484 37324 15596 37380
rect 15596 37314 15652 37324
rect 14924 37156 14980 37166
rect 14924 36706 14980 37100
rect 14924 36654 14926 36706
rect 14978 36654 14980 36706
rect 14924 36642 14980 36654
rect 15708 36708 15764 38108
rect 15932 38052 15988 38062
rect 15932 37958 15988 37996
rect 16044 38050 16100 38612
rect 16044 37998 16046 38050
rect 16098 37998 16100 38050
rect 16044 37986 16100 37998
rect 16380 38052 16436 38782
rect 16604 38668 16660 40350
rect 17388 40292 17444 41804
rect 17500 41860 17556 41870
rect 17500 40964 17556 41804
rect 17612 41748 17668 41758
rect 17612 41746 17780 41748
rect 17612 41694 17614 41746
rect 17666 41694 17780 41746
rect 17612 41692 17780 41694
rect 17612 41682 17668 41692
rect 17724 41298 17780 41692
rect 17724 41246 17726 41298
rect 17778 41246 17780 41298
rect 17724 41234 17780 41246
rect 17500 40898 17556 40908
rect 17612 41186 17668 41198
rect 17612 41134 17614 41186
rect 17666 41134 17668 41186
rect 17500 40740 17556 40750
rect 17500 40626 17556 40684
rect 17500 40574 17502 40626
rect 17554 40574 17556 40626
rect 17500 40562 17556 40574
rect 16828 40236 17444 40292
rect 17612 40404 17668 41134
rect 18172 41188 18228 41198
rect 18172 41094 18228 41132
rect 17948 40962 18004 40974
rect 17948 40910 17950 40962
rect 18002 40910 18004 40962
rect 17948 40740 18004 40910
rect 18284 40852 18340 41916
rect 18284 40786 18340 40796
rect 17948 40674 18004 40684
rect 18396 40628 18452 42028
rect 18956 41972 19012 42030
rect 18508 41916 19012 41972
rect 18508 41858 18564 41916
rect 18508 41806 18510 41858
rect 18562 41806 18564 41858
rect 18508 41524 18564 41806
rect 18620 41748 18676 41758
rect 18620 41654 18676 41692
rect 18508 41468 18788 41524
rect 18508 41074 18564 41086
rect 18508 41022 18510 41074
rect 18562 41022 18564 41074
rect 18508 40964 18564 41022
rect 18732 41076 18788 41468
rect 18732 40982 18788 41020
rect 18844 41300 18900 41310
rect 18844 41186 18900 41244
rect 18844 41134 18846 41186
rect 18898 41134 18900 41186
rect 18564 40908 18676 40964
rect 18508 40898 18564 40908
rect 18284 40572 18452 40628
rect 18620 40628 18676 40908
rect 17724 40404 17780 40414
rect 17612 40402 17780 40404
rect 17612 40350 17726 40402
rect 17778 40350 17780 40402
rect 17612 40348 17780 40350
rect 16716 39396 16772 39406
rect 16716 39302 16772 39340
rect 16604 38612 16772 38668
rect 16380 37986 16436 37996
rect 15820 37938 15876 37950
rect 15820 37886 15822 37938
rect 15874 37886 15876 37938
rect 15820 37716 15876 37886
rect 15820 37154 15876 37660
rect 16156 37828 16212 37838
rect 16492 37828 16548 37838
rect 16156 37378 16212 37772
rect 16156 37326 16158 37378
rect 16210 37326 16212 37378
rect 16156 37314 16212 37326
rect 16380 37826 16548 37828
rect 16380 37774 16494 37826
rect 16546 37774 16548 37826
rect 16380 37772 16548 37774
rect 16380 37378 16436 37772
rect 16492 37762 16548 37772
rect 16380 37326 16382 37378
rect 16434 37326 16436 37378
rect 15820 37102 15822 37154
rect 15874 37102 15876 37154
rect 15820 37090 15876 37102
rect 16268 37156 16324 37166
rect 16268 37062 16324 37100
rect 15708 36652 15988 36708
rect 14364 36484 14420 36494
rect 14700 36484 14756 36494
rect 14252 36482 14756 36484
rect 14252 36430 14366 36482
rect 14418 36430 14702 36482
rect 14754 36430 14756 36482
rect 14252 36428 14756 36430
rect 14140 35746 14196 35756
rect 13020 34962 13076 34972
rect 14252 35028 14308 35038
rect 14252 34934 14308 34972
rect 13468 34914 13524 34926
rect 13468 34862 13470 34914
rect 13522 34862 13524 34914
rect 13132 33348 13188 33358
rect 13020 33292 13132 33348
rect 13020 30996 13076 33292
rect 13132 33282 13188 33292
rect 13468 33348 13524 34862
rect 14252 34356 14308 34366
rect 14364 34356 14420 36428
rect 14700 36418 14756 36428
rect 15260 36484 15316 36494
rect 15820 36484 15876 36494
rect 15260 36482 15876 36484
rect 15260 36430 15262 36482
rect 15314 36430 15822 36482
rect 15874 36430 15876 36482
rect 15260 36428 15876 36430
rect 15260 36418 15316 36428
rect 15820 36418 15876 36428
rect 15596 36260 15652 36270
rect 15596 36166 15652 36204
rect 14812 35924 14868 35934
rect 15932 35924 15988 36652
rect 14812 35698 14868 35868
rect 15820 35868 15988 35924
rect 15260 35812 15316 35822
rect 15260 35718 15316 35756
rect 14812 35646 14814 35698
rect 14866 35646 14868 35698
rect 14812 35634 14868 35646
rect 14252 34354 14420 34356
rect 14252 34302 14254 34354
rect 14306 34302 14420 34354
rect 14252 34300 14420 34302
rect 14252 34290 14308 34300
rect 13468 33282 13524 33292
rect 14588 34130 14644 34142
rect 14588 34078 14590 34130
rect 14642 34078 14644 34130
rect 13804 33236 13860 33246
rect 13804 33142 13860 33180
rect 13468 33124 13524 33134
rect 13132 33122 13524 33124
rect 13132 33070 13470 33122
rect 13522 33070 13524 33122
rect 13132 33068 13524 33070
rect 13132 32674 13188 33068
rect 13468 33058 13524 33068
rect 14588 33012 14644 34078
rect 14588 32946 14644 32956
rect 15148 33346 15204 33358
rect 15148 33294 15150 33346
rect 15202 33294 15204 33346
rect 13132 32622 13134 32674
rect 13186 32622 13188 32674
rect 13132 32610 13188 32622
rect 15148 32452 15204 33294
rect 15708 33236 15764 33246
rect 15708 33142 15764 33180
rect 15372 33124 15428 33134
rect 15372 33030 15428 33068
rect 15708 32788 15764 32798
rect 15708 32694 15764 32732
rect 15260 32452 15316 32462
rect 15596 32452 15652 32462
rect 15148 32450 15652 32452
rect 15148 32398 15262 32450
rect 15314 32398 15598 32450
rect 15650 32398 15652 32450
rect 15148 32396 15652 32398
rect 15260 32386 15316 32396
rect 15596 32386 15652 32396
rect 15820 32116 15876 35868
rect 15932 35698 15988 35710
rect 15932 35646 15934 35698
rect 15986 35646 15988 35698
rect 15932 34132 15988 35646
rect 15932 34038 15988 34076
rect 16156 35588 16212 35598
rect 16380 35588 16436 37326
rect 16156 35586 16436 35588
rect 16156 35534 16158 35586
rect 16210 35534 16436 35586
rect 16156 35532 16436 35534
rect 16716 35924 16772 38612
rect 16828 36708 16884 40236
rect 17612 40180 17668 40348
rect 17724 40338 17780 40348
rect 18172 40402 18228 40414
rect 18172 40350 18174 40402
rect 18226 40350 18228 40402
rect 18060 40292 18116 40302
rect 16940 40124 17668 40180
rect 17948 40290 18116 40292
rect 17948 40238 18062 40290
rect 18114 40238 18116 40290
rect 17948 40236 18116 40238
rect 16940 39618 16996 40124
rect 17948 40068 18004 40236
rect 18060 40226 18116 40236
rect 18172 40180 18228 40350
rect 18172 40114 18228 40124
rect 17948 40002 18004 40012
rect 16940 39566 16942 39618
rect 16994 39566 16996 39618
rect 16940 39554 16996 39566
rect 17724 39956 17780 39966
rect 18284 39956 18340 40572
rect 17052 39508 17108 39518
rect 16940 38052 16996 38062
rect 16940 37958 16996 37996
rect 16828 36642 16884 36652
rect 16716 35588 16772 35868
rect 16716 35586 16884 35588
rect 16716 35534 16718 35586
rect 16770 35534 16884 35586
rect 16716 35532 16884 35534
rect 16156 34130 16212 35532
rect 16716 35522 16772 35532
rect 16156 34078 16158 34130
rect 16210 34078 16212 34130
rect 16156 34066 16212 34078
rect 16380 35026 16436 35038
rect 16380 34974 16382 35026
rect 16434 34974 16436 35026
rect 16380 34132 16436 34974
rect 16828 34916 16884 35532
rect 17052 35140 17108 39452
rect 17724 39508 17780 39900
rect 17724 39414 17780 39452
rect 18060 39900 18340 39956
rect 18396 40402 18452 40414
rect 18396 40350 18398 40402
rect 18450 40350 18452 40402
rect 17500 39396 17556 39406
rect 17500 39302 17556 39340
rect 17612 39394 17668 39406
rect 17612 39342 17614 39394
rect 17666 39342 17668 39394
rect 17612 39284 17668 39342
rect 17612 39218 17668 39228
rect 18060 38834 18116 39900
rect 18396 39508 18452 40350
rect 18620 39732 18676 40572
rect 18844 40404 18900 41134
rect 19068 40628 19124 42252
rect 19180 41970 19236 42252
rect 19180 41918 19182 41970
rect 19234 41918 19236 41970
rect 19180 41906 19236 41918
rect 20076 41858 20132 41870
rect 20076 41806 20078 41858
rect 20130 41806 20132 41858
rect 19292 41748 19348 41758
rect 19964 41748 20020 41758
rect 19348 41692 19572 41748
rect 19292 41682 19348 41692
rect 19516 41186 19572 41692
rect 19516 41134 19518 41186
rect 19570 41134 19572 41186
rect 19516 41122 19572 41134
rect 19628 41746 20020 41748
rect 19628 41694 19966 41746
rect 20018 41694 20020 41746
rect 19628 41692 20020 41694
rect 19628 40628 19684 41692
rect 19964 41682 20020 41692
rect 20076 41524 20132 41806
rect 19852 41468 20132 41524
rect 20188 41636 20244 42924
rect 21196 42868 21252 43374
rect 21532 43426 21588 43438
rect 21532 43374 21534 43426
rect 21586 43374 21588 43426
rect 21532 42980 21588 43374
rect 21532 42914 21588 42924
rect 21196 42802 21252 42812
rect 21868 42868 21924 42878
rect 21868 42754 21924 42812
rect 21868 42702 21870 42754
rect 21922 42702 21924 42754
rect 21868 42690 21924 42702
rect 21644 42530 21700 42542
rect 21644 42478 21646 42530
rect 21698 42478 21700 42530
rect 21644 42420 21700 42478
rect 21644 42354 21700 42364
rect 22092 42532 22148 44044
rect 22204 44034 22260 44044
rect 22428 44100 22484 44110
rect 22428 44006 22484 44044
rect 22540 44098 22596 44110
rect 22540 44046 22542 44098
rect 22594 44046 22596 44098
rect 22316 42756 22372 42766
rect 22204 42644 22260 42654
rect 22204 42550 22260 42588
rect 20188 41580 20916 41636
rect 19740 41076 19796 41086
rect 19852 41076 19908 41468
rect 19796 41020 19908 41076
rect 20076 41298 20132 41310
rect 20076 41246 20078 41298
rect 20130 41246 20132 41298
rect 19740 40982 19796 41020
rect 19964 40964 20020 41002
rect 20076 40964 20132 41246
rect 20188 41186 20244 41580
rect 20636 41300 20692 41310
rect 20636 41206 20692 41244
rect 20188 41134 20190 41186
rect 20242 41134 20244 41186
rect 20188 41122 20244 41134
rect 20524 41074 20580 41086
rect 20524 41022 20526 41074
rect 20578 41022 20580 41074
rect 20412 40964 20468 40974
rect 20524 40964 20580 41022
rect 20076 40908 20244 40964
rect 19964 40898 20020 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19852 40628 19908 40638
rect 19068 40572 19572 40628
rect 19628 40626 19908 40628
rect 19628 40574 19854 40626
rect 19906 40574 19908 40626
rect 19628 40572 19908 40574
rect 19516 40404 19572 40572
rect 19852 40562 19908 40572
rect 20076 40628 20132 40638
rect 20076 40534 20132 40572
rect 19628 40404 19684 40414
rect 19516 40402 19684 40404
rect 19516 40350 19630 40402
rect 19682 40350 19684 40402
rect 19516 40348 19684 40350
rect 18844 40338 18900 40348
rect 19628 40338 19684 40348
rect 19740 40404 19796 40414
rect 20188 40404 20244 40908
rect 20468 40908 20580 40964
rect 18732 39732 18788 39742
rect 18620 39730 18788 39732
rect 18620 39678 18734 39730
rect 18786 39678 18788 39730
rect 18620 39676 18788 39678
rect 18732 39666 18788 39676
rect 19628 39730 19684 39742
rect 19628 39678 19630 39730
rect 19682 39678 19684 39730
rect 19180 39620 19236 39630
rect 19516 39620 19572 39630
rect 19180 39618 19572 39620
rect 19180 39566 19182 39618
rect 19234 39566 19518 39618
rect 19570 39566 19572 39618
rect 19180 39564 19572 39566
rect 19180 39554 19236 39564
rect 19516 39554 19572 39564
rect 18620 39508 18676 39518
rect 18396 39452 18620 39508
rect 18620 39414 18676 39452
rect 19068 39506 19124 39518
rect 19068 39454 19070 39506
rect 19122 39454 19124 39506
rect 19068 39396 19124 39454
rect 19068 39330 19124 39340
rect 18060 38782 18062 38834
rect 18114 38782 18116 38834
rect 17836 38722 17892 38734
rect 17836 38670 17838 38722
rect 17890 38670 17892 38722
rect 17836 38668 17892 38670
rect 18060 38668 18116 38782
rect 17388 38612 17892 38668
rect 17948 38612 18116 38668
rect 18732 38722 18788 38734
rect 18732 38670 18734 38722
rect 18786 38670 18788 38722
rect 17164 38052 17220 38062
rect 17164 37958 17220 37996
rect 17276 37828 17332 37838
rect 17276 37734 17332 37772
rect 17388 37826 17444 38612
rect 17948 38276 18004 38612
rect 17612 38220 18004 38276
rect 18396 38610 18452 38622
rect 18396 38558 18398 38610
rect 18450 38558 18452 38610
rect 17612 38050 17668 38220
rect 18172 38164 18228 38174
rect 17612 37998 17614 38050
rect 17666 37998 17668 38050
rect 17612 37986 17668 37998
rect 17724 38052 17780 38062
rect 17388 37774 17390 37826
rect 17442 37774 17444 37826
rect 17388 37716 17444 37774
rect 17388 37650 17444 37660
rect 17388 37380 17444 37390
rect 17388 37286 17444 37324
rect 17612 37268 17668 37278
rect 17724 37268 17780 37996
rect 17948 38050 18004 38062
rect 18172 38052 18228 38108
rect 17948 37998 17950 38050
rect 18002 37998 18004 38050
rect 17948 37828 18004 37998
rect 17948 37762 18004 37772
rect 18060 38050 18228 38052
rect 18060 37998 18174 38050
rect 18226 37998 18228 38050
rect 18060 37996 18228 37998
rect 17948 37492 18004 37502
rect 18060 37492 18116 37996
rect 18172 37986 18228 37996
rect 17948 37490 18116 37492
rect 17948 37438 17950 37490
rect 18002 37438 18116 37490
rect 17948 37436 18116 37438
rect 18284 37940 18340 37950
rect 18396 37940 18452 38558
rect 18732 38164 18788 38670
rect 18844 38612 18900 38622
rect 18844 38610 19460 38612
rect 18844 38558 18846 38610
rect 18898 38558 19460 38610
rect 18844 38556 19460 38558
rect 18844 38546 18900 38556
rect 18732 38098 18788 38108
rect 18284 37938 18452 37940
rect 18284 37886 18286 37938
rect 18338 37886 18452 37938
rect 18284 37884 18452 37886
rect 18732 37940 18788 37950
rect 19068 37940 19124 37950
rect 18732 37938 19124 37940
rect 18732 37886 18734 37938
rect 18786 37886 19070 37938
rect 19122 37886 19124 37938
rect 18732 37884 19124 37886
rect 17948 37426 18004 37436
rect 17612 37266 17780 37268
rect 17612 37214 17614 37266
rect 17666 37214 17780 37266
rect 17612 37212 17780 37214
rect 18284 37268 18340 37884
rect 18732 37874 18788 37884
rect 19068 37874 19124 37884
rect 17612 37202 17668 37212
rect 18284 37202 18340 37212
rect 18508 37828 18564 37838
rect 18508 37266 18564 37772
rect 18956 37492 19012 37502
rect 18956 37398 19012 37436
rect 19180 37492 19236 37502
rect 19404 37492 19460 38556
rect 19180 37490 19460 37492
rect 19180 37438 19182 37490
rect 19234 37438 19460 37490
rect 19180 37436 19460 37438
rect 19516 38050 19572 38062
rect 19516 37998 19518 38050
rect 19570 37998 19572 38050
rect 19180 37426 19236 37436
rect 18508 37214 18510 37266
rect 18562 37214 18564 37266
rect 18508 37202 18564 37214
rect 19292 37268 19348 37278
rect 19068 37154 19124 37166
rect 19068 37102 19070 37154
rect 19122 37102 19124 37154
rect 19068 36820 19124 37102
rect 19068 36764 19236 36820
rect 17612 36708 17668 36718
rect 17612 36594 17668 36652
rect 17612 36542 17614 36594
rect 17666 36542 17668 36594
rect 17612 35476 17668 36542
rect 17836 36484 17892 36494
rect 17836 36482 18340 36484
rect 17836 36430 17838 36482
rect 17890 36430 18340 36482
rect 17836 36428 18340 36430
rect 17836 36418 17892 36428
rect 18172 36258 18228 36270
rect 18172 36206 18174 36258
rect 18226 36206 18228 36258
rect 17612 35410 17668 35420
rect 17724 35698 17780 35710
rect 17724 35646 17726 35698
rect 17778 35646 17780 35698
rect 17052 35074 17108 35084
rect 16940 34916 16996 34926
rect 16828 34860 16940 34916
rect 16940 34850 16996 34860
rect 17724 34244 17780 35646
rect 18172 35252 18228 36206
rect 18172 35186 18228 35196
rect 18060 35140 18116 35150
rect 17836 35028 17892 35038
rect 17836 34914 17892 34972
rect 17836 34862 17838 34914
rect 17890 34862 17892 34914
rect 17836 34850 17892 34862
rect 18060 34914 18116 35084
rect 18284 35026 18340 36428
rect 19180 36370 19236 36764
rect 19292 36482 19348 37212
rect 19292 36430 19294 36482
rect 19346 36430 19348 36482
rect 19292 36418 19348 36430
rect 19180 36318 19182 36370
rect 19234 36318 19236 36370
rect 19180 36306 19236 36318
rect 19516 36260 19572 37998
rect 19628 37492 19684 39678
rect 19740 39618 19796 40348
rect 20076 40348 20244 40404
rect 20300 40404 20356 40414
rect 19964 40292 20020 40302
rect 19964 40198 20020 40236
rect 19740 39566 19742 39618
rect 19794 39566 19796 39618
rect 19740 39554 19796 39566
rect 19964 39620 20020 39630
rect 20076 39620 20132 40348
rect 20300 40310 20356 40348
rect 20300 39844 20356 39854
rect 19964 39618 20076 39620
rect 19964 39566 19966 39618
rect 20018 39566 20076 39618
rect 19964 39564 20076 39566
rect 19964 39554 20020 39564
rect 20076 39526 20132 39564
rect 20188 39788 20300 39844
rect 20188 39618 20244 39788
rect 20300 39778 20356 39788
rect 20188 39566 20190 39618
rect 20242 39566 20244 39618
rect 20188 39554 20244 39566
rect 20188 39396 20244 39406
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20188 38388 20244 39340
rect 20300 38612 20356 38622
rect 20300 38518 20356 38556
rect 20188 38332 20356 38388
rect 20300 38162 20356 38332
rect 20300 38110 20302 38162
rect 20354 38110 20356 38162
rect 20300 38098 20356 38110
rect 20412 38050 20468 40908
rect 20524 40402 20580 40414
rect 20524 40350 20526 40402
rect 20578 40350 20580 40402
rect 20524 40292 20580 40350
rect 20524 39618 20580 40236
rect 20524 39566 20526 39618
rect 20578 39566 20580 39618
rect 20524 39554 20580 39566
rect 20636 39620 20692 39630
rect 20860 39620 20916 41580
rect 21308 41298 21364 41310
rect 21308 41246 21310 41298
rect 21362 41246 21364 41298
rect 21308 41076 21364 41246
rect 21308 40852 21364 41020
rect 22092 40964 22148 42476
rect 22316 42530 22372 42700
rect 22540 42754 22596 44046
rect 22540 42702 22542 42754
rect 22594 42702 22596 42754
rect 22540 42644 22596 42702
rect 22876 42980 22932 42990
rect 22876 42754 22932 42924
rect 22988 42868 23044 44158
rect 23100 44098 23156 44110
rect 23100 44046 23102 44098
rect 23154 44046 23156 44098
rect 23100 43652 23156 44046
rect 23100 43586 23156 43596
rect 23212 42868 23268 42878
rect 22988 42866 23268 42868
rect 22988 42814 23214 42866
rect 23266 42814 23268 42866
rect 22988 42812 23268 42814
rect 23212 42802 23268 42812
rect 22876 42702 22878 42754
rect 22930 42702 22932 42754
rect 22876 42690 22932 42702
rect 22540 42578 22596 42588
rect 22988 42644 23044 42654
rect 22316 42478 22318 42530
rect 22370 42478 22372 42530
rect 22316 42194 22372 42478
rect 22316 42142 22318 42194
rect 22370 42142 22372 42194
rect 22316 42130 22372 42142
rect 22540 41858 22596 41870
rect 22540 41806 22542 41858
rect 22594 41806 22596 41858
rect 22540 41076 22596 41806
rect 22652 41748 22708 41758
rect 22876 41748 22932 41758
rect 22652 41746 22932 41748
rect 22652 41694 22654 41746
rect 22706 41694 22878 41746
rect 22930 41694 22932 41746
rect 22652 41692 22932 41694
rect 22988 41748 23044 42588
rect 23436 42644 23492 42654
rect 23436 42550 23492 42588
rect 23100 42532 23156 42542
rect 23100 42438 23156 42476
rect 23324 42532 23380 42542
rect 23324 42438 23380 42476
rect 23548 42084 23604 45054
rect 23884 44324 23940 46620
rect 25228 46676 25284 46686
rect 25228 46582 25284 46620
rect 25004 46452 25060 46462
rect 24556 44436 24612 44446
rect 24556 44342 24612 44380
rect 23884 44322 24388 44324
rect 23884 44270 23886 44322
rect 23938 44270 24388 44322
rect 23884 44268 24388 44270
rect 23884 44258 23940 44268
rect 23660 43652 23716 43662
rect 23660 43558 23716 43596
rect 24332 43540 24388 44268
rect 23436 42028 23604 42084
rect 24108 43538 24388 43540
rect 24108 43486 24334 43538
rect 24386 43486 24388 43538
rect 24108 43484 24388 43486
rect 24108 42754 24164 43484
rect 24332 43474 24388 43484
rect 24108 42702 24110 42754
rect 24162 42702 24164 42754
rect 23100 41972 23156 41982
rect 23436 41972 23492 42028
rect 23100 41970 23436 41972
rect 23100 41918 23102 41970
rect 23154 41918 23436 41970
rect 23100 41916 23436 41918
rect 23100 41906 23156 41916
rect 23436 41878 23492 41916
rect 23548 41858 23604 41870
rect 23548 41806 23550 41858
rect 23602 41806 23604 41858
rect 22988 41692 23268 41748
rect 22652 41682 22708 41692
rect 22876 41682 22932 41692
rect 23100 41524 23156 41534
rect 22540 41020 23044 41076
rect 22092 40908 22596 40964
rect 21308 40786 21364 40796
rect 20972 40628 21028 40638
rect 21532 40628 21588 40638
rect 20972 40626 21588 40628
rect 20972 40574 20974 40626
rect 21026 40574 21534 40626
rect 21586 40574 21588 40626
rect 20972 40572 21588 40574
rect 20972 40562 21028 40572
rect 21196 40402 21252 40414
rect 21196 40350 21198 40402
rect 21250 40350 21252 40402
rect 21084 40290 21140 40302
rect 21084 40238 21086 40290
rect 21138 40238 21140 40290
rect 21084 39844 21140 40238
rect 21196 39956 21252 40350
rect 21196 39890 21252 39900
rect 21084 39778 21140 39788
rect 21308 39732 21364 40572
rect 21532 40562 21588 40572
rect 22092 40516 22148 40526
rect 21980 40404 22036 40414
rect 21980 40310 22036 40348
rect 21644 40290 21700 40302
rect 21644 40238 21646 40290
rect 21698 40238 21700 40290
rect 21196 39676 21364 39732
rect 21420 40180 21476 40190
rect 20860 39564 21028 39620
rect 20636 39506 20692 39564
rect 20636 39454 20638 39506
rect 20690 39454 20692 39506
rect 20636 39442 20692 39454
rect 20860 39396 20916 39406
rect 20748 39394 20916 39396
rect 20748 39342 20862 39394
rect 20914 39342 20916 39394
rect 20748 39340 20916 39342
rect 20748 38834 20804 39340
rect 20860 39330 20916 39340
rect 20972 39396 21028 39564
rect 20972 39330 21028 39340
rect 20748 38782 20750 38834
rect 20802 38782 20804 38834
rect 20748 38770 20804 38782
rect 20972 38834 21028 38846
rect 20972 38782 20974 38834
rect 21026 38782 21028 38834
rect 20412 37998 20414 38050
rect 20466 37998 20468 38050
rect 20412 37986 20468 37998
rect 20524 38612 20580 38622
rect 20076 37940 20132 37950
rect 20076 37846 20132 37884
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37426 19684 37436
rect 19740 37266 19796 37278
rect 19740 37214 19742 37266
rect 19794 37214 19796 37266
rect 19740 36594 19796 37214
rect 20524 37268 20580 38556
rect 20972 38164 21028 38782
rect 21196 38834 21252 39676
rect 21196 38782 21198 38834
rect 21250 38782 21252 38834
rect 21196 38770 21252 38782
rect 21420 39618 21476 40124
rect 21644 39730 21700 40238
rect 21644 39678 21646 39730
rect 21698 39678 21700 39730
rect 21644 39666 21700 39678
rect 21420 39566 21422 39618
rect 21474 39566 21476 39618
rect 21420 38668 21476 39566
rect 21868 39620 21924 39630
rect 22092 39620 22148 40460
rect 22428 40516 22484 40526
rect 21868 39618 22148 39620
rect 21868 39566 21870 39618
rect 21922 39566 22148 39618
rect 21868 39564 22148 39566
rect 22204 39956 22260 39966
rect 21868 39554 21924 39564
rect 21756 39508 21812 39518
rect 21756 39414 21812 39452
rect 21532 39396 21588 39406
rect 21532 39302 21588 39340
rect 22204 39060 22260 39900
rect 22428 39730 22484 40460
rect 22540 40292 22596 40908
rect 22652 40852 22708 40862
rect 22652 40514 22708 40796
rect 22988 40626 23044 41020
rect 22988 40574 22990 40626
rect 23042 40574 23044 40626
rect 22988 40562 23044 40574
rect 23100 40626 23156 41468
rect 23100 40574 23102 40626
rect 23154 40574 23156 40626
rect 23100 40562 23156 40574
rect 23212 40628 23268 41692
rect 23436 41746 23492 41758
rect 23436 41694 23438 41746
rect 23490 41694 23492 41746
rect 23436 41298 23492 41694
rect 23548 41748 23604 41806
rect 23548 41682 23604 41692
rect 24108 41860 24164 42702
rect 24556 43428 24612 43438
rect 24556 41970 24612 43372
rect 24780 42644 24836 42654
rect 24668 42642 24836 42644
rect 24668 42590 24782 42642
rect 24834 42590 24836 42642
rect 24668 42588 24836 42590
rect 24668 42194 24724 42588
rect 24780 42578 24836 42588
rect 24668 42142 24670 42194
rect 24722 42142 24724 42194
rect 24668 42130 24724 42142
rect 24556 41918 24558 41970
rect 24610 41918 24612 41970
rect 24556 41906 24612 41918
rect 24332 41860 24388 41870
rect 23436 41246 23438 41298
rect 23490 41246 23492 41298
rect 23436 41234 23492 41246
rect 24108 41188 24164 41804
rect 24108 41094 24164 41132
rect 24220 41858 24388 41860
rect 24220 41806 24334 41858
rect 24386 41806 24388 41858
rect 24220 41804 24388 41806
rect 23660 40628 23716 40638
rect 23212 40626 23716 40628
rect 23212 40574 23214 40626
rect 23266 40574 23662 40626
rect 23714 40574 23716 40626
rect 23212 40572 23716 40574
rect 23212 40562 23268 40572
rect 23660 40562 23716 40572
rect 23996 40628 24052 40638
rect 24220 40628 24276 41804
rect 24332 41794 24388 41804
rect 24780 41188 24836 41198
rect 24780 41094 24836 41132
rect 23996 40626 24388 40628
rect 23996 40574 23998 40626
rect 24050 40574 24388 40626
rect 23996 40572 24388 40574
rect 23996 40562 24052 40572
rect 22652 40462 22654 40514
rect 22706 40462 22708 40514
rect 22652 40450 22708 40462
rect 22876 40402 22932 40414
rect 22876 40350 22878 40402
rect 22930 40350 22932 40402
rect 22876 40292 22932 40350
rect 22540 40236 22932 40292
rect 22428 39678 22430 39730
rect 22482 39678 22484 39730
rect 22428 39666 22484 39678
rect 22092 39004 22260 39060
rect 22652 39396 22708 39406
rect 20972 38098 21028 38108
rect 21308 38612 21476 38668
rect 21644 38834 21700 38846
rect 21644 38782 21646 38834
rect 21698 38782 21700 38834
rect 20524 37202 20580 37212
rect 20748 37154 20804 37166
rect 20748 37102 20750 37154
rect 20802 37102 20804 37154
rect 19740 36542 19742 36594
rect 19794 36542 19796 36594
rect 19740 36530 19796 36542
rect 20076 37044 20132 37054
rect 20076 36482 20132 36988
rect 20636 37042 20692 37054
rect 20636 36990 20638 37042
rect 20690 36990 20692 37042
rect 20076 36430 20078 36482
rect 20130 36430 20132 36482
rect 20076 36260 20132 36430
rect 19516 36194 19572 36204
rect 19628 36204 20132 36260
rect 20524 36596 20580 36606
rect 18396 35586 18452 35598
rect 18396 35534 18398 35586
rect 18450 35534 18452 35586
rect 18396 35140 18452 35534
rect 18844 35252 18900 35262
rect 18396 35084 18676 35140
rect 18284 34974 18286 35026
rect 18338 34974 18340 35026
rect 18284 34962 18340 34974
rect 18060 34862 18062 34914
rect 18114 34862 18116 34914
rect 18060 34850 18116 34862
rect 18172 34916 18228 34926
rect 18060 34356 18116 34366
rect 18172 34356 18228 34860
rect 18620 34802 18676 35084
rect 18844 34914 18900 35196
rect 18844 34862 18846 34914
rect 18898 34862 18900 34914
rect 18844 34850 18900 34862
rect 18620 34750 18622 34802
rect 18674 34750 18676 34802
rect 18620 34738 18676 34750
rect 18060 34354 18228 34356
rect 18060 34302 18062 34354
rect 18114 34302 18228 34354
rect 18060 34300 18228 34302
rect 19628 34356 19684 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20524 35586 20580 36540
rect 20524 35534 20526 35586
rect 20578 35534 20580 35586
rect 20412 35028 20468 35038
rect 20412 34934 20468 34972
rect 20524 34914 20580 35534
rect 20524 34862 20526 34914
rect 20578 34862 20580 34914
rect 20524 34850 20580 34862
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19852 34356 19908 34366
rect 19628 34354 19908 34356
rect 19628 34302 19854 34354
rect 19906 34302 19908 34354
rect 19628 34300 19908 34302
rect 18060 34290 18116 34300
rect 19852 34290 19908 34300
rect 17724 34178 17780 34188
rect 16380 34066 16436 34076
rect 17388 34132 17444 34142
rect 17388 34038 17444 34076
rect 18620 34020 18676 34030
rect 18620 33926 18676 33964
rect 18844 34018 18900 34030
rect 18844 33966 18846 34018
rect 18898 33966 18900 34018
rect 16492 33908 16548 33918
rect 16492 33906 16772 33908
rect 16492 33854 16494 33906
rect 16546 33854 16772 33906
rect 16492 33852 16772 33854
rect 16492 33842 16548 33852
rect 16716 33684 16772 33852
rect 17500 33906 17556 33918
rect 17500 33854 17502 33906
rect 17554 33854 17556 33906
rect 16716 33628 16996 33684
rect 16940 33572 16996 33628
rect 17164 33572 17220 33582
rect 16940 33516 17164 33572
rect 17164 33478 17220 33516
rect 16828 33460 16884 33470
rect 16268 33458 16884 33460
rect 16268 33406 16830 33458
rect 16882 33406 16884 33458
rect 16268 33404 16884 33406
rect 16268 33346 16324 33404
rect 16828 33394 16884 33404
rect 16268 33294 16270 33346
rect 16322 33294 16324 33346
rect 16268 33282 16324 33294
rect 17500 33348 17556 33854
rect 17500 33282 17556 33292
rect 17836 33572 17892 33582
rect 18844 33572 18900 33966
rect 19292 34018 19348 34030
rect 19292 33966 19294 34018
rect 19346 33966 19348 34018
rect 18956 33908 19012 33918
rect 18956 33906 19236 33908
rect 18956 33854 18958 33906
rect 19010 33854 19236 33906
rect 18956 33852 19236 33854
rect 18956 33842 19012 33852
rect 18844 33516 19012 33572
rect 16156 33236 16212 33246
rect 16156 33142 16212 33180
rect 16380 33234 16436 33246
rect 16380 33182 16382 33234
rect 16434 33182 16436 33234
rect 16380 33124 16436 33182
rect 17388 33234 17444 33246
rect 17388 33182 17390 33234
rect 17442 33182 17444 33234
rect 17388 33124 17444 33182
rect 16380 33068 16772 33124
rect 16380 33012 16436 33068
rect 16380 32946 16436 32956
rect 16492 32564 16548 32574
rect 16268 32562 16548 32564
rect 16268 32510 16494 32562
rect 16546 32510 16548 32562
rect 16268 32508 16548 32510
rect 15596 32060 15876 32116
rect 16044 32338 16100 32350
rect 16044 32286 16046 32338
rect 16098 32286 16100 32338
rect 13580 31780 13636 31790
rect 13580 31686 13636 31724
rect 13468 30996 13524 31006
rect 13076 30994 13972 30996
rect 13076 30942 13470 30994
rect 13522 30942 13972 30994
rect 13076 30940 13972 30942
rect 13020 30902 13076 30940
rect 13468 30930 13524 30940
rect 13804 30772 13860 30782
rect 13804 30210 13860 30716
rect 13804 30158 13806 30210
rect 13858 30158 13860 30210
rect 13804 30146 13860 30158
rect 13916 30324 13972 30940
rect 14252 30884 14308 30894
rect 13916 29426 13972 30268
rect 14140 30882 14308 30884
rect 14140 30830 14254 30882
rect 14306 30830 14308 30882
rect 14140 30828 14308 30830
rect 14140 30098 14196 30828
rect 14252 30818 14308 30828
rect 14476 30548 14532 30558
rect 14532 30492 14644 30548
rect 14476 30482 14532 30492
rect 14140 30046 14142 30098
rect 14194 30046 14196 30098
rect 14140 30034 14196 30046
rect 14476 30210 14532 30222
rect 14476 30158 14478 30210
rect 14530 30158 14532 30210
rect 13916 29374 13918 29426
rect 13970 29374 13972 29426
rect 13916 29362 13972 29374
rect 14476 29316 14532 30158
rect 14476 29250 14532 29260
rect 14028 28756 14084 28766
rect 13468 28084 13524 28094
rect 13132 27748 13188 27758
rect 12908 26852 13076 26908
rect 9212 26226 9268 26236
rect 9548 26292 9604 26302
rect 9548 26198 9604 26236
rect 12460 26292 12516 26302
rect 10332 26180 10388 26190
rect 8652 26178 9044 26180
rect 8652 26126 8990 26178
rect 9042 26126 9044 26178
rect 8652 26124 9044 26126
rect 7980 25454 7982 25506
rect 8034 25454 8036 25506
rect 7980 25442 8036 25454
rect 8428 25508 8484 25518
rect 8428 25414 8484 25452
rect 8652 25506 8708 26124
rect 8988 26114 9044 26124
rect 10108 26178 10388 26180
rect 10108 26126 10334 26178
rect 10386 26126 10388 26178
rect 10108 26124 10388 26126
rect 8652 25454 8654 25506
rect 8706 25454 8708 25506
rect 8652 25442 8708 25454
rect 9772 25508 9828 25518
rect 9772 25414 9828 25452
rect 8316 25396 8372 25406
rect 8316 25302 8372 25340
rect 10108 25394 10164 26124
rect 10332 26114 10388 26124
rect 12460 26178 12516 26236
rect 12460 26126 12462 26178
rect 12514 26126 12516 26178
rect 12460 26114 12516 26126
rect 12684 26068 12740 26078
rect 12572 26066 12740 26068
rect 12572 26014 12686 26066
rect 12738 26014 12740 26066
rect 12572 26012 12740 26014
rect 10444 25508 10500 25518
rect 10444 25414 10500 25452
rect 10780 25508 10836 25518
rect 10780 25414 10836 25452
rect 11004 25506 11060 25518
rect 11004 25454 11006 25506
rect 11058 25454 11060 25506
rect 10108 25342 10110 25394
rect 10162 25342 10164 25394
rect 10108 25330 10164 25342
rect 7868 25228 8260 25284
rect 7644 24836 7700 24846
rect 6636 24670 6638 24722
rect 6690 24670 6692 24722
rect 6636 24658 6692 24670
rect 6860 24834 7700 24836
rect 6860 24782 7646 24834
rect 7698 24782 7700 24834
rect 6860 24780 7700 24782
rect 6188 24612 6244 24622
rect 6188 24518 6244 24556
rect 6524 24500 6580 24510
rect 6412 24498 6580 24500
rect 6412 24446 6526 24498
rect 6578 24446 6580 24498
rect 6412 24444 6580 24446
rect 6412 24164 6468 24444
rect 6524 24434 6580 24444
rect 5404 24098 5460 24108
rect 6076 24108 6468 24164
rect 5964 24052 6020 24062
rect 5628 23940 5684 23950
rect 5628 23846 5684 23884
rect 5852 23826 5908 23838
rect 5852 23774 5854 23826
rect 5906 23774 5908 23826
rect 5852 23492 5908 23774
rect 5292 23436 5460 23492
rect 4620 23156 4676 23166
rect 4508 23154 4676 23156
rect 4508 23102 4622 23154
rect 4674 23102 4676 23154
rect 4508 23100 4676 23102
rect 4620 23090 4676 23100
rect 4844 23156 4900 23212
rect 5068 23156 5124 23166
rect 4844 23154 5124 23156
rect 4844 23102 4846 23154
rect 4898 23102 5070 23154
rect 5122 23102 5124 23154
rect 4844 23100 5124 23102
rect 4844 23090 4900 23100
rect 5068 23090 5124 23100
rect 5292 23156 5348 23166
rect 5292 23062 5348 23100
rect 5404 23156 5460 23436
rect 5628 23436 5908 23492
rect 5628 23156 5684 23436
rect 5740 23268 5796 23278
rect 5964 23268 6020 23996
rect 6076 24050 6132 24108
rect 6076 23998 6078 24050
rect 6130 23998 6132 24050
rect 6076 23986 6132 23998
rect 6636 24052 6692 24062
rect 6636 23958 6692 23996
rect 6300 23940 6356 23950
rect 6188 23828 6244 23838
rect 6188 23734 6244 23772
rect 5740 23266 6020 23268
rect 5740 23214 5742 23266
rect 5794 23214 6020 23266
rect 5740 23212 6020 23214
rect 5740 23202 5796 23212
rect 5404 23154 5684 23156
rect 5404 23102 5406 23154
rect 5458 23102 5684 23154
rect 5404 23100 5684 23102
rect 6188 23156 6244 23166
rect 6300 23156 6356 23884
rect 6860 23266 6916 24780
rect 7644 24770 7700 24780
rect 7868 24052 7924 25228
rect 8204 25172 8260 25228
rect 8204 25116 8484 25172
rect 8428 24946 8484 25116
rect 8428 24894 8430 24946
rect 8482 24894 8484 24946
rect 8428 24882 8484 24894
rect 9996 24834 10052 24846
rect 9996 24782 9998 24834
rect 10050 24782 10052 24834
rect 7980 24724 8036 24734
rect 7980 24722 8260 24724
rect 7980 24670 7982 24722
rect 8034 24670 8260 24722
rect 7980 24668 8260 24670
rect 7980 24658 8036 24668
rect 7868 23958 7924 23996
rect 8204 24050 8260 24668
rect 8204 23998 8206 24050
rect 8258 23998 8260 24050
rect 8204 23986 8260 23998
rect 9884 24052 9940 24062
rect 9996 24052 10052 24782
rect 10332 24724 10388 24734
rect 10332 24722 10500 24724
rect 10332 24670 10334 24722
rect 10386 24670 10500 24722
rect 10332 24668 10500 24670
rect 10332 24658 10388 24668
rect 9884 24050 10052 24052
rect 9884 23998 9886 24050
rect 9938 23998 10052 24050
rect 9884 23996 10052 23998
rect 9884 23986 9940 23996
rect 7756 23938 7812 23950
rect 7756 23886 7758 23938
rect 7810 23886 7812 23938
rect 7756 23828 7812 23886
rect 7756 23762 7812 23772
rect 9100 23940 9156 23950
rect 6860 23214 6862 23266
rect 6914 23214 6916 23266
rect 6860 23202 6916 23214
rect 8764 23716 8820 23726
rect 6188 23154 6356 23156
rect 6188 23102 6190 23154
rect 6242 23102 6356 23154
rect 6188 23100 6356 23102
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 3612 22530 3668 22540
rect 4620 22596 4676 22606
rect 4620 22482 4676 22540
rect 5404 22596 5460 23100
rect 5404 22530 5460 22540
rect 4620 22430 4622 22482
rect 4674 22430 4676 22482
rect 4620 22418 4676 22430
rect 2828 21646 2830 21698
rect 2882 21646 2884 21698
rect 2828 21634 2884 21646
rect 3948 21812 4004 21822
rect 1820 20710 1876 20748
rect 3948 20804 4004 21756
rect 5516 21812 5572 21822
rect 5516 21586 5572 21756
rect 6188 21812 6244 23100
rect 8764 23044 8820 23660
rect 8988 23044 9044 23054
rect 8764 23042 9044 23044
rect 8764 22990 8990 23042
rect 9042 22990 9044 23042
rect 8764 22988 9044 22990
rect 8988 22708 9044 22988
rect 8988 22642 9044 22652
rect 9100 22482 9156 23884
rect 10444 23378 10500 24668
rect 10444 23326 10446 23378
rect 10498 23326 10500 23378
rect 10444 23314 10500 23326
rect 10780 24612 10836 24622
rect 10780 23154 10836 24556
rect 10780 23102 10782 23154
rect 10834 23102 10836 23154
rect 10780 23090 10836 23102
rect 11004 24052 11060 25454
rect 12236 25508 12292 25518
rect 12236 25414 12292 25452
rect 12460 25508 12516 25518
rect 12460 25414 12516 25452
rect 12124 25396 12180 25406
rect 12012 25394 12180 25396
rect 12012 25342 12126 25394
rect 12178 25342 12180 25394
rect 12012 25340 12180 25342
rect 11900 24612 11956 24622
rect 11900 24518 11956 24556
rect 11004 23156 11060 23996
rect 11676 24500 11732 24510
rect 11676 23266 11732 24444
rect 11788 24498 11844 24510
rect 11788 24446 11790 24498
rect 11842 24446 11844 24498
rect 11788 23378 11844 24446
rect 12012 24500 12068 25340
rect 12124 25330 12180 25340
rect 12012 24434 12068 24444
rect 12124 24722 12180 24734
rect 12124 24670 12126 24722
rect 12178 24670 12180 24722
rect 12124 24276 12180 24670
rect 12572 24722 12628 26012
rect 12684 26002 12740 26012
rect 12572 24670 12574 24722
rect 12626 24670 12628 24722
rect 12012 24050 12068 24062
rect 12012 23998 12014 24050
rect 12066 23998 12068 24050
rect 12012 23940 12068 23998
rect 12012 23874 12068 23884
rect 11788 23326 11790 23378
rect 11842 23326 11844 23378
rect 11788 23314 11844 23326
rect 11676 23214 11678 23266
rect 11730 23214 11732 23266
rect 11676 23202 11732 23214
rect 12012 23268 12068 23278
rect 12012 23174 12068 23212
rect 11004 23154 11508 23156
rect 11004 23102 11006 23154
rect 11058 23102 11508 23154
rect 11004 23100 11508 23102
rect 11004 23090 11060 23100
rect 9100 22430 9102 22482
rect 9154 22430 9156 22482
rect 9100 22418 9156 22430
rect 11004 22708 11060 22718
rect 6636 22372 6692 22382
rect 6636 22278 6692 22316
rect 10332 22372 10388 22382
rect 6188 21746 6244 21756
rect 6748 21812 6804 21822
rect 8764 21812 8820 21822
rect 5516 21534 5518 21586
rect 5570 21534 5572 21586
rect 5516 21522 5572 21534
rect 6188 21474 6244 21486
rect 6188 21422 6190 21474
rect 6242 21422 6244 21474
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 2492 20692 2548 20702
rect 2492 20690 3108 20692
rect 2492 20638 2494 20690
rect 2546 20638 3108 20690
rect 2492 20636 3108 20638
rect 2492 20626 2548 20636
rect 3052 20242 3108 20636
rect 3052 20190 3054 20242
rect 3106 20190 3108 20242
rect 3052 20178 3108 20190
rect 2492 20132 2548 20142
rect 2492 20038 2548 20076
rect 2716 20132 2772 20142
rect 2716 20130 2884 20132
rect 2716 20078 2718 20130
rect 2770 20078 2884 20130
rect 2716 20076 2884 20078
rect 2716 20066 2772 20076
rect 2380 20018 2436 20030
rect 2380 19966 2382 20018
rect 2434 19966 2436 20018
rect 2380 19684 2436 19966
rect 2828 20018 2884 20076
rect 2828 19966 2830 20018
rect 2882 19966 2884 20018
rect 2828 19954 2884 19966
rect 3164 20018 3220 20030
rect 3164 19966 3166 20018
rect 3218 19966 3220 20018
rect 2380 19628 2884 19684
rect 1820 19234 1876 19246
rect 1820 19182 1822 19234
rect 1874 19182 1876 19234
rect 1708 18116 1764 18126
rect 1708 16994 1764 18060
rect 1708 16942 1710 16994
rect 1762 16942 1764 16994
rect 1708 16930 1764 16942
rect 1820 17666 1876 19182
rect 2492 19124 2548 19134
rect 2492 19122 2772 19124
rect 2492 19070 2494 19122
rect 2546 19070 2772 19122
rect 2492 19068 2772 19070
rect 2492 19058 2548 19068
rect 2604 18676 2660 18686
rect 2492 18562 2548 18574
rect 2492 18510 2494 18562
rect 2546 18510 2548 18562
rect 2268 18452 2324 18462
rect 2268 18358 2324 18396
rect 2492 17780 2548 18510
rect 2604 18562 2660 18620
rect 2604 18510 2606 18562
rect 2658 18510 2660 18562
rect 2604 17780 2660 18510
rect 2716 18340 2772 19068
rect 2828 18564 2884 19628
rect 2940 18564 2996 18574
rect 2828 18562 2996 18564
rect 2828 18510 2942 18562
rect 2994 18510 2996 18562
rect 2828 18508 2996 18510
rect 2716 18274 2772 18284
rect 2940 17892 2996 18508
rect 3052 18564 3108 18574
rect 3052 18470 3108 18508
rect 3164 18228 3220 19966
rect 3500 20018 3556 20030
rect 3500 19966 3502 20018
rect 3554 19966 3556 20018
rect 3276 18562 3332 18574
rect 3276 18510 3278 18562
rect 3330 18510 3332 18562
rect 3276 18452 3332 18510
rect 3388 18452 3444 18462
rect 3276 18450 3444 18452
rect 3276 18398 3390 18450
rect 3442 18398 3444 18450
rect 3276 18396 3444 18398
rect 3388 18386 3444 18396
rect 3164 18162 3220 18172
rect 3500 18116 3556 19966
rect 3948 20018 4004 20748
rect 4620 20914 4676 20926
rect 4620 20862 4622 20914
rect 4674 20862 4676 20914
rect 4620 20132 4676 20862
rect 5852 20690 5908 20702
rect 5852 20638 5854 20690
rect 5906 20638 5908 20690
rect 4620 20066 4676 20076
rect 5068 20132 5124 20142
rect 3948 19966 3950 20018
rect 4002 19966 4004 20018
rect 3948 19954 4004 19966
rect 4620 19908 4676 19918
rect 4620 19814 4676 19852
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4620 19348 4676 19358
rect 4508 19346 4676 19348
rect 4508 19294 4622 19346
rect 4674 19294 4676 19346
rect 4508 19292 4676 19294
rect 4284 18564 4340 18574
rect 3724 18452 3780 18462
rect 3724 18358 3780 18396
rect 3948 18452 4004 18462
rect 3612 18340 3668 18350
rect 3612 18246 3668 18284
rect 3500 18050 3556 18060
rect 3948 18116 4004 18396
rect 3948 18050 4004 18060
rect 4284 18452 4340 18508
rect 4508 18562 4564 19292
rect 4620 19282 4676 19292
rect 4508 18510 4510 18562
rect 4562 18510 4564 18562
rect 4508 18452 4564 18510
rect 4620 18676 4676 18686
rect 4620 18564 4676 18620
rect 5068 18674 5124 20076
rect 5852 19348 5908 20638
rect 6076 20690 6132 20702
rect 6076 20638 6078 20690
rect 6130 20638 6132 20690
rect 5068 18622 5070 18674
rect 5122 18622 5124 18674
rect 5068 18610 5124 18622
rect 5292 19292 5796 19348
rect 5292 18674 5348 19292
rect 5628 19124 5684 19134
rect 5292 18622 5294 18674
rect 5346 18622 5348 18674
rect 5292 18610 5348 18622
rect 5516 19122 5684 19124
rect 5516 19070 5630 19122
rect 5682 19070 5684 19122
rect 5516 19068 5684 19070
rect 5740 19124 5796 19292
rect 5852 19282 5908 19292
rect 5964 19908 6020 19918
rect 5852 19124 5908 19134
rect 5740 19122 5908 19124
rect 5740 19070 5854 19122
rect 5906 19070 5908 19122
rect 5740 19068 5908 19070
rect 4956 18564 5012 18574
rect 4620 18562 5012 18564
rect 4620 18510 4622 18562
rect 4674 18510 4958 18562
rect 5010 18510 5012 18562
rect 4620 18508 5012 18510
rect 4620 18498 4676 18508
rect 4956 18498 5012 18508
rect 5516 18562 5572 19068
rect 5628 19058 5684 19068
rect 5852 19058 5908 19068
rect 5964 19010 6020 19852
rect 6076 19236 6132 20638
rect 6188 20578 6244 21422
rect 6524 21364 6580 21374
rect 6524 20802 6580 21308
rect 6524 20750 6526 20802
rect 6578 20750 6580 20802
rect 6524 20738 6580 20750
rect 6748 20802 6804 21756
rect 8428 21756 8764 21812
rect 8316 21476 8372 21486
rect 8428 21476 8484 21756
rect 8764 21718 8820 21756
rect 9660 21812 9716 21822
rect 9660 21718 9716 21756
rect 10220 21700 10276 21710
rect 10220 21606 10276 21644
rect 8316 21474 8484 21476
rect 8316 21422 8318 21474
rect 8370 21422 8484 21474
rect 8316 21420 8484 21422
rect 8316 21410 8372 21420
rect 6748 20750 6750 20802
rect 6802 20750 6804 20802
rect 6748 20738 6804 20750
rect 6188 20526 6190 20578
rect 6242 20526 6244 20578
rect 6188 20514 6244 20526
rect 7532 20690 7588 20702
rect 7532 20638 7534 20690
rect 7586 20638 7588 20690
rect 7420 20132 7476 20142
rect 7420 20038 7476 20076
rect 7308 20020 7364 20030
rect 6748 20018 7364 20020
rect 6748 19966 7310 20018
rect 7362 19966 7364 20018
rect 6748 19964 7364 19966
rect 6748 19908 6804 19964
rect 6076 19170 6132 19180
rect 6636 19906 6804 19908
rect 6636 19854 6750 19906
rect 6802 19854 6804 19906
rect 6636 19852 6804 19854
rect 6188 19124 6244 19134
rect 6412 19124 6468 19134
rect 6188 19122 6468 19124
rect 6188 19070 6190 19122
rect 6242 19070 6414 19122
rect 6466 19070 6468 19122
rect 6188 19068 6468 19070
rect 6188 19058 6244 19068
rect 6412 19058 6468 19068
rect 6636 19122 6692 19852
rect 6748 19842 6804 19852
rect 7308 19460 7364 19964
rect 7532 19796 7588 20638
rect 8316 20244 8372 20282
rect 8316 20178 8372 20188
rect 8428 20018 8484 21420
rect 8428 19966 8430 20018
rect 8482 19966 8484 20018
rect 8428 19954 8484 19966
rect 8540 21586 8596 21598
rect 8540 21534 8542 21586
rect 8594 21534 8596 21586
rect 7532 19730 7588 19740
rect 7308 19404 7700 19460
rect 7420 19236 7476 19246
rect 7420 19142 7476 19180
rect 6636 19070 6638 19122
rect 6690 19070 6692 19122
rect 6636 19058 6692 19070
rect 6748 19124 6804 19134
rect 5964 18958 5966 19010
rect 6018 18958 6020 19010
rect 5964 18946 6020 18958
rect 6636 18676 6692 18686
rect 6748 18676 6804 19068
rect 7644 19122 7700 19404
rect 8316 19348 8372 19358
rect 8316 19234 8372 19292
rect 8316 19182 8318 19234
rect 8370 19182 8372 19234
rect 7644 19070 7646 19122
rect 7698 19070 7700 19122
rect 7644 19058 7700 19070
rect 7756 19122 7812 19134
rect 7756 19070 7758 19122
rect 7810 19070 7812 19122
rect 6636 18674 6804 18676
rect 6636 18622 6638 18674
rect 6690 18622 6804 18674
rect 6636 18620 6804 18622
rect 6636 18610 6692 18620
rect 5516 18510 5518 18562
rect 5570 18510 5572 18562
rect 4284 18396 4564 18452
rect 5516 18452 5572 18510
rect 7756 18562 7812 19070
rect 7756 18510 7758 18562
rect 7810 18510 7812 18562
rect 2940 17836 3108 17892
rect 2604 17724 2996 17780
rect 2492 17714 2548 17724
rect 1820 17614 1822 17666
rect 1874 17614 1876 17666
rect 1820 16996 1876 17614
rect 2492 17554 2548 17566
rect 2492 17502 2494 17554
rect 2546 17502 2548 17554
rect 2268 16996 2324 17006
rect 1820 16098 1876 16940
rect 2044 16994 2324 16996
rect 2044 16942 2270 16994
rect 2322 16942 2324 16994
rect 2044 16940 2324 16942
rect 1820 16046 1822 16098
rect 1874 16046 1876 16098
rect 1820 14530 1876 16046
rect 1932 16882 1988 16894
rect 1932 16830 1934 16882
rect 1986 16830 1988 16882
rect 1932 15204 1988 16830
rect 2044 15538 2100 16940
rect 2268 16930 2324 16940
rect 2156 16772 2212 16782
rect 2492 16772 2548 17502
rect 2828 16996 2884 17006
rect 2828 16902 2884 16940
rect 2156 16770 2548 16772
rect 2156 16718 2158 16770
rect 2210 16718 2548 16770
rect 2156 16716 2548 16718
rect 2604 16772 2660 16782
rect 2156 16706 2212 16716
rect 2604 16660 2660 16716
rect 2380 16604 2660 16660
rect 2044 15486 2046 15538
rect 2098 15486 2100 15538
rect 2044 15474 2100 15486
rect 2268 15540 2324 15550
rect 2268 15446 2324 15484
rect 2380 15426 2436 16604
rect 2492 15988 2548 15998
rect 2492 15894 2548 15932
rect 2380 15374 2382 15426
rect 2434 15374 2436 15426
rect 2380 15362 2436 15374
rect 2828 15428 2884 15438
rect 2828 15334 2884 15372
rect 2604 15314 2660 15326
rect 2604 15262 2606 15314
rect 2658 15262 2660 15314
rect 2604 15204 2660 15262
rect 1932 15148 2660 15204
rect 2940 15314 2996 17724
rect 3052 16772 3108 17836
rect 3052 16706 3108 16716
rect 4172 17780 4228 17790
rect 3388 15988 3444 15998
rect 3388 15538 3444 15932
rect 3388 15486 3390 15538
rect 3442 15486 3444 15538
rect 3388 15474 3444 15486
rect 4172 15540 4228 17724
rect 2940 15262 2942 15314
rect 2994 15262 2996 15314
rect 1820 14478 1822 14530
rect 1874 14478 1876 14530
rect 1820 14466 1876 14478
rect 2492 14418 2548 14430
rect 2492 14366 2494 14418
rect 2546 14366 2548 14418
rect 2492 13860 2548 14366
rect 2940 14308 2996 15262
rect 3276 15316 3332 15326
rect 3276 15222 3332 15260
rect 3612 15314 3668 15326
rect 3612 15262 3614 15314
rect 3666 15262 3668 15314
rect 3612 14756 3668 15262
rect 3836 15314 3892 15326
rect 3836 15262 3838 15314
rect 3890 15262 3892 15314
rect 3836 15204 3892 15262
rect 4172 15314 4228 15484
rect 4284 15426 4340 18396
rect 5516 18386 5572 18396
rect 5852 18450 5908 18462
rect 6860 18452 6916 18462
rect 5852 18398 5854 18450
rect 5906 18398 5908 18450
rect 4508 18228 4564 18266
rect 4508 18162 4564 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4620 17780 4676 17790
rect 4620 17686 4676 17724
rect 5852 16884 5908 18398
rect 6300 18450 6916 18452
rect 6300 18398 6862 18450
rect 6914 18398 6916 18450
rect 6300 18396 6916 18398
rect 6300 17668 6356 18396
rect 6860 18386 6916 18396
rect 7420 18450 7476 18462
rect 7420 18398 7422 18450
rect 7474 18398 7476 18450
rect 6300 17574 6356 17612
rect 6860 17554 6916 17566
rect 6860 17502 6862 17554
rect 6914 17502 6916 17554
rect 5852 16818 5908 16828
rect 5964 17442 6020 17454
rect 5964 17390 5966 17442
rect 6018 17390 6020 17442
rect 5964 16772 6020 17390
rect 6524 17444 6580 17454
rect 6524 17350 6580 17388
rect 6748 17442 6804 17454
rect 6748 17390 6750 17442
rect 6802 17390 6804 17442
rect 5964 16706 6020 16716
rect 6524 16884 6580 16894
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4284 15374 4286 15426
rect 4338 15374 4340 15426
rect 4284 15362 4340 15374
rect 4620 16210 4676 16222
rect 4620 16158 4622 16210
rect 4674 16158 4676 16210
rect 4620 15428 4676 16158
rect 5964 16210 6020 16222
rect 5964 16158 5966 16210
rect 6018 16158 6020 16210
rect 4620 15362 4676 15372
rect 5628 15538 5684 15550
rect 5628 15486 5630 15538
rect 5682 15486 5684 15538
rect 4172 15262 4174 15314
rect 4226 15262 4228 15314
rect 4172 15250 4228 15262
rect 3836 15138 3892 15148
rect 4844 15204 4900 15214
rect 4900 15148 5012 15204
rect 4844 15138 4900 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4844 14868 4900 14878
rect 3612 14690 3668 14700
rect 2940 14242 2996 14252
rect 4620 14644 4676 14654
rect 4844 14644 4900 14812
rect 4620 14642 4900 14644
rect 4620 14590 4622 14642
rect 4674 14590 4900 14642
rect 4620 14588 4900 14590
rect 3724 14028 4564 14084
rect 2492 13794 2548 13804
rect 3164 13972 3220 13982
rect 3164 13858 3220 13916
rect 3500 13972 3556 13982
rect 3724 13972 3780 14028
rect 3500 13970 3780 13972
rect 3500 13918 3502 13970
rect 3554 13918 3780 13970
rect 3500 13916 3780 13918
rect 3500 13906 3556 13916
rect 3164 13806 3166 13858
rect 3218 13806 3220 13858
rect 3164 13794 3220 13806
rect 3276 13858 3332 13870
rect 3276 13806 3278 13858
rect 3330 13806 3332 13858
rect 3276 13188 3332 13806
rect 3836 13858 3892 13870
rect 3836 13806 3838 13858
rect 3890 13806 3892 13858
rect 3724 13746 3780 13758
rect 3724 13694 3726 13746
rect 3778 13694 3780 13746
rect 3724 13636 3780 13694
rect 3836 13748 3892 13806
rect 4060 13860 4116 13870
rect 4396 13860 4452 13870
rect 4060 13858 4228 13860
rect 4060 13806 4062 13858
rect 4114 13806 4228 13858
rect 4060 13804 4228 13806
rect 4060 13794 4116 13804
rect 3836 13682 3892 13692
rect 4172 13746 4228 13804
rect 4396 13766 4452 13804
rect 4172 13694 4174 13746
rect 4226 13694 4228 13746
rect 4172 13682 4228 13694
rect 4508 13746 4564 14028
rect 4508 13694 4510 13746
rect 4562 13694 4564 13746
rect 4508 13682 4564 13694
rect 4620 13748 4676 14588
rect 4844 13860 4900 13870
rect 4956 13860 5012 15148
rect 5628 14532 5684 15486
rect 5964 15540 6020 16158
rect 5964 15474 6020 15484
rect 6412 16100 6468 16110
rect 5740 15426 5796 15438
rect 5740 15374 5742 15426
rect 5794 15374 5796 15426
rect 5740 14868 5796 15374
rect 5852 15428 5908 15438
rect 5852 15314 5908 15372
rect 5852 15262 5854 15314
rect 5906 15262 5908 15314
rect 5852 15250 5908 15262
rect 6188 15426 6244 15438
rect 6188 15374 6190 15426
rect 6242 15374 6244 15426
rect 6188 15204 6244 15374
rect 6188 15138 6244 15148
rect 5740 14802 5796 14812
rect 5628 14476 6244 14532
rect 5628 14308 5684 14318
rect 5628 14214 5684 14252
rect 5964 14306 6020 14318
rect 5964 14254 5966 14306
rect 6018 14254 6020 14306
rect 4844 13858 5012 13860
rect 4844 13806 4846 13858
rect 4898 13806 5012 13858
rect 4844 13804 5012 13806
rect 4844 13794 4900 13804
rect 4620 13682 4676 13692
rect 3276 13122 3332 13132
rect 3388 13580 3724 13636
rect 2492 13076 2548 13086
rect 2492 12982 2548 13020
rect 1820 12962 1876 12974
rect 1820 12910 1822 12962
rect 1874 12910 1876 12962
rect 1820 11508 1876 12910
rect 3388 12290 3444 13580
rect 3724 13570 3780 13580
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4620 13188 4676 13198
rect 4620 13076 4676 13132
rect 4620 13074 4900 13076
rect 4620 13022 4622 13074
rect 4674 13022 4900 13074
rect 4620 13020 4900 13022
rect 4620 13010 4676 13020
rect 4508 12964 4564 12974
rect 3500 12404 3556 12414
rect 3500 12310 3556 12348
rect 3388 12238 3390 12290
rect 3442 12238 3444 12290
rect 3388 12226 3444 12238
rect 3724 12290 3780 12302
rect 3724 12238 3726 12290
rect 3778 12238 3780 12290
rect 3724 12180 3780 12238
rect 4508 12290 4564 12908
rect 4508 12238 4510 12290
rect 4562 12238 4564 12290
rect 4508 12226 4564 12238
rect 4844 12740 4900 13020
rect 4956 12964 5012 13804
rect 5516 13972 5572 13982
rect 5516 13858 5572 13916
rect 5964 13972 6020 14254
rect 5964 13906 6020 13916
rect 6188 13970 6244 14476
rect 6188 13918 6190 13970
rect 6242 13918 6244 13970
rect 6188 13906 6244 13918
rect 6300 14306 6356 14318
rect 6300 14254 6302 14306
rect 6354 14254 6356 14306
rect 6300 14084 6356 14254
rect 5516 13806 5518 13858
rect 5570 13806 5572 13858
rect 5516 13794 5572 13806
rect 5628 13858 5684 13870
rect 5628 13806 5630 13858
rect 5682 13806 5684 13858
rect 5628 13188 5684 13806
rect 4956 12898 5012 12908
rect 5068 13132 5684 13188
rect 5852 13746 5908 13758
rect 5852 13694 5854 13746
rect 5906 13694 5908 13746
rect 3836 12180 3892 12190
rect 3724 12178 3892 12180
rect 3724 12126 3838 12178
rect 3890 12126 3892 12178
rect 3724 12124 3892 12126
rect 3836 12114 3892 12124
rect 4284 12178 4340 12190
rect 4284 12126 4286 12178
rect 4338 12126 4340 12178
rect 1820 11394 1876 11452
rect 2492 12068 2548 12078
rect 2492 11506 2548 12012
rect 4060 12068 4116 12078
rect 4060 11974 4116 12012
rect 2492 11454 2494 11506
rect 2546 11454 2548 11506
rect 2492 11442 2548 11454
rect 1820 11342 1822 11394
rect 1874 11342 1876 11394
rect 1820 11330 1876 11342
rect 4284 10836 4340 12126
rect 4844 12178 4900 12684
rect 5068 12404 5124 13132
rect 5628 12964 5684 12974
rect 5628 12870 5684 12908
rect 5852 12962 5908 13694
rect 6076 13746 6132 13758
rect 6076 13694 6078 13746
rect 6130 13694 6132 13746
rect 5852 12910 5854 12962
rect 5906 12910 5908 12962
rect 5852 12898 5908 12910
rect 5964 13076 6020 13086
rect 5180 12738 5236 12750
rect 5180 12686 5182 12738
rect 5234 12686 5236 12738
rect 5180 12628 5236 12686
rect 5964 12738 6020 13020
rect 5964 12686 5966 12738
rect 6018 12686 6020 12738
rect 5964 12674 6020 12686
rect 5180 12562 5236 12572
rect 5068 12180 5124 12348
rect 5628 12292 5684 12302
rect 6076 12292 6132 13694
rect 6300 13188 6356 14028
rect 6412 13970 6468 16044
rect 6524 15314 6580 16828
rect 6748 15540 6804 17390
rect 6748 15474 6804 15484
rect 6524 15262 6526 15314
rect 6578 15262 6580 15314
rect 6524 15204 6580 15262
rect 6748 15316 6804 15326
rect 6748 15222 6804 15260
rect 6524 15138 6580 15148
rect 6860 15092 6916 17502
rect 7196 17554 7252 17566
rect 7196 17502 7198 17554
rect 7250 17502 7252 17554
rect 7196 16884 7252 17502
rect 7196 16818 7252 16828
rect 7084 16772 7140 16782
rect 6972 15428 7028 15438
rect 6972 15334 7028 15372
rect 7084 15426 7140 16716
rect 7420 15652 7476 18398
rect 7756 18452 7812 18510
rect 7756 18386 7812 18396
rect 8316 18562 8372 19182
rect 8540 19234 8596 21534
rect 8876 21586 8932 21598
rect 8876 21534 8878 21586
rect 8930 21534 8932 21586
rect 8876 20356 8932 21534
rect 9772 21586 9828 21598
rect 9772 21534 9774 21586
rect 9826 21534 9828 21586
rect 9660 21364 9716 21374
rect 9660 21270 9716 21308
rect 8764 20300 8932 20356
rect 9660 20914 9716 20926
rect 9660 20862 9662 20914
rect 9714 20862 9716 20914
rect 8540 19182 8542 19234
rect 8594 19182 8596 19234
rect 8540 19170 8596 19182
rect 8652 19796 8708 19806
rect 8652 19010 8708 19740
rect 8764 19236 8820 20300
rect 9660 20242 9716 20862
rect 9660 20190 9662 20242
rect 9714 20190 9716 20242
rect 9660 20188 9716 20190
rect 8876 20132 9716 20188
rect 8876 20130 8932 20132
rect 8876 20078 8878 20130
rect 8930 20078 8932 20130
rect 8876 20066 8932 20078
rect 9436 20020 9492 20030
rect 8988 20018 9492 20020
rect 8988 19966 9438 20018
rect 9490 19966 9492 20018
rect 8988 19964 9492 19966
rect 8876 19236 8932 19246
rect 8764 19180 8876 19236
rect 8876 19170 8932 19180
rect 8988 19234 9044 19964
rect 9436 19954 9492 19964
rect 9548 19796 9604 20132
rect 8988 19182 8990 19234
rect 9042 19182 9044 19234
rect 8988 19170 9044 19182
rect 9324 19740 9604 19796
rect 9772 20018 9828 21534
rect 10108 20804 10164 20814
rect 10108 20710 10164 20748
rect 10332 20188 10388 22316
rect 10556 21700 10612 21710
rect 10892 21700 10948 21710
rect 10556 21698 10836 21700
rect 10556 21646 10558 21698
rect 10610 21646 10836 21698
rect 10556 21644 10836 21646
rect 10556 21634 10612 21644
rect 10780 20914 10836 21644
rect 10892 21606 10948 21644
rect 10780 20862 10782 20914
rect 10834 20862 10836 20914
rect 10780 20850 10836 20862
rect 9772 19966 9774 20018
rect 9826 19966 9828 20018
rect 9324 19122 9380 19740
rect 9324 19070 9326 19122
rect 9378 19070 9380 19122
rect 9324 19058 9380 19070
rect 9436 19236 9492 19246
rect 9436 19124 9492 19180
rect 9772 19124 9828 19966
rect 9436 19122 9604 19124
rect 9436 19070 9438 19122
rect 9490 19070 9604 19122
rect 9436 19068 9604 19070
rect 9436 19058 9492 19068
rect 9100 19012 9156 19022
rect 8652 18958 8654 19010
rect 8706 18958 8708 19010
rect 8652 18946 8708 18958
rect 8988 19010 9156 19012
rect 8988 18958 9102 19010
rect 9154 18958 9156 19010
rect 8988 18956 9156 18958
rect 8988 18676 9044 18956
rect 9100 18946 9156 18956
rect 8316 18510 8318 18562
rect 8370 18510 8372 18562
rect 7868 18340 7924 18350
rect 7532 18228 7588 18238
rect 7532 17554 7588 18172
rect 7532 17502 7534 17554
rect 7586 17502 7588 17554
rect 7532 17490 7588 17502
rect 7756 17668 7812 17678
rect 7084 15374 7086 15426
rect 7138 15374 7140 15426
rect 7084 15362 7140 15374
rect 7196 15596 7476 15652
rect 7756 15652 7812 17612
rect 7868 16882 7924 18284
rect 8316 18228 8372 18510
rect 8540 18620 9044 18676
rect 8540 18562 8596 18620
rect 8540 18510 8542 18562
rect 8594 18510 8596 18562
rect 8540 18498 8596 18510
rect 8988 18452 9044 18462
rect 9436 18452 9492 18462
rect 8988 18450 9492 18452
rect 8988 18398 8990 18450
rect 9042 18398 9438 18450
rect 9490 18398 9492 18450
rect 8988 18396 9492 18398
rect 8988 18386 9044 18396
rect 9436 18386 9492 18396
rect 9548 18452 9604 19068
rect 8764 18340 8820 18350
rect 8652 18338 8820 18340
rect 8652 18286 8766 18338
rect 8818 18286 8820 18338
rect 8652 18284 8820 18286
rect 8372 18172 8596 18228
rect 8316 18134 8372 18172
rect 7868 16830 7870 16882
rect 7922 16830 7924 16882
rect 7868 16818 7924 16830
rect 7980 17666 8036 17678
rect 7980 17614 7982 17666
rect 8034 17614 8036 17666
rect 7980 16212 8036 17614
rect 8092 17444 8148 17454
rect 8092 16882 8148 17388
rect 8540 17108 8596 18172
rect 8652 17778 8708 18284
rect 8764 18274 8820 18284
rect 8652 17726 8654 17778
rect 8706 17726 8708 17778
rect 8652 17714 8708 17726
rect 9436 17444 9492 17454
rect 8540 17052 8708 17108
rect 8092 16830 8094 16882
rect 8146 16830 8148 16882
rect 8092 16818 8148 16830
rect 8540 16884 8596 16894
rect 8540 16790 8596 16828
rect 8652 16882 8708 17052
rect 8652 16830 8654 16882
rect 8706 16830 8708 16882
rect 8652 16818 8708 16830
rect 8316 16770 8372 16782
rect 8316 16718 8318 16770
rect 8370 16718 8372 16770
rect 8316 16324 8372 16718
rect 7980 16146 8036 16156
rect 8092 16268 8372 16324
rect 8092 16210 8148 16268
rect 8092 16158 8094 16210
rect 8146 16158 8148 16210
rect 8092 16146 8148 16158
rect 8876 16100 8932 16110
rect 7756 15596 8372 15652
rect 7196 15148 7252 15596
rect 7756 15540 7812 15596
rect 6860 15026 6916 15036
rect 6972 15092 7252 15148
rect 7308 15538 7812 15540
rect 7308 15486 7758 15538
rect 7810 15486 7812 15538
rect 7308 15484 7812 15486
rect 6860 14756 6916 14766
rect 6860 14530 6916 14700
rect 6860 14478 6862 14530
rect 6914 14478 6916 14530
rect 6860 14466 6916 14478
rect 6636 14308 6692 14318
rect 6972 14308 7028 15092
rect 7084 14868 7140 14878
rect 7084 14418 7140 14812
rect 7084 14366 7086 14418
rect 7138 14366 7140 14418
rect 7084 14354 7140 14366
rect 7196 14418 7252 14430
rect 7196 14366 7198 14418
rect 7250 14366 7252 14418
rect 6636 14306 7028 14308
rect 6636 14254 6638 14306
rect 6690 14254 7028 14306
rect 6636 14252 7028 14254
rect 6636 14242 6692 14252
rect 6412 13918 6414 13970
rect 6466 13918 6468 13970
rect 6412 13906 6468 13918
rect 6748 13972 6804 14252
rect 6972 14084 7028 14252
rect 7196 14084 7252 14366
rect 6972 14028 7140 14084
rect 6748 13906 6804 13916
rect 6636 13858 6692 13870
rect 6636 13806 6638 13858
rect 6690 13806 6692 13858
rect 6636 13636 6692 13806
rect 6300 13132 6580 13188
rect 6188 13020 6468 13076
rect 6188 12962 6244 13020
rect 6188 12910 6190 12962
rect 6242 12910 6244 12962
rect 6188 12898 6244 12910
rect 6412 12962 6468 13020
rect 6412 12910 6414 12962
rect 6466 12910 6468 12962
rect 6412 12898 6468 12910
rect 5628 12290 6132 12292
rect 5628 12238 5630 12290
rect 5682 12238 6132 12290
rect 5628 12236 6132 12238
rect 5628 12226 5684 12236
rect 4844 12126 4846 12178
rect 4898 12126 4900 12178
rect 4844 12114 4900 12126
rect 4956 12178 5124 12180
rect 4956 12126 5070 12178
rect 5122 12126 5124 12178
rect 4956 12124 5124 12126
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4956 11620 5012 12124
rect 5068 12114 5124 12124
rect 5964 12066 6020 12078
rect 5964 12014 5966 12066
rect 6018 12014 6020 12066
rect 5292 11956 5348 11966
rect 5516 11956 5572 11966
rect 5292 11954 5460 11956
rect 5292 11902 5294 11954
rect 5346 11902 5460 11954
rect 5292 11900 5460 11902
rect 5292 11890 5348 11900
rect 5404 11732 5460 11900
rect 5516 11862 5572 11900
rect 5964 11732 6020 12014
rect 5404 11676 6020 11732
rect 4620 11564 5012 11620
rect 4620 11506 4676 11564
rect 4620 11454 4622 11506
rect 4674 11454 4676 11506
rect 4620 11442 4676 11454
rect 5292 11508 5348 11518
rect 5348 11452 5460 11508
rect 5292 11442 5348 11452
rect 4284 10770 4340 10780
rect 5068 11170 5124 11182
rect 5068 11118 5070 11170
rect 5122 11118 5124 11170
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4732 9828 4788 9838
rect 4732 9734 4788 9772
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4620 8484 4676 8494
rect 4620 7474 4676 8428
rect 5068 8260 5124 11118
rect 5292 10500 5348 10510
rect 5180 10498 5348 10500
rect 5180 10446 5294 10498
rect 5346 10446 5348 10498
rect 5180 10444 5348 10446
rect 5180 9716 5236 10444
rect 5292 10434 5348 10444
rect 5180 9622 5236 9660
rect 5292 9044 5348 9054
rect 5404 9044 5460 11452
rect 5516 10836 5572 10846
rect 5516 10742 5572 10780
rect 5740 10836 5796 11676
rect 6524 11620 6580 13132
rect 6636 12964 6692 13580
rect 6972 13746 7028 13758
rect 6972 13694 6974 13746
rect 7026 13694 7028 13746
rect 6972 13412 7028 13694
rect 6972 13346 7028 13356
rect 6636 12908 6804 12964
rect 6748 12850 6804 12908
rect 7084 12962 7140 14028
rect 7196 14018 7252 14028
rect 7308 13970 7364 15484
rect 7756 15474 7812 15484
rect 8092 15426 8148 15438
rect 8092 15374 8094 15426
rect 8146 15374 8148 15426
rect 8092 15092 8148 15374
rect 8092 14532 8148 15036
rect 8092 14466 8148 14476
rect 8204 15428 8260 15438
rect 8092 14306 8148 14318
rect 8092 14254 8094 14306
rect 8146 14254 8148 14306
rect 8092 14196 8148 14254
rect 8092 14130 8148 14140
rect 7308 13918 7310 13970
rect 7362 13918 7364 13970
rect 7308 13906 7364 13918
rect 8204 13970 8260 15372
rect 8316 14530 8372 15596
rect 8428 15540 8484 15550
rect 8428 15426 8484 15484
rect 8428 15374 8430 15426
rect 8482 15374 8484 15426
rect 8428 15362 8484 15374
rect 8652 15538 8708 15550
rect 8652 15486 8654 15538
rect 8706 15486 8708 15538
rect 8652 14754 8708 15486
rect 8764 15428 8820 15438
rect 8764 15334 8820 15372
rect 8876 15204 8932 16044
rect 9324 16100 9380 16110
rect 9436 16100 9492 17388
rect 9548 16994 9604 18396
rect 9660 18562 9716 18574
rect 9660 18510 9662 18562
rect 9714 18510 9716 18562
rect 9660 17780 9716 18510
rect 9772 18562 9828 19068
rect 10220 20132 10388 20188
rect 10556 20244 10612 20254
rect 9772 18510 9774 18562
rect 9826 18510 9828 18562
rect 9772 18498 9828 18510
rect 9996 19010 10052 19022
rect 9996 18958 9998 19010
rect 10050 18958 10052 19010
rect 9996 18226 10052 18958
rect 10220 18340 10276 20132
rect 10220 18246 10276 18284
rect 9996 18174 9998 18226
rect 10050 18174 10052 18226
rect 9996 18162 10052 18174
rect 9660 17108 9716 17724
rect 9660 17106 10052 17108
rect 9660 17054 9662 17106
rect 9714 17054 10052 17106
rect 9660 17052 10052 17054
rect 9660 17042 9716 17052
rect 9548 16942 9550 16994
rect 9602 16942 9604 16994
rect 9548 16930 9604 16942
rect 9884 16884 9940 16894
rect 9884 16790 9940 16828
rect 9548 16548 9604 16558
rect 9548 16322 9604 16492
rect 9548 16270 9550 16322
rect 9602 16270 9604 16322
rect 9548 16258 9604 16270
rect 9884 16324 9940 16334
rect 9772 16100 9828 16110
rect 9436 16098 9828 16100
rect 9436 16046 9774 16098
rect 9826 16046 9828 16098
rect 9436 16044 9828 16046
rect 9324 16006 9380 16044
rect 8988 15876 9044 15886
rect 8988 15426 9044 15820
rect 8988 15374 8990 15426
rect 9042 15374 9044 15426
rect 8988 15362 9044 15374
rect 9772 15148 9828 16044
rect 8876 15138 8932 15148
rect 9548 15092 9828 15148
rect 9884 15540 9940 16268
rect 9996 16322 10052 17052
rect 10108 16770 10164 16782
rect 10108 16718 10110 16770
rect 10162 16718 10164 16770
rect 10108 16548 10164 16718
rect 10108 16482 10164 16492
rect 9996 16270 9998 16322
rect 10050 16270 10052 16322
rect 9996 16258 10052 16270
rect 10556 16100 10612 20188
rect 10668 18338 10724 18350
rect 10668 18286 10670 18338
rect 10722 18286 10724 18338
rect 10668 18226 10724 18286
rect 10668 18174 10670 18226
rect 10722 18174 10724 18226
rect 10668 16324 10724 18174
rect 10780 17780 10836 17790
rect 10780 17686 10836 17724
rect 10668 16258 10724 16268
rect 10668 16100 10724 16110
rect 10556 16098 10724 16100
rect 10556 16046 10670 16098
rect 10722 16046 10724 16098
rect 10556 16044 10724 16046
rect 10668 16034 10724 16044
rect 10892 16098 10948 16110
rect 10892 16046 10894 16098
rect 10946 16046 10948 16098
rect 10108 15988 10164 15998
rect 10444 15988 10500 15998
rect 10108 15986 10500 15988
rect 10108 15934 10110 15986
rect 10162 15934 10446 15986
rect 10498 15934 10500 15986
rect 10108 15932 10500 15934
rect 10108 15922 10164 15932
rect 10444 15922 10500 15932
rect 10556 15876 10612 15886
rect 10556 15782 10612 15820
rect 8652 14702 8654 14754
rect 8706 14702 8708 14754
rect 8652 14690 8708 14702
rect 9212 14980 9268 14990
rect 9212 14642 9268 14924
rect 9212 14590 9214 14642
rect 9266 14590 9268 14642
rect 9212 14578 9268 14590
rect 9548 14644 9604 15092
rect 8316 14478 8318 14530
rect 8370 14478 8372 14530
rect 8316 14466 8372 14478
rect 9436 14532 9492 14542
rect 9436 14438 9492 14476
rect 9548 14418 9604 14588
rect 9548 14366 9550 14418
rect 9602 14366 9604 14418
rect 9548 14354 9604 14366
rect 8540 14306 8596 14318
rect 8540 14254 8542 14306
rect 8594 14254 8596 14306
rect 8204 13918 8206 13970
rect 8258 13918 8260 13970
rect 8204 13906 8260 13918
rect 8316 14084 8372 14094
rect 8316 13858 8372 14028
rect 8316 13806 8318 13858
rect 8370 13806 8372 13858
rect 8316 13794 8372 13806
rect 7644 13746 7700 13758
rect 7644 13694 7646 13746
rect 7698 13694 7700 13746
rect 7644 13412 7700 13694
rect 7980 13748 8036 13758
rect 8540 13748 8596 14254
rect 9772 14308 9828 14318
rect 9772 14214 9828 14252
rect 8876 14084 8932 14094
rect 8764 14028 8876 14084
rect 8652 13748 8708 13758
rect 8540 13746 8708 13748
rect 8540 13694 8654 13746
rect 8706 13694 8708 13746
rect 8540 13692 8708 13694
rect 7980 13654 8036 13692
rect 8652 13682 8708 13692
rect 7644 13346 7700 13356
rect 7644 13074 7700 13086
rect 7644 13022 7646 13074
rect 7698 13022 7700 13074
rect 7644 12964 7700 13022
rect 8764 13076 8820 14028
rect 8876 14018 8932 14028
rect 9772 13972 9828 13982
rect 9884 13972 9940 15484
rect 10892 15428 10948 16046
rect 10892 15362 10948 15372
rect 10108 15204 10164 15214
rect 10108 14530 10164 15148
rect 10108 14478 10110 14530
rect 10162 14478 10164 14530
rect 9772 13970 9940 13972
rect 9772 13918 9774 13970
rect 9826 13918 9940 13970
rect 9772 13916 9940 13918
rect 9996 13972 10052 13982
rect 9772 13906 9828 13916
rect 9996 13878 10052 13916
rect 8876 13634 8932 13646
rect 8876 13582 8878 13634
rect 8930 13582 8932 13634
rect 8876 13188 8932 13582
rect 8988 13524 9044 13534
rect 8988 13522 9716 13524
rect 8988 13470 8990 13522
rect 9042 13470 9716 13522
rect 8988 13468 9716 13470
rect 8988 13458 9044 13468
rect 9660 13300 9716 13468
rect 9660 13244 9940 13300
rect 8876 13132 9828 13188
rect 8764 13020 9604 13076
rect 7084 12910 7086 12962
rect 7138 12910 7140 12962
rect 7084 12898 7140 12910
rect 7196 12908 7700 12964
rect 6748 12798 6750 12850
rect 6802 12798 6804 12850
rect 6636 12740 6692 12750
rect 6636 12646 6692 12684
rect 5740 10742 5796 10780
rect 5852 11564 6580 11620
rect 5852 10722 5908 11564
rect 6412 10836 6468 10846
rect 6636 10836 6692 10846
rect 6468 10834 6692 10836
rect 6468 10782 6638 10834
rect 6690 10782 6692 10834
rect 6468 10780 6692 10782
rect 6412 10770 6468 10780
rect 6636 10770 6692 10780
rect 5852 10670 5854 10722
rect 5906 10670 5908 10722
rect 5852 10658 5908 10670
rect 6524 10612 6580 10622
rect 6748 10612 6804 12798
rect 7196 12850 7252 12908
rect 7196 12798 7198 12850
rect 7250 12798 7252 12850
rect 7196 11956 7252 12798
rect 7196 11890 7252 11900
rect 7420 12738 7476 12750
rect 7420 12686 7422 12738
rect 7474 12686 7476 12738
rect 6524 10610 6804 10612
rect 6524 10558 6526 10610
rect 6578 10558 6804 10610
rect 6524 10556 6804 10558
rect 6860 10722 6916 10734
rect 6860 10670 6862 10722
rect 6914 10670 6916 10722
rect 6860 10612 6916 10670
rect 7420 10722 7476 12686
rect 7644 12404 7700 12908
rect 7644 12338 7700 12348
rect 9548 12402 9604 13020
rect 9772 13074 9828 13132
rect 9772 13022 9774 13074
rect 9826 13022 9828 13074
rect 9772 13010 9828 13022
rect 9884 12740 9940 13244
rect 10108 12964 10164 14478
rect 10780 14418 10836 14430
rect 10780 14366 10782 14418
rect 10834 14366 10836 14418
rect 10556 14308 10612 14318
rect 10332 13860 10388 13870
rect 10332 13766 10388 13804
rect 10556 13746 10612 14252
rect 10780 13970 10836 14366
rect 10780 13918 10782 13970
rect 10834 13918 10836 13970
rect 10780 13906 10836 13918
rect 10556 13694 10558 13746
rect 10610 13694 10612 13746
rect 10556 13682 10612 13694
rect 10892 13748 10948 13758
rect 10892 13654 10948 13692
rect 10556 12964 10612 12974
rect 10108 12962 10612 12964
rect 10108 12910 10558 12962
rect 10610 12910 10612 12962
rect 10108 12908 10612 12910
rect 9548 12350 9550 12402
rect 9602 12350 9604 12402
rect 9548 12338 9604 12350
rect 9660 12684 9940 12740
rect 9660 12402 9716 12684
rect 9660 12350 9662 12402
rect 9714 12350 9716 12402
rect 9660 12338 9716 12350
rect 9772 12404 9828 12414
rect 9772 12310 9828 12348
rect 8764 12178 8820 12190
rect 8764 12126 8766 12178
rect 8818 12126 8820 12178
rect 8092 12068 8148 12078
rect 7420 10670 7422 10722
rect 7474 10670 7476 10722
rect 7420 10658 7476 10670
rect 7532 12066 8148 12068
rect 7532 12014 8094 12066
rect 8146 12014 8148 12066
rect 7532 12012 8148 12014
rect 6972 10612 7028 10622
rect 6860 10610 7028 10612
rect 6860 10558 6974 10610
rect 7026 10558 7028 10610
rect 6860 10556 7028 10558
rect 6524 10546 6580 10556
rect 6972 10546 7028 10556
rect 7196 10500 7252 10510
rect 7532 10500 7588 12012
rect 8092 12002 8148 12012
rect 8764 11508 8820 12126
rect 10220 12178 10276 12190
rect 10220 12126 10222 12178
rect 10274 12126 10276 12178
rect 8764 11414 8820 11452
rect 9100 11732 9156 11742
rect 9100 10834 9156 11676
rect 9100 10782 9102 10834
rect 9154 10782 9156 10834
rect 9100 10770 9156 10782
rect 9996 11732 10052 11742
rect 7196 10498 7588 10500
rect 7196 10446 7198 10498
rect 7250 10446 7588 10498
rect 7196 10444 7588 10446
rect 7644 10610 7700 10622
rect 7644 10558 7646 10610
rect 7698 10558 7700 10610
rect 7196 10434 7252 10444
rect 5852 10052 5908 10062
rect 5852 9938 5908 9996
rect 7644 10052 7700 10558
rect 7644 9986 7700 9996
rect 7980 10498 8036 10510
rect 7980 10446 7982 10498
rect 8034 10446 8036 10498
rect 5852 9886 5854 9938
rect 5906 9886 5908 9938
rect 5852 9874 5908 9886
rect 7308 9828 7364 9838
rect 7756 9828 7812 9838
rect 7308 9826 7812 9828
rect 7308 9774 7310 9826
rect 7362 9774 7758 9826
rect 7810 9774 7812 9826
rect 7308 9772 7812 9774
rect 7308 9762 7364 9772
rect 7756 9762 7812 9772
rect 7868 9828 7924 9838
rect 7980 9828 8036 10446
rect 9772 10500 9828 10510
rect 8204 10386 8260 10398
rect 8204 10334 8206 10386
rect 8258 10334 8260 10386
rect 8204 10164 8260 10334
rect 8540 10388 8596 10398
rect 9436 10388 9492 10398
rect 8540 10386 8708 10388
rect 8540 10334 8542 10386
rect 8594 10334 8708 10386
rect 8540 10332 8708 10334
rect 8540 10322 8596 10332
rect 7868 9826 8036 9828
rect 7868 9774 7870 9826
rect 7922 9774 8036 9826
rect 7868 9772 8036 9774
rect 7868 9762 7924 9772
rect 5964 9604 6020 9614
rect 5964 9154 6020 9548
rect 6300 9604 6356 9614
rect 6300 9602 6580 9604
rect 6300 9550 6302 9602
rect 6354 9550 6580 9602
rect 6300 9548 6580 9550
rect 6300 9538 6356 9548
rect 5964 9102 5966 9154
rect 6018 9102 6020 9154
rect 5964 9090 6020 9102
rect 5292 9042 5460 9044
rect 5292 8990 5294 9042
rect 5346 8990 5460 9042
rect 5292 8988 5460 8990
rect 4620 7422 4622 7474
rect 4674 7422 4676 7474
rect 4620 7410 4676 7422
rect 4956 8204 5124 8260
rect 5180 8596 5236 8606
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4732 6468 4788 6478
rect 4956 6468 5012 8204
rect 4620 6466 5012 6468
rect 4620 6414 4734 6466
rect 4786 6414 5012 6466
rect 4620 6412 5012 6414
rect 5068 8034 5124 8046
rect 5068 7982 5070 8034
rect 5122 7982 5124 8034
rect 5068 6804 5124 7982
rect 4620 5908 4676 6412
rect 4732 6402 4788 6412
rect 5068 6244 5124 6748
rect 5180 6690 5236 8540
rect 5292 8484 5348 8988
rect 6524 8484 6580 9548
rect 6636 9602 6692 9614
rect 6636 9550 6638 9602
rect 6690 9550 6692 9602
rect 6636 8708 6692 9550
rect 6636 8642 6692 8652
rect 7084 9602 7140 9614
rect 7084 9550 7086 9602
rect 7138 9550 7140 9602
rect 6524 8428 6916 8484
rect 5292 8418 5348 8428
rect 5292 8036 5348 8046
rect 5292 7586 5348 7980
rect 6076 8034 6132 8046
rect 6076 7982 6078 8034
rect 6130 7982 6132 8034
rect 6076 7588 6132 7982
rect 5292 7534 5294 7586
rect 5346 7534 5348 7586
rect 5292 7522 5348 7534
rect 5964 7532 6076 7588
rect 5964 6802 6020 7532
rect 6076 7522 6132 7532
rect 6636 8034 6692 8046
rect 6636 7982 6638 8034
rect 6690 7982 6692 8034
rect 6524 7476 6580 7486
rect 6412 7420 6524 7476
rect 5964 6750 5966 6802
rect 6018 6750 6020 6802
rect 5964 6738 6020 6750
rect 6188 6916 6244 6926
rect 5180 6638 5182 6690
rect 5234 6638 5236 6690
rect 5180 6626 5236 6638
rect 4732 6188 5124 6244
rect 4732 6130 4788 6188
rect 4732 6078 4734 6130
rect 4786 6078 4788 6130
rect 4732 6066 4788 6078
rect 6188 6018 6244 6860
rect 6300 6692 6356 6702
rect 6300 6598 6356 6636
rect 6188 5966 6190 6018
rect 6242 5966 6244 6018
rect 6188 5954 6244 5966
rect 4620 5852 4900 5908
rect 4284 5794 4340 5806
rect 4284 5742 4286 5794
rect 4338 5742 4340 5794
rect 4284 5682 4340 5742
rect 4284 5630 4286 5682
rect 4338 5630 4340 5682
rect 4284 5618 4340 5630
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4844 5348 4900 5852
rect 5516 5906 5572 5918
rect 5516 5854 5518 5906
rect 5570 5854 5572 5906
rect 5180 5796 5236 5806
rect 5180 5702 5236 5740
rect 5068 5682 5124 5694
rect 5068 5630 5070 5682
rect 5122 5630 5124 5682
rect 5068 5460 5124 5630
rect 5180 5460 5236 5470
rect 5068 5404 5180 5460
rect 4844 4562 4900 5292
rect 5180 5234 5236 5404
rect 5180 5182 5182 5234
rect 5234 5182 5236 5234
rect 5180 5170 5236 5182
rect 4844 4510 4846 4562
rect 4898 4510 4900 4562
rect 4844 4498 4900 4510
rect 5068 5012 5124 5022
rect 5068 4338 5124 4956
rect 5516 5012 5572 5854
rect 6076 5796 6132 5806
rect 6076 5234 6132 5740
rect 6076 5182 6078 5234
rect 6130 5182 6132 5234
rect 6076 5170 6132 5182
rect 5516 4946 5572 4956
rect 5068 4286 5070 4338
rect 5122 4286 5124 4338
rect 5068 4274 5124 4286
rect 5852 4228 5908 4238
rect 5852 4134 5908 4172
rect 5068 4116 5124 4126
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 5068 3666 5124 4060
rect 5068 3614 5070 3666
rect 5122 3614 5124 3666
rect 5068 3602 5124 3614
rect 6412 3668 6468 7420
rect 6524 7410 6580 7420
rect 6636 7028 6692 7982
rect 6636 6962 6692 6972
rect 6636 6804 6692 6814
rect 6636 6692 6692 6748
rect 6748 6692 6804 6702
rect 6636 6690 6804 6692
rect 6636 6638 6750 6690
rect 6802 6638 6804 6690
rect 6636 6636 6804 6638
rect 6748 6626 6804 6636
rect 6860 6468 6916 8428
rect 7084 8372 7140 9550
rect 7196 9604 7252 9614
rect 7196 9510 7252 9548
rect 7644 9604 7700 9614
rect 7644 9510 7700 9548
rect 7980 8932 8036 9772
rect 8092 10108 8204 10164
rect 8092 9604 8148 10108
rect 8204 10098 8260 10108
rect 8092 9538 8148 9548
rect 8204 9940 8260 9950
rect 8092 8932 8148 8942
rect 7980 8930 8148 8932
rect 7980 8878 8094 8930
rect 8146 8878 8148 8930
rect 7980 8876 8148 8878
rect 8092 8866 8148 8876
rect 8204 8708 8260 9884
rect 7084 8306 7140 8316
rect 8092 8652 8260 8708
rect 8316 9826 8372 9838
rect 8316 9774 8318 9826
rect 8370 9774 8372 9826
rect 8316 9604 8372 9774
rect 7196 8260 7252 8270
rect 7644 8260 7700 8270
rect 7196 8258 7700 8260
rect 7196 8206 7198 8258
rect 7250 8206 7646 8258
rect 7698 8206 7700 8258
rect 7196 8204 7700 8206
rect 7196 8194 7252 8204
rect 7644 8194 7700 8204
rect 7756 8260 7812 8270
rect 6972 8148 7028 8158
rect 6972 8054 7028 8092
rect 7084 8036 7140 8046
rect 7084 7942 7140 7980
rect 7532 8036 7588 8046
rect 7532 7942 7588 7980
rect 7756 7812 7812 8204
rect 7420 7756 7812 7812
rect 7868 8036 7924 8046
rect 8092 8036 8148 8652
rect 8204 8260 8260 8270
rect 8316 8260 8372 9548
rect 8540 9380 8596 9390
rect 8540 9266 8596 9324
rect 8540 9214 8542 9266
rect 8594 9214 8596 9266
rect 8204 8258 8372 8260
rect 8204 8206 8206 8258
rect 8258 8206 8372 8258
rect 8204 8204 8372 8206
rect 8428 8260 8484 8270
rect 8204 8194 8260 8204
rect 8428 8166 8484 8204
rect 8092 7980 8484 8036
rect 7420 7362 7476 7756
rect 7420 7310 7422 7362
rect 7474 7310 7476 7362
rect 7420 7298 7476 7310
rect 7756 7588 7812 7598
rect 7868 7588 7924 7980
rect 7756 7586 7924 7588
rect 7756 7534 7758 7586
rect 7810 7534 7924 7586
rect 7756 7532 7924 7534
rect 7756 7252 7812 7532
rect 7980 7476 8036 7486
rect 7980 7474 8260 7476
rect 7980 7422 7982 7474
rect 8034 7422 8260 7474
rect 7980 7420 8260 7422
rect 7980 7410 8036 7420
rect 7756 7186 7812 7196
rect 7868 7362 7924 7374
rect 7868 7310 7870 7362
rect 7922 7310 7924 7362
rect 7868 7028 7924 7310
rect 7420 6972 7924 7028
rect 8092 7252 8148 7262
rect 7084 6916 7140 6926
rect 7084 6822 7140 6860
rect 7420 6914 7476 6972
rect 7420 6862 7422 6914
rect 7474 6862 7476 6914
rect 7420 6850 7476 6862
rect 8092 6914 8148 7196
rect 8092 6862 8094 6914
rect 8146 6862 8148 6914
rect 8092 6850 8148 6862
rect 8204 6804 8260 7420
rect 8316 7474 8372 7486
rect 8316 7422 8318 7474
rect 8370 7422 8372 7474
rect 8316 7028 8372 7422
rect 8428 7476 8484 7980
rect 8428 7410 8484 7420
rect 8316 6972 8484 7028
rect 8316 6804 8372 6814
rect 8204 6802 8372 6804
rect 8204 6750 8318 6802
rect 8370 6750 8372 6802
rect 8204 6748 8372 6750
rect 7196 6468 7252 6478
rect 7756 6468 7812 6478
rect 6860 6412 7028 6468
rect 6524 5348 6580 5358
rect 6524 5234 6580 5292
rect 6524 5182 6526 5234
rect 6578 5182 6580 5234
rect 6524 5170 6580 5182
rect 6860 4900 6916 4910
rect 6860 4806 6916 4844
rect 6524 3668 6580 3678
rect 6412 3666 6580 3668
rect 6412 3614 6526 3666
rect 6578 3614 6580 3666
rect 6412 3612 6580 3614
rect 6524 3602 6580 3612
rect 1708 3332 1764 3342
rect 3164 3332 3220 3342
rect 1148 3330 1764 3332
rect 1148 3278 1710 3330
rect 1762 3278 1764 3330
rect 1148 3276 1764 3278
rect 1148 800 1204 3276
rect 1708 3266 1764 3276
rect 2940 3330 3220 3332
rect 2940 3278 3166 3330
rect 3218 3278 3220 3330
rect 2940 3276 3220 3278
rect 2940 800 2996 3276
rect 3164 3266 3220 3276
rect 4732 3332 4788 3342
rect 4732 800 4788 3276
rect 5516 3332 5572 3342
rect 6748 3332 6804 3342
rect 5516 3238 5572 3276
rect 6636 3330 6804 3332
rect 6636 3278 6750 3330
rect 6802 3278 6804 3330
rect 6636 3276 6804 3278
rect 6636 1652 6692 3276
rect 6748 3266 6804 3276
rect 6972 2772 7028 6412
rect 7196 6466 7812 6468
rect 7196 6414 7198 6466
rect 7250 6414 7758 6466
rect 7810 6414 7812 6466
rect 7196 6412 7812 6414
rect 7196 5348 7252 6412
rect 7756 6402 7812 6412
rect 8316 5794 8372 6748
rect 8316 5742 8318 5794
rect 8370 5742 8372 5794
rect 8316 5730 8372 5742
rect 8428 6580 8484 6972
rect 8540 6804 8596 9214
rect 8652 8372 8708 10332
rect 9436 9938 9492 10332
rect 9436 9886 9438 9938
rect 9490 9886 9492 9938
rect 9436 9874 9492 9886
rect 8764 9826 8820 9838
rect 8764 9774 8766 9826
rect 8818 9774 8820 9826
rect 8764 9716 8820 9774
rect 9772 9716 9828 10444
rect 8764 9660 9828 9716
rect 8988 9268 9044 9278
rect 8652 7924 8708 8316
rect 8652 7858 8708 7868
rect 8764 9212 8988 9268
rect 8540 6738 8596 6748
rect 8764 6692 8820 9212
rect 8988 9174 9044 9212
rect 9548 8370 9604 8382
rect 9548 8318 9550 8370
rect 9602 8318 9604 8370
rect 8988 8036 9044 8046
rect 8988 7942 9044 7980
rect 8988 7476 9044 7486
rect 8988 7382 9044 7420
rect 9548 6802 9604 8318
rect 9660 8034 9716 8046
rect 9660 7982 9662 8034
rect 9714 7982 9716 8034
rect 9660 7700 9716 7982
rect 9660 7634 9716 7644
rect 9772 7474 9828 9660
rect 9884 10498 9940 10510
rect 9884 10446 9886 10498
rect 9938 10446 9940 10498
rect 9884 8820 9940 10446
rect 9996 9266 10052 11676
rect 10220 10836 10276 12126
rect 10556 12180 10612 12908
rect 10780 12180 10836 12190
rect 10556 12178 10836 12180
rect 10556 12126 10782 12178
rect 10834 12126 10836 12178
rect 10556 12124 10836 12126
rect 10780 12114 10836 12124
rect 9996 9214 9998 9266
rect 10050 9214 10052 9266
rect 9996 9202 10052 9214
rect 10108 10834 10276 10836
rect 10108 10782 10222 10834
rect 10274 10782 10276 10834
rect 10108 10780 10276 10782
rect 9884 8754 9940 8764
rect 9884 8148 9940 8158
rect 9884 8054 9940 8092
rect 9772 7422 9774 7474
rect 9826 7422 9828 7474
rect 9772 7410 9828 7422
rect 9548 6750 9550 6802
rect 9602 6750 9604 6802
rect 9548 6738 9604 6750
rect 8764 6626 8820 6636
rect 8876 6690 8932 6702
rect 8876 6638 8878 6690
rect 8930 6638 8932 6690
rect 7196 5346 7364 5348
rect 7196 5294 7198 5346
rect 7250 5294 7364 5346
rect 7196 5292 7364 5294
rect 7196 5282 7252 5292
rect 7308 4900 7364 5292
rect 7420 5124 7476 5134
rect 7980 5124 8036 5134
rect 7420 5122 8036 5124
rect 7420 5070 7422 5122
rect 7474 5070 7982 5122
rect 8034 5070 8036 5122
rect 7420 5068 8036 5070
rect 7420 5058 7476 5068
rect 7756 4900 7812 4910
rect 7308 4898 7812 4900
rect 7308 4846 7758 4898
rect 7810 4846 7812 4898
rect 7308 4844 7812 4846
rect 7756 4834 7812 4844
rect 7868 4898 7924 4910
rect 7868 4846 7870 4898
rect 7922 4846 7924 4898
rect 7868 4004 7924 4846
rect 7980 4226 8036 5068
rect 8428 5124 8484 6524
rect 8428 5030 8484 5068
rect 8652 5906 8708 5918
rect 8652 5854 8654 5906
rect 8706 5854 8708 5906
rect 8540 4900 8596 4910
rect 8540 4562 8596 4844
rect 8540 4510 8542 4562
rect 8594 4510 8596 4562
rect 8540 4498 8596 4510
rect 7980 4174 7982 4226
rect 8034 4174 8036 4226
rect 7980 4162 8036 4174
rect 8428 4228 8484 4238
rect 8428 4134 8484 4172
rect 8316 4114 8372 4126
rect 8316 4062 8318 4114
rect 8370 4062 8372 4114
rect 8316 4004 8372 4062
rect 7868 3948 8372 4004
rect 8652 3780 8708 5854
rect 8876 5796 8932 6638
rect 10108 6580 10164 10780
rect 10220 10770 10276 10780
rect 10780 11394 10836 11406
rect 10780 11342 10782 11394
rect 10834 11342 10836 11394
rect 10556 10612 10612 10622
rect 10556 10518 10612 10556
rect 10780 9268 10836 11342
rect 11004 10948 11060 22652
rect 11340 22372 11396 22382
rect 11340 22278 11396 22316
rect 11452 21812 11508 23100
rect 11452 21586 11508 21756
rect 11452 21534 11454 21586
rect 11506 21534 11508 21586
rect 11452 21522 11508 21534
rect 11228 21476 11284 21486
rect 11228 21382 11284 21420
rect 11788 21476 11844 21486
rect 11788 21382 11844 21420
rect 12124 21474 12180 24220
rect 12460 24610 12516 24622
rect 12460 24558 12462 24610
rect 12514 24558 12516 24610
rect 12460 24164 12516 24558
rect 12572 24500 12628 24670
rect 13020 24724 13076 26852
rect 13132 26290 13188 27692
rect 13244 27300 13300 27310
rect 13244 26402 13300 27244
rect 13468 27186 13524 28028
rect 13804 27972 13860 27982
rect 13804 27878 13860 27916
rect 14028 27970 14084 28700
rect 14028 27918 14030 27970
rect 14082 27918 14084 27970
rect 14028 27906 14084 27918
rect 13692 27748 13748 27758
rect 14588 27748 14644 30492
rect 14700 30212 14756 30222
rect 14700 30210 14980 30212
rect 14700 30158 14702 30210
rect 14754 30158 14980 30210
rect 14700 30156 14980 30158
rect 14700 30146 14756 30156
rect 14700 29316 14756 29326
rect 14700 29222 14756 29260
rect 14924 29092 14980 30156
rect 15036 29988 15092 29998
rect 15036 29894 15092 29932
rect 15484 29316 15540 29326
rect 14924 29036 15092 29092
rect 14924 28756 14980 28766
rect 15036 28756 15092 29036
rect 15148 28756 15204 28766
rect 15036 28754 15204 28756
rect 15036 28702 15150 28754
rect 15202 28702 15204 28754
rect 15036 28700 15204 28702
rect 14700 28642 14756 28654
rect 14700 28590 14702 28642
rect 14754 28590 14756 28642
rect 14700 27972 14756 28590
rect 14700 27906 14756 27916
rect 14924 28642 14980 28700
rect 15148 28690 15204 28700
rect 14924 28590 14926 28642
rect 14978 28590 14980 28642
rect 14588 27692 14868 27748
rect 13692 27654 13748 27692
rect 14476 27634 14532 27646
rect 14476 27582 14478 27634
rect 14530 27582 14532 27634
rect 13468 27134 13470 27186
rect 13522 27134 13524 27186
rect 13468 27122 13524 27134
rect 14364 27188 14420 27198
rect 14476 27188 14532 27582
rect 14364 27186 14532 27188
rect 14364 27134 14366 27186
rect 14418 27134 14532 27186
rect 14364 27132 14532 27134
rect 14364 27122 14420 27132
rect 13916 27076 13972 27086
rect 13804 27074 13972 27076
rect 13804 27022 13918 27074
rect 13970 27022 13972 27074
rect 13804 27020 13972 27022
rect 13804 26908 13860 27020
rect 13916 27010 13972 27020
rect 13244 26350 13246 26402
rect 13298 26350 13300 26402
rect 13244 26338 13300 26350
rect 13580 26852 13860 26908
rect 13916 26852 13972 26862
rect 14476 26852 14532 27132
rect 14812 27076 14868 27692
rect 14924 27746 14980 28590
rect 15484 28530 15540 29260
rect 15484 28478 15486 28530
rect 15538 28478 15540 28530
rect 15484 28466 15540 28478
rect 15260 27972 15316 27982
rect 15036 27860 15092 27870
rect 15036 27766 15092 27804
rect 15260 27858 15316 27916
rect 15260 27806 15262 27858
rect 15314 27806 15316 27858
rect 15260 27794 15316 27806
rect 14924 27694 14926 27746
rect 14978 27694 14980 27746
rect 14924 27682 14980 27694
rect 15260 27300 15316 27310
rect 14812 27074 15204 27076
rect 14812 27022 14814 27074
rect 14866 27022 15204 27074
rect 14812 27020 15204 27022
rect 14812 27010 14868 27020
rect 13580 26404 13636 26852
rect 13580 26310 13636 26348
rect 13132 26238 13134 26290
rect 13186 26238 13188 26290
rect 13132 26226 13188 26238
rect 13692 26292 13748 26302
rect 13692 26198 13748 26236
rect 13916 24948 13972 26796
rect 14028 26796 14532 26852
rect 15036 26850 15092 26862
rect 15036 26798 15038 26850
rect 15090 26798 15092 26850
rect 14028 26402 14084 26796
rect 14924 26516 14980 26526
rect 14476 26514 14980 26516
rect 14476 26462 14926 26514
rect 14978 26462 14980 26514
rect 14476 26460 14980 26462
rect 14028 26350 14030 26402
rect 14082 26350 14084 26402
rect 14028 26338 14084 26350
rect 14140 26404 14196 26414
rect 14476 26404 14532 26460
rect 14924 26450 14980 26460
rect 14196 26348 14532 26404
rect 14140 26338 14196 26348
rect 14252 26290 14308 26348
rect 14252 26238 14254 26290
rect 14306 26238 14308 26290
rect 14252 26226 14308 26238
rect 14140 26178 14196 26190
rect 14140 26126 14142 26178
rect 14194 26126 14196 26178
rect 14140 25508 14196 26126
rect 14364 25618 14420 26348
rect 14588 26292 14644 26302
rect 14588 26198 14644 26236
rect 14476 25732 14532 25742
rect 14476 25638 14532 25676
rect 14924 25732 14980 25742
rect 15036 25732 15092 26798
rect 15148 26290 15204 27020
rect 15260 27074 15316 27244
rect 15372 27188 15428 27198
rect 15372 27186 15540 27188
rect 15372 27134 15374 27186
rect 15426 27134 15540 27186
rect 15372 27132 15540 27134
rect 15372 27122 15428 27132
rect 15260 27022 15262 27074
rect 15314 27022 15316 27074
rect 15260 27010 15316 27022
rect 15484 26964 15540 27132
rect 15484 26898 15540 26908
rect 15148 26238 15150 26290
rect 15202 26238 15204 26290
rect 15148 26226 15204 26238
rect 15372 26850 15428 26862
rect 15372 26798 15374 26850
rect 15426 26798 15428 26850
rect 14924 25730 15092 25732
rect 14924 25678 14926 25730
rect 14978 25678 15092 25730
rect 14924 25676 15092 25678
rect 15260 25956 15316 25966
rect 14924 25666 14980 25676
rect 14364 25566 14366 25618
rect 14418 25566 14420 25618
rect 14364 25554 14420 25566
rect 15260 25618 15316 25900
rect 15372 25730 15428 26798
rect 15596 25956 15652 32060
rect 16044 30996 16100 32286
rect 16044 30930 16100 30940
rect 16268 30772 16324 32508
rect 16492 32498 16548 32508
rect 16604 32564 16660 32574
rect 16716 32564 16772 33068
rect 17388 33058 17444 33068
rect 17612 33236 17668 33246
rect 17500 32674 17556 32686
rect 17500 32622 17502 32674
rect 17554 32622 17556 32674
rect 16828 32564 16884 32574
rect 16716 32562 16884 32564
rect 16716 32510 16830 32562
rect 16882 32510 16884 32562
rect 16716 32508 16884 32510
rect 16604 32470 16660 32508
rect 16828 32452 16884 32508
rect 17276 32564 17332 32574
rect 17276 32470 17332 32508
rect 16828 32386 16884 32396
rect 17276 32116 17332 32126
rect 16828 31892 16884 31902
rect 16716 31220 16772 31230
rect 16716 31108 16772 31164
rect 16828 31218 16884 31836
rect 16828 31166 16830 31218
rect 16882 31166 16884 31218
rect 16828 31154 16884 31166
rect 16380 31106 16772 31108
rect 16380 31054 16718 31106
rect 16770 31054 16772 31106
rect 16380 31052 16772 31054
rect 16380 30882 16436 31052
rect 16716 31042 16772 31052
rect 16380 30830 16382 30882
rect 16434 30830 16436 30882
rect 16380 30818 16436 30830
rect 16268 30706 16324 30716
rect 15708 29988 15764 29998
rect 15708 28642 15764 29932
rect 16828 29316 16884 29326
rect 16716 29314 16884 29316
rect 16716 29262 16830 29314
rect 16882 29262 16884 29314
rect 16716 29260 16884 29262
rect 15708 28590 15710 28642
rect 15762 28590 15764 28642
rect 15708 28578 15764 28590
rect 16268 28644 16324 28654
rect 16268 28082 16324 28588
rect 16716 28530 16772 29260
rect 16828 29250 16884 29260
rect 17052 28644 17108 28654
rect 17052 28550 17108 28588
rect 16716 28478 16718 28530
rect 16770 28478 16772 28530
rect 16604 28418 16660 28430
rect 16604 28366 16606 28418
rect 16658 28366 16660 28418
rect 16268 28030 16270 28082
rect 16322 28030 16324 28082
rect 16268 28018 16324 28030
rect 16380 28084 16436 28094
rect 16380 27990 16436 28028
rect 16604 27972 16660 28366
rect 16716 28308 16772 28478
rect 16716 28242 16772 28252
rect 17164 28418 17220 28430
rect 17164 28366 17166 28418
rect 17218 28366 17220 28418
rect 16604 27878 16660 27916
rect 15932 27860 15988 27870
rect 15820 27300 15876 27310
rect 15820 27186 15876 27244
rect 15932 27298 15988 27804
rect 15932 27246 15934 27298
rect 15986 27246 15988 27298
rect 15932 27234 15988 27246
rect 16044 27858 16100 27870
rect 16044 27806 16046 27858
rect 16098 27806 16100 27858
rect 15820 27134 15822 27186
rect 15874 27134 15876 27186
rect 15820 27122 15876 27134
rect 15708 26404 15764 26414
rect 15708 26310 15764 26348
rect 15820 26292 15876 26302
rect 15820 26198 15876 26236
rect 15372 25678 15374 25730
rect 15426 25678 15428 25730
rect 15372 25666 15428 25678
rect 15484 25900 15652 25956
rect 16044 25956 16100 27806
rect 16156 27860 16212 27870
rect 16156 27766 16212 27804
rect 16492 27860 16548 27870
rect 16380 26964 16436 27002
rect 16492 26964 16548 27804
rect 16828 27412 16884 27422
rect 16604 27076 16660 27086
rect 16604 26982 16660 27020
rect 16436 26908 16548 26964
rect 16828 26962 16884 27356
rect 17164 27186 17220 28366
rect 17164 27134 17166 27186
rect 17218 27134 17220 27186
rect 17164 27076 17220 27134
rect 17164 27010 17220 27020
rect 16828 26910 16830 26962
rect 16882 26910 16884 26962
rect 16380 26898 16436 26908
rect 16828 26898 16884 26910
rect 16716 26852 16772 26862
rect 16716 26758 16772 26796
rect 16492 26516 16548 26526
rect 16492 26422 16548 26460
rect 15260 25566 15262 25618
rect 15314 25566 15316 25618
rect 15260 25554 15316 25566
rect 14140 25442 14196 25452
rect 14812 25394 14868 25406
rect 14812 25342 14814 25394
rect 14866 25342 14868 25394
rect 14812 25284 14868 25342
rect 14812 25218 14868 25228
rect 15484 24948 15540 25900
rect 16044 25890 16100 25900
rect 16156 26290 16212 26302
rect 16156 26238 16158 26290
rect 16210 26238 16212 26290
rect 16156 25732 16212 26238
rect 16156 25666 16212 25676
rect 16380 26290 16436 26302
rect 16380 26238 16382 26290
rect 16434 26238 16436 26290
rect 16268 25508 16324 25518
rect 16156 25506 16324 25508
rect 16156 25454 16270 25506
rect 16322 25454 16324 25506
rect 16156 25452 16324 25454
rect 16044 25396 16100 25406
rect 16044 25302 16100 25340
rect 15932 25284 15988 25294
rect 13916 24892 14196 24948
rect 13804 24836 13860 24846
rect 13356 24834 13860 24836
rect 13356 24782 13806 24834
rect 13858 24782 13860 24834
rect 13356 24780 13860 24782
rect 13020 24658 13076 24668
rect 13132 24722 13188 24734
rect 13132 24670 13134 24722
rect 13186 24670 13188 24722
rect 12572 24434 12628 24444
rect 12572 24164 12628 24174
rect 12460 24162 12628 24164
rect 12460 24110 12574 24162
rect 12626 24110 12628 24162
rect 12460 24108 12628 24110
rect 12572 24098 12628 24108
rect 12908 24164 12964 24174
rect 12908 24070 12964 24108
rect 12348 24052 12404 24062
rect 12348 23958 12404 23996
rect 12236 23940 12292 23950
rect 12236 23266 12292 23884
rect 12236 23214 12238 23266
rect 12290 23214 12292 23266
rect 12236 23202 12292 23214
rect 13132 23828 13188 24670
rect 13132 23268 13188 23772
rect 13132 23202 13188 23212
rect 13356 23266 13412 24780
rect 13804 24770 13860 24780
rect 14028 24722 14084 24734
rect 14028 24670 14030 24722
rect 14082 24670 14084 24722
rect 13916 24500 13972 24510
rect 13356 23214 13358 23266
rect 13410 23214 13412 23266
rect 13356 23202 13412 23214
rect 13468 24276 13524 24286
rect 13468 24162 13524 24220
rect 13468 24110 13470 24162
rect 13522 24110 13524 24162
rect 12684 23154 12740 23166
rect 12684 23102 12686 23154
rect 12738 23102 12740 23154
rect 12124 21422 12126 21474
rect 12178 21422 12180 21474
rect 12124 21410 12180 21422
rect 12460 21586 12516 21598
rect 12460 21534 12462 21586
rect 12514 21534 12516 21586
rect 11116 20804 11172 20814
rect 11116 18450 11172 20748
rect 12460 20580 12516 21534
rect 12684 20804 12740 23102
rect 13468 23044 13524 24110
rect 13916 23938 13972 24444
rect 14028 24164 14084 24670
rect 14028 24098 14084 24108
rect 13916 23886 13918 23938
rect 13970 23886 13972 23938
rect 13916 23874 13972 23886
rect 14028 23828 14084 23838
rect 14028 23734 14084 23772
rect 13356 22988 13524 23044
rect 13356 21586 13412 22988
rect 14028 21812 14084 21822
rect 14028 21718 14084 21756
rect 13356 21534 13358 21586
rect 13410 21534 13412 21586
rect 13356 21522 13412 21534
rect 14140 21588 14196 24892
rect 15372 24892 15540 24948
rect 15596 25282 15988 25284
rect 15596 25230 15934 25282
rect 15986 25230 15988 25282
rect 15596 25228 15988 25230
rect 15596 24946 15652 25228
rect 15596 24894 15598 24946
rect 15650 24894 15652 24946
rect 14588 24836 14644 24846
rect 14588 24742 14644 24780
rect 15036 24722 15092 24734
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 14700 24612 14756 24622
rect 14700 24164 14756 24556
rect 14812 24164 14868 24174
rect 14700 24162 14868 24164
rect 14700 24110 14814 24162
rect 14866 24110 14868 24162
rect 14700 24108 14868 24110
rect 14812 24098 14868 24108
rect 14252 23940 14308 23950
rect 14252 23846 14308 23884
rect 14588 23826 14644 23838
rect 14588 23774 14590 23826
rect 14642 23774 14644 23826
rect 14588 23044 14644 23774
rect 15036 23828 15092 24670
rect 15260 24722 15316 24734
rect 15260 24670 15262 24722
rect 15314 24670 15316 24722
rect 15260 24612 15316 24670
rect 15260 24546 15316 24556
rect 15036 23492 15092 23772
rect 15260 23828 15316 23838
rect 15148 23716 15204 23726
rect 15260 23716 15316 23772
rect 15148 23714 15316 23716
rect 15148 23662 15150 23714
rect 15202 23662 15316 23714
rect 15148 23660 15316 23662
rect 15148 23650 15204 23660
rect 15036 23426 15092 23436
rect 14588 22978 14644 22988
rect 14252 21588 14308 21598
rect 14140 21586 14308 21588
rect 14140 21534 14254 21586
rect 14306 21534 14308 21586
rect 14140 21532 14308 21534
rect 13132 21474 13188 21486
rect 13132 21422 13134 21474
rect 13186 21422 13188 21474
rect 12684 20738 12740 20748
rect 12908 20916 12964 20926
rect 13132 20916 13188 21422
rect 12908 20914 13188 20916
rect 12908 20862 12910 20914
rect 12962 20862 13188 20914
rect 12908 20860 13188 20862
rect 13692 21362 13748 21374
rect 13692 21310 13694 21362
rect 13746 21310 13748 21362
rect 12908 20580 12964 20860
rect 12460 20524 12964 20580
rect 12908 20188 12964 20524
rect 13692 20188 13748 21310
rect 14140 20804 14196 20814
rect 14140 20710 14196 20748
rect 14252 20188 14308 21532
rect 14924 20690 14980 20702
rect 14924 20638 14926 20690
rect 14978 20638 14980 20690
rect 14924 20580 14980 20638
rect 14924 20514 14980 20524
rect 15372 20356 15428 24892
rect 15596 24882 15652 24894
rect 15484 24722 15540 24734
rect 15484 24670 15486 24722
rect 15538 24670 15540 24722
rect 15484 24050 15540 24670
rect 15596 24612 15652 24622
rect 15596 24518 15652 24556
rect 15708 24162 15764 25228
rect 15932 25218 15988 25228
rect 16156 24834 16212 25452
rect 16268 25442 16324 25452
rect 16380 25284 16436 26238
rect 16604 26292 16660 26302
rect 16604 26198 16660 26236
rect 16828 26290 16884 26302
rect 16828 26238 16830 26290
rect 16882 26238 16884 26290
rect 16828 25620 16884 26238
rect 16828 25554 16884 25564
rect 16716 25508 16772 25518
rect 16716 25414 16772 25452
rect 16940 25508 16996 25518
rect 16940 25506 17220 25508
rect 16940 25454 16942 25506
rect 16994 25454 17220 25506
rect 16940 25452 17220 25454
rect 16940 25442 16996 25452
rect 16380 25218 16436 25228
rect 16828 25282 16884 25294
rect 16828 25230 16830 25282
rect 16882 25230 16884 25282
rect 16828 25060 16884 25230
rect 16716 25004 16884 25060
rect 17052 25284 17108 25294
rect 16156 24782 16158 24834
rect 16210 24782 16212 24834
rect 16156 24612 16212 24782
rect 16268 24892 16660 24948
rect 16268 24834 16324 24892
rect 16268 24782 16270 24834
rect 16322 24782 16324 24834
rect 16268 24770 16324 24782
rect 16156 24546 16212 24556
rect 16380 24722 16436 24734
rect 16380 24670 16382 24722
rect 16434 24670 16436 24722
rect 15708 24110 15710 24162
rect 15762 24110 15764 24162
rect 15708 24098 15764 24110
rect 15484 23998 15486 24050
rect 15538 23998 15540 24050
rect 15484 23940 15540 23998
rect 16044 24050 16100 24062
rect 16044 23998 16046 24050
rect 16098 23998 16100 24050
rect 16044 23940 16100 23998
rect 16380 23940 16436 24670
rect 16044 23938 16436 23940
rect 16044 23886 16382 23938
rect 16434 23886 16436 23938
rect 16044 23884 16436 23886
rect 15484 23874 15540 23884
rect 16380 23874 16436 23884
rect 16492 24164 16548 24174
rect 15820 23492 15876 23502
rect 15820 23378 15876 23436
rect 15820 23326 15822 23378
rect 15874 23326 15876 23378
rect 15820 23314 15876 23326
rect 16492 23378 16548 24108
rect 16492 23326 16494 23378
rect 16546 23326 16548 23378
rect 16492 23314 16548 23326
rect 16604 23828 16660 24892
rect 16604 23266 16660 23772
rect 16716 23826 16772 25004
rect 16828 24836 16884 24846
rect 17052 24836 17108 25228
rect 16828 24834 17108 24836
rect 16828 24782 16830 24834
rect 16882 24782 17108 24834
rect 16828 24780 17108 24782
rect 16828 24770 16884 24780
rect 17164 24164 17220 25452
rect 17276 24948 17332 32060
rect 17500 31892 17556 32622
rect 17612 32674 17668 33180
rect 17612 32622 17614 32674
rect 17666 32622 17668 32674
rect 17612 32228 17668 32622
rect 17612 32162 17668 32172
rect 17724 33124 17780 33134
rect 17500 31826 17556 31836
rect 17500 31666 17556 31678
rect 17500 31614 17502 31666
rect 17554 31614 17556 31666
rect 17388 31220 17444 31230
rect 17388 31126 17444 31164
rect 17500 30324 17556 31614
rect 17612 31220 17668 31230
rect 17724 31220 17780 33068
rect 17612 31218 17780 31220
rect 17612 31166 17614 31218
rect 17666 31166 17780 31218
rect 17612 31164 17780 31166
rect 17612 31154 17668 31164
rect 17724 31108 17780 31164
rect 17724 31042 17780 31052
rect 17836 32004 17892 33516
rect 18620 33460 18676 33470
rect 18620 33458 18900 33460
rect 18620 33406 18622 33458
rect 18674 33406 18900 33458
rect 18620 33404 18900 33406
rect 18620 33394 18676 33404
rect 18172 33348 18228 33358
rect 18172 33254 18228 33292
rect 18060 33124 18116 33134
rect 18284 33124 18340 33134
rect 18060 32674 18116 33068
rect 18060 32622 18062 32674
rect 18114 32622 18116 32674
rect 18060 32610 18116 32622
rect 18172 33068 18284 33124
rect 17836 31106 17892 31948
rect 18060 32228 18116 32238
rect 18060 31218 18116 32172
rect 18172 32116 18228 33068
rect 18284 33030 18340 33068
rect 18508 33122 18564 33134
rect 18508 33070 18510 33122
rect 18562 33070 18564 33122
rect 18508 32788 18564 33070
rect 18620 33124 18676 33134
rect 18620 33122 18788 33124
rect 18620 33070 18622 33122
rect 18674 33070 18788 33122
rect 18620 33068 18788 33070
rect 18620 33058 18676 33068
rect 18508 32722 18564 32732
rect 18732 32788 18788 33068
rect 18732 32722 18788 32732
rect 18620 32676 18676 32686
rect 18172 32050 18228 32060
rect 18284 32562 18340 32574
rect 18284 32510 18286 32562
rect 18338 32510 18340 32562
rect 18060 31166 18062 31218
rect 18114 31166 18116 31218
rect 18060 31154 18116 31166
rect 18172 31780 18228 31790
rect 17836 31054 17838 31106
rect 17890 31054 17892 31106
rect 17836 31042 17892 31054
rect 17724 30772 17780 30782
rect 17724 30678 17780 30716
rect 17500 29426 17556 30268
rect 18172 30100 18228 31724
rect 18284 31444 18340 32510
rect 18508 32562 18564 32574
rect 18508 32510 18510 32562
rect 18562 32510 18564 32562
rect 18284 31378 18340 31388
rect 18396 32004 18452 32014
rect 18284 31108 18340 31118
rect 18284 31014 18340 31052
rect 18396 31106 18452 31948
rect 18508 31220 18564 32510
rect 18620 32450 18676 32620
rect 18620 32398 18622 32450
rect 18674 32398 18676 32450
rect 18620 32386 18676 32398
rect 18732 32562 18788 32574
rect 18732 32510 18734 32562
rect 18786 32510 18788 32562
rect 18508 31154 18564 31164
rect 18732 31218 18788 32510
rect 18844 32564 18900 33404
rect 18956 32676 19012 33516
rect 19068 33124 19124 33134
rect 19068 33030 19124 33068
rect 18956 32610 19012 32620
rect 19068 32788 19124 32798
rect 19180 32788 19236 33852
rect 19292 33458 19348 33966
rect 20412 34020 20468 34030
rect 20468 33964 20580 34020
rect 20412 33926 20468 33964
rect 19516 33906 19572 33918
rect 19516 33854 19518 33906
rect 19570 33854 19572 33906
rect 19292 33406 19294 33458
rect 19346 33406 19348 33458
rect 19292 33394 19348 33406
rect 19404 33460 19460 33470
rect 19292 33236 19348 33246
rect 19292 33142 19348 33180
rect 19404 33234 19460 33404
rect 19404 33182 19406 33234
rect 19458 33182 19460 33234
rect 19404 33170 19460 33182
rect 19404 33012 19460 33022
rect 19292 32788 19348 32798
rect 19180 32786 19348 32788
rect 19180 32734 19294 32786
rect 19346 32734 19348 32786
rect 19180 32732 19348 32734
rect 18844 32498 18900 32508
rect 18732 31166 18734 31218
rect 18786 31166 18788 31218
rect 18732 31154 18788 31166
rect 18956 31556 19012 31566
rect 18396 31054 18398 31106
rect 18450 31054 18452 31106
rect 18396 31042 18452 31054
rect 18844 30884 18900 30894
rect 18844 30790 18900 30828
rect 18620 30772 18676 30782
rect 18396 30100 18452 30110
rect 18172 30044 18396 30100
rect 18396 30006 18452 30044
rect 17500 29374 17502 29426
rect 17554 29374 17556 29426
rect 17500 29362 17556 29374
rect 18172 29316 18228 29326
rect 18172 29314 18452 29316
rect 18172 29262 18174 29314
rect 18226 29262 18452 29314
rect 18172 29260 18452 29262
rect 18172 29250 18228 29260
rect 17724 28530 17780 28542
rect 17724 28478 17726 28530
rect 17778 28478 17780 28530
rect 17724 28420 17780 28478
rect 17836 28532 17892 28542
rect 17836 28438 17892 28476
rect 18284 28530 18340 28542
rect 18284 28478 18286 28530
rect 18338 28478 18340 28530
rect 17724 28354 17780 28364
rect 18060 28418 18116 28430
rect 18060 28366 18062 28418
rect 18114 28366 18116 28418
rect 17500 27972 17556 27982
rect 17500 27970 17780 27972
rect 17500 27918 17502 27970
rect 17554 27918 17780 27970
rect 17500 27916 17780 27918
rect 17500 27906 17556 27916
rect 17388 27860 17444 27870
rect 17388 27766 17444 27804
rect 17500 27634 17556 27646
rect 17500 27582 17502 27634
rect 17554 27582 17556 27634
rect 17388 27300 17444 27310
rect 17500 27300 17556 27582
rect 17612 27300 17668 27310
rect 17500 27298 17668 27300
rect 17500 27246 17614 27298
rect 17666 27246 17668 27298
rect 17500 27244 17668 27246
rect 17388 27206 17444 27244
rect 17612 27234 17668 27244
rect 17388 26852 17444 26862
rect 17388 26402 17444 26796
rect 17612 26516 17668 26526
rect 17724 26516 17780 27916
rect 17948 27860 18004 27870
rect 17836 27858 18004 27860
rect 17836 27806 17950 27858
rect 18002 27806 18004 27858
rect 17836 27804 18004 27806
rect 17836 26852 17892 27804
rect 17948 27794 18004 27804
rect 17836 26786 17892 26796
rect 17948 27636 18004 27646
rect 17668 26460 17780 26516
rect 17612 26422 17668 26460
rect 17388 26350 17390 26402
rect 17442 26350 17444 26402
rect 17388 26338 17444 26350
rect 17836 26404 17892 26414
rect 17836 26310 17892 26348
rect 17500 26292 17556 26302
rect 17500 25506 17556 26236
rect 17500 25454 17502 25506
rect 17554 25454 17556 25506
rect 17500 25442 17556 25454
rect 17724 26178 17780 26190
rect 17724 26126 17726 26178
rect 17778 26126 17780 26178
rect 17724 25508 17780 26126
rect 17948 26068 18004 27580
rect 18060 27076 18116 28366
rect 18172 27860 18228 27870
rect 18172 27766 18228 27804
rect 18284 27524 18340 28478
rect 18396 28082 18452 29260
rect 18396 28030 18398 28082
rect 18450 28030 18452 28082
rect 18396 28018 18452 28030
rect 18508 28418 18564 28430
rect 18508 28366 18510 28418
rect 18562 28366 18564 28418
rect 18396 27636 18452 27646
rect 18396 27542 18452 27580
rect 18284 27458 18340 27468
rect 18060 27010 18116 27020
rect 18284 27300 18340 27310
rect 18508 27300 18564 28366
rect 18620 27970 18676 30716
rect 18620 27918 18622 27970
rect 18674 27918 18676 27970
rect 18620 27906 18676 27918
rect 18732 28642 18788 28654
rect 18732 28590 18734 28642
rect 18786 28590 18788 28642
rect 18732 28308 18788 28590
rect 18284 27074 18340 27244
rect 18284 27022 18286 27074
rect 18338 27022 18340 27074
rect 18284 27010 18340 27022
rect 18396 27244 18564 27300
rect 18620 27412 18676 27422
rect 18060 26852 18116 26862
rect 18060 26850 18228 26852
rect 18060 26798 18062 26850
rect 18114 26798 18228 26850
rect 18060 26796 18228 26798
rect 18060 26786 18116 26796
rect 18172 26516 18228 26796
rect 18396 26628 18452 27244
rect 18620 27186 18676 27356
rect 18620 27134 18622 27186
rect 18674 27134 18676 27186
rect 18620 27122 18676 27134
rect 18508 27076 18564 27086
rect 18508 26962 18564 27020
rect 18732 27074 18788 28252
rect 18956 27858 19012 31500
rect 19068 30884 19124 32732
rect 19292 32722 19348 32732
rect 19404 32786 19460 32956
rect 19404 32734 19406 32786
rect 19458 32734 19460 32786
rect 19404 32722 19460 32734
rect 19516 32788 19572 33854
rect 20188 33460 20244 33470
rect 20188 33346 20244 33404
rect 20188 33294 20190 33346
rect 20242 33294 20244 33346
rect 19516 32722 19572 32732
rect 19628 33234 19684 33246
rect 19628 33182 19630 33234
rect 19682 33182 19684 33234
rect 19628 32788 19684 33182
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19740 32788 19796 32798
rect 19628 32786 19796 32788
rect 19628 32734 19742 32786
rect 19794 32734 19796 32786
rect 19628 32732 19796 32734
rect 19516 32564 19572 32574
rect 19516 32470 19572 32508
rect 19180 31892 19236 31902
rect 19180 31778 19236 31836
rect 19628 31890 19684 32732
rect 19740 32722 19796 32732
rect 20076 32788 20132 32798
rect 20076 32694 20132 32732
rect 20188 32002 20244 33294
rect 20412 33346 20468 33358
rect 20412 33294 20414 33346
rect 20466 33294 20468 33346
rect 20412 33124 20468 33294
rect 20412 33058 20468 33068
rect 20300 32674 20356 32686
rect 20300 32622 20302 32674
rect 20354 32622 20356 32674
rect 20300 32564 20356 32622
rect 20412 32676 20468 32686
rect 20412 32582 20468 32620
rect 20300 32498 20356 32508
rect 20524 32116 20580 33964
rect 20188 31950 20190 32002
rect 20242 31950 20244 32002
rect 20188 31938 20244 31950
rect 20412 32060 20580 32116
rect 19628 31838 19630 31890
rect 19682 31838 19684 31890
rect 19628 31826 19684 31838
rect 19180 31726 19182 31778
rect 19234 31726 19236 31778
rect 19180 31714 19236 31726
rect 19404 31780 19460 31790
rect 19404 31554 19460 31724
rect 19852 31778 19908 31790
rect 19852 31726 19854 31778
rect 19906 31726 19908 31778
rect 19852 31668 19908 31726
rect 20412 31780 20468 32060
rect 20412 31714 20468 31724
rect 20524 31778 20580 31790
rect 20524 31726 20526 31778
rect 20578 31726 20580 31778
rect 19852 31602 19908 31612
rect 20524 31668 20580 31726
rect 19404 31502 19406 31554
rect 19458 31502 19460 31554
rect 19180 31444 19236 31454
rect 19180 31218 19236 31388
rect 19404 31332 19460 31502
rect 19628 31556 19684 31566
rect 19628 31462 19684 31500
rect 20188 31444 20244 31454
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19404 31276 19684 31332
rect 19836 31322 20100 31332
rect 19180 31166 19182 31218
rect 19234 31166 19236 31218
rect 19180 31154 19236 31166
rect 19292 30884 19348 30894
rect 19628 30884 19684 31276
rect 19068 30882 19572 30884
rect 19068 30830 19294 30882
rect 19346 30830 19572 30882
rect 19068 30828 19572 30830
rect 19292 30818 19348 30828
rect 19404 29652 19460 29662
rect 19404 28644 19460 29596
rect 18956 27806 18958 27858
rect 19010 27806 19012 27858
rect 18956 27794 19012 27806
rect 19180 28642 19460 28644
rect 19180 28590 19406 28642
rect 19458 28590 19460 28642
rect 19180 28588 19460 28590
rect 19180 28532 19236 28588
rect 19404 28578 19460 28588
rect 19180 27858 19236 28476
rect 19404 28420 19460 28430
rect 19180 27806 19182 27858
rect 19234 27806 19236 27858
rect 19180 27794 19236 27806
rect 19292 27972 19348 27982
rect 19292 27636 19348 27916
rect 19404 27858 19460 28364
rect 19404 27806 19406 27858
rect 19458 27806 19460 27858
rect 19404 27794 19460 27806
rect 19292 27580 19460 27636
rect 19180 27524 19236 27534
rect 19236 27468 19348 27524
rect 19180 27458 19236 27468
rect 18732 27022 18734 27074
rect 18786 27022 18788 27074
rect 18732 27010 18788 27022
rect 18956 27074 19012 27086
rect 18956 27022 18958 27074
rect 19010 27022 19012 27074
rect 18508 26910 18510 26962
rect 18562 26910 18564 26962
rect 18508 26898 18564 26910
rect 18956 26964 19012 27022
rect 19292 27074 19348 27468
rect 19404 27186 19460 27580
rect 19404 27134 19406 27186
rect 19458 27134 19460 27186
rect 19404 27122 19460 27134
rect 19292 27022 19294 27074
rect 19346 27022 19348 27074
rect 19292 26964 19348 27022
rect 18956 26908 19348 26964
rect 19292 26628 19348 26638
rect 18396 26572 18788 26628
rect 18172 26460 18676 26516
rect 18060 26292 18116 26302
rect 18396 26292 18452 26302
rect 18060 26290 18452 26292
rect 18060 26238 18062 26290
rect 18114 26238 18398 26290
rect 18450 26238 18452 26290
rect 18060 26236 18452 26238
rect 18060 26226 18116 26236
rect 18396 26226 18452 26236
rect 18508 26178 18564 26190
rect 18508 26126 18510 26178
rect 18562 26126 18564 26178
rect 17948 26012 18116 26068
rect 17948 25620 18004 25630
rect 17948 25526 18004 25564
rect 17724 25442 17780 25452
rect 17836 25172 17892 25182
rect 17276 24892 17444 24948
rect 17164 24098 17220 24108
rect 17052 24052 17108 24062
rect 17052 23958 17108 23996
rect 16716 23774 16718 23826
rect 16770 23774 16772 23826
rect 16716 23762 16772 23774
rect 16604 23214 16606 23266
rect 16658 23214 16660 23266
rect 16604 23202 16660 23214
rect 16044 23154 16100 23166
rect 16044 23102 16046 23154
rect 16098 23102 16100 23154
rect 15484 23044 15540 23054
rect 15484 22950 15540 22988
rect 16044 23044 16100 23102
rect 16044 22978 16100 22988
rect 17276 22932 17332 22942
rect 17052 22596 17108 22606
rect 17052 22482 17108 22540
rect 17052 22430 17054 22482
rect 17106 22430 17108 22482
rect 17052 22418 17108 22430
rect 17276 22482 17332 22876
rect 17276 22430 17278 22482
rect 17330 22430 17332 22482
rect 17276 22418 17332 22430
rect 16044 21588 16100 21598
rect 16044 21494 16100 21532
rect 16492 21476 16548 21486
rect 16492 21382 16548 21420
rect 16828 21474 16884 21486
rect 16828 21422 16830 21474
rect 16882 21422 16884 21474
rect 16828 21252 16884 21422
rect 17388 21474 17444 24892
rect 17836 24836 17892 25116
rect 17836 24050 17892 24780
rect 18060 24500 18116 26012
rect 18508 25620 18564 26126
rect 18508 25554 18564 25564
rect 18396 25508 18452 25518
rect 18172 25394 18228 25406
rect 18172 25342 18174 25394
rect 18226 25342 18228 25394
rect 18172 24722 18228 25342
rect 18284 25394 18340 25406
rect 18284 25342 18286 25394
rect 18338 25342 18340 25394
rect 18284 25284 18340 25342
rect 18284 25218 18340 25228
rect 18172 24670 18174 24722
rect 18226 24670 18228 24722
rect 18172 24658 18228 24670
rect 18060 24444 18340 24500
rect 17836 23998 17838 24050
rect 17890 23998 17892 24050
rect 17836 23986 17892 23998
rect 17388 21422 17390 21474
rect 17442 21422 17444 21474
rect 17388 21364 17444 21422
rect 17388 21298 17444 21308
rect 17500 23940 17556 23950
rect 16828 21186 16884 21196
rect 17052 20914 17108 20926
rect 17052 20862 17054 20914
rect 17106 20862 17108 20914
rect 17052 20804 17108 20862
rect 17052 20738 17108 20748
rect 17388 20802 17444 20814
rect 17388 20750 17390 20802
rect 17442 20750 17444 20802
rect 16604 20692 16660 20702
rect 15372 20290 15428 20300
rect 16044 20300 16436 20356
rect 16044 20188 16100 20300
rect 12908 20132 13524 20188
rect 13692 20132 13860 20188
rect 13468 20130 13524 20132
rect 13468 20078 13470 20130
rect 13522 20078 13524 20130
rect 13468 20066 13524 20078
rect 13804 20066 13860 20076
rect 14140 20132 14196 20142
rect 14252 20132 14756 20188
rect 15372 20132 15428 20142
rect 13692 20020 13748 20030
rect 12796 19796 12852 19806
rect 12124 19122 12180 19134
rect 12124 19070 12126 19122
rect 12178 19070 12180 19122
rect 11788 19010 11844 19022
rect 11788 18958 11790 19010
rect 11842 18958 11844 19010
rect 11788 18562 11844 18958
rect 12124 19012 12180 19070
rect 12684 19012 12740 19022
rect 12124 18946 12180 18956
rect 12572 19010 12740 19012
rect 12572 18958 12686 19010
rect 12738 18958 12740 19010
rect 12572 18956 12740 18958
rect 11788 18510 11790 18562
rect 11842 18510 11844 18562
rect 11788 18498 11844 18510
rect 11116 18398 11118 18450
rect 11170 18398 11172 18450
rect 11116 17780 11172 18398
rect 11116 17714 11172 17724
rect 11116 17554 11172 17566
rect 11116 17502 11118 17554
rect 11170 17502 11172 17554
rect 11116 15988 11172 17502
rect 11900 17556 11956 17566
rect 11900 17554 12516 17556
rect 11900 17502 11902 17554
rect 11954 17502 12516 17554
rect 11900 17500 12516 17502
rect 11900 17490 11956 17500
rect 11228 17444 11284 17454
rect 11228 17350 11284 17388
rect 11452 17442 11508 17454
rect 11452 17390 11454 17442
rect 11506 17390 11508 17442
rect 11228 16324 11284 16334
rect 11228 16098 11284 16268
rect 11228 16046 11230 16098
rect 11282 16046 11284 16098
rect 11228 16034 11284 16046
rect 11116 15922 11172 15932
rect 11452 15876 11508 17390
rect 11564 17442 11620 17454
rect 11564 17390 11566 17442
rect 11618 17390 11620 17442
rect 11564 16098 11620 17390
rect 11788 17442 11844 17454
rect 11788 17390 11790 17442
rect 11842 17390 11844 17442
rect 11788 17108 11844 17390
rect 11788 17052 12404 17108
rect 12236 16884 12292 16894
rect 11676 16882 12292 16884
rect 11676 16830 12238 16882
rect 12290 16830 12292 16882
rect 11676 16828 12292 16830
rect 11676 16210 11732 16828
rect 12236 16818 12292 16828
rect 12348 16548 12404 17052
rect 12348 16482 12404 16492
rect 11676 16158 11678 16210
rect 11730 16158 11732 16210
rect 11676 16146 11732 16158
rect 11564 16046 11566 16098
rect 11618 16046 11620 16098
rect 11564 16034 11620 16046
rect 11788 16098 11844 16110
rect 11788 16046 11790 16098
rect 11842 16046 11844 16098
rect 11788 15876 11844 16046
rect 11452 15820 11844 15876
rect 12124 15986 12180 15998
rect 12124 15934 12126 15986
rect 12178 15934 12180 15986
rect 12124 15764 12180 15934
rect 11788 15092 11844 15102
rect 11116 14196 11172 14206
rect 11116 13746 11172 14140
rect 11564 13860 11620 13870
rect 11116 13694 11118 13746
rect 11170 13694 11172 13746
rect 11116 13682 11172 13694
rect 11340 13804 11564 13860
rect 11116 13300 11172 13310
rect 11116 13074 11172 13244
rect 11340 13186 11396 13804
rect 11564 13766 11620 13804
rect 11340 13134 11342 13186
rect 11394 13134 11396 13186
rect 11340 13122 11396 13134
rect 11116 13022 11118 13074
rect 11170 13022 11172 13074
rect 11116 13010 11172 13022
rect 11676 12964 11732 12974
rect 11676 12870 11732 12908
rect 11564 12066 11620 12078
rect 11564 12014 11566 12066
rect 11618 12014 11620 12066
rect 11340 11618 11396 11630
rect 11340 11566 11342 11618
rect 11394 11566 11396 11618
rect 11340 11506 11396 11566
rect 11340 11454 11342 11506
rect 11394 11454 11396 11506
rect 11340 11442 11396 11454
rect 11564 11284 11620 12014
rect 11788 11508 11844 15036
rect 12124 14196 12180 15708
rect 12124 14130 12180 14140
rect 12460 14532 12516 17500
rect 12572 16884 12628 18956
rect 12684 18946 12740 18956
rect 12684 17668 12740 17678
rect 12796 17668 12852 19740
rect 13580 19794 13636 19806
rect 13580 19742 13582 19794
rect 13634 19742 13636 19794
rect 13580 18676 13636 19742
rect 13692 19234 13748 19964
rect 13916 19796 13972 19806
rect 13916 19702 13972 19740
rect 13692 19182 13694 19234
rect 13746 19182 13748 19234
rect 13692 19170 13748 19182
rect 14028 19236 14084 19246
rect 14028 19142 14084 19180
rect 13804 19124 13860 19134
rect 13804 19030 13860 19068
rect 13580 18610 13636 18620
rect 13916 18564 13972 18574
rect 13916 18338 13972 18508
rect 14140 18452 14196 20076
rect 14364 20020 14420 20030
rect 14364 19926 14420 19964
rect 14476 20018 14532 20030
rect 14476 19966 14478 20018
rect 14530 19966 14532 20018
rect 14252 19012 14308 19022
rect 14252 18918 14308 18956
rect 14476 18788 14532 19966
rect 14700 20020 14756 20132
rect 15148 20130 15428 20132
rect 15148 20078 15374 20130
rect 15426 20078 15428 20130
rect 15148 20076 15428 20078
rect 14700 20018 14980 20020
rect 14700 19966 14702 20018
rect 14754 19966 14980 20018
rect 14700 19964 14980 19966
rect 14700 19954 14756 19964
rect 14700 19684 14756 19694
rect 14700 19234 14756 19628
rect 14700 19182 14702 19234
rect 14754 19182 14756 19234
rect 14700 19170 14756 19182
rect 14812 19236 14868 19246
rect 14812 19142 14868 19180
rect 14924 19234 14980 19964
rect 14924 19182 14926 19234
rect 14978 19182 14980 19234
rect 14924 19170 14980 19182
rect 15148 19908 15204 20076
rect 15372 20066 15428 20076
rect 15932 20132 16100 20188
rect 16268 20132 16324 20142
rect 15596 20020 15652 20030
rect 15484 20018 15652 20020
rect 15484 19966 15598 20018
rect 15650 19966 15652 20018
rect 15484 19964 15652 19966
rect 14252 18732 14532 18788
rect 14252 18674 14308 18732
rect 14252 18622 14254 18674
rect 14306 18622 14308 18674
rect 14252 18610 14308 18622
rect 15148 18564 15204 19852
rect 15372 19906 15428 19918
rect 15372 19854 15374 19906
rect 15426 19854 15428 19906
rect 15372 19684 15428 19854
rect 15372 19618 15428 19628
rect 15484 19796 15540 19964
rect 15596 19954 15652 19964
rect 15932 20018 15988 20076
rect 16156 20130 16324 20132
rect 16156 20078 16270 20130
rect 16322 20078 16324 20130
rect 16156 20076 16324 20078
rect 15932 19966 15934 20018
rect 15986 19966 15988 20018
rect 15932 19954 15988 19966
rect 16044 20020 16100 20030
rect 16044 19926 16100 19964
rect 15484 19460 15540 19740
rect 16044 19796 16100 19806
rect 16156 19796 16212 20076
rect 16268 20066 16324 20076
rect 16380 20130 16436 20300
rect 16380 20078 16382 20130
rect 16434 20078 16436 20130
rect 16380 20066 16436 20078
rect 16100 19740 16212 19796
rect 16268 19796 16324 19806
rect 16044 19730 16100 19740
rect 15148 18498 15204 18508
rect 15260 19404 15540 19460
rect 14588 18452 14644 18462
rect 14140 18450 14644 18452
rect 14140 18398 14590 18450
rect 14642 18398 14644 18450
rect 14140 18396 14644 18398
rect 14588 18386 14644 18396
rect 14812 18452 14868 18462
rect 14812 18358 14868 18396
rect 15260 18452 15316 19404
rect 16268 19124 16324 19740
rect 15708 18564 15764 18574
rect 15596 18508 15708 18564
rect 13916 18286 13918 18338
rect 13970 18286 13972 18338
rect 13916 18274 13972 18286
rect 15036 18340 15092 18350
rect 12908 17780 12964 17790
rect 13692 17780 13748 17790
rect 12964 17724 13076 17780
rect 12908 17714 12964 17724
rect 12684 17666 12852 17668
rect 12684 17614 12686 17666
rect 12738 17614 12852 17666
rect 12684 17612 12852 17614
rect 12684 17602 12740 17612
rect 12908 17444 12964 17454
rect 12908 17350 12964 17388
rect 13020 16884 13076 17724
rect 13748 17724 13972 17780
rect 13692 17686 13748 17724
rect 13356 16884 13412 16894
rect 12572 16828 12964 16884
rect 12796 16548 12852 16558
rect 11900 13972 11956 13982
rect 11900 13878 11956 13916
rect 12460 13858 12516 14476
rect 12572 16324 12628 16334
rect 12572 13970 12628 16268
rect 12572 13918 12574 13970
rect 12626 13918 12628 13970
rect 12572 13906 12628 13918
rect 12684 15988 12740 15998
rect 12684 13972 12740 15932
rect 12796 15986 12852 16492
rect 12796 15934 12798 15986
rect 12850 15934 12852 15986
rect 12796 15922 12852 15934
rect 12796 15764 12852 15774
rect 12908 15764 12964 16828
rect 13020 16882 13412 16884
rect 13020 16830 13022 16882
rect 13074 16830 13358 16882
rect 13410 16830 13412 16882
rect 13020 16828 13412 16830
rect 13020 16818 13076 16828
rect 13356 16818 13412 16828
rect 13356 16100 13412 16110
rect 13132 16098 13412 16100
rect 13132 16046 13358 16098
rect 13410 16046 13412 16098
rect 13132 16044 13412 16046
rect 13020 15988 13076 15998
rect 13020 15894 13076 15932
rect 12852 15708 12964 15764
rect 12796 15698 12852 15708
rect 13132 15148 13188 16044
rect 13356 16034 13412 16044
rect 13692 16098 13748 16110
rect 13692 16046 13694 16098
rect 13746 16046 13748 16098
rect 13692 15988 13748 16046
rect 13692 15922 13748 15932
rect 13580 15874 13636 15886
rect 13580 15822 13582 15874
rect 13634 15822 13636 15874
rect 13580 15316 13636 15822
rect 13804 15764 13860 15774
rect 13580 15250 13636 15260
rect 13692 15708 13804 15764
rect 13692 15148 13748 15708
rect 13804 15698 13860 15708
rect 12684 13906 12740 13916
rect 12796 15092 13188 15148
rect 13580 15092 13748 15148
rect 12796 13970 12852 15092
rect 12908 14644 12964 14654
rect 12908 14550 12964 14588
rect 13580 14642 13636 15092
rect 13580 14590 13582 14642
rect 13634 14590 13636 14642
rect 13580 14578 13636 14590
rect 13916 14530 13972 17724
rect 14140 17444 14196 17454
rect 14140 16994 14196 17388
rect 14140 16942 14142 16994
rect 14194 16942 14196 16994
rect 14140 16930 14196 16942
rect 14028 15986 14084 15998
rect 14028 15934 14030 15986
rect 14082 15934 14084 15986
rect 14028 15764 14084 15934
rect 14476 15876 14532 15886
rect 14028 15698 14084 15708
rect 14364 15820 14476 15876
rect 14252 15428 14308 15438
rect 14364 15428 14420 15820
rect 14476 15782 14532 15820
rect 14812 15874 14868 15886
rect 14812 15822 14814 15874
rect 14866 15822 14868 15874
rect 14812 15764 14868 15822
rect 14812 15698 14868 15708
rect 14308 15372 14420 15428
rect 15036 15540 15092 18284
rect 15260 17444 15316 18396
rect 15372 18450 15428 18462
rect 15372 18398 15374 18450
rect 15426 18398 15428 18450
rect 15372 17668 15428 18398
rect 15596 18450 15652 18508
rect 15708 18498 15764 18508
rect 15596 18398 15598 18450
rect 15650 18398 15652 18450
rect 15596 18386 15652 18398
rect 15820 18450 15876 18462
rect 15820 18398 15822 18450
rect 15874 18398 15876 18450
rect 15708 18338 15764 18350
rect 15708 18286 15710 18338
rect 15762 18286 15764 18338
rect 15708 18004 15764 18286
rect 15820 18228 15876 18398
rect 16268 18450 16324 19068
rect 16604 18674 16660 20636
rect 17388 20692 17444 20750
rect 17388 20626 17444 20636
rect 16828 19908 16884 19918
rect 16828 19814 16884 19852
rect 17500 19906 17556 23884
rect 18060 23042 18116 23054
rect 18060 22990 18062 23042
rect 18114 22990 18116 23042
rect 17948 21252 18004 21262
rect 17948 21026 18004 21196
rect 17948 20974 17950 21026
rect 18002 20974 18004 21026
rect 17948 20962 18004 20974
rect 17500 19854 17502 19906
rect 17554 19854 17556 19906
rect 17500 19842 17556 19854
rect 17724 20690 17780 20702
rect 17724 20638 17726 20690
rect 17778 20638 17780 20690
rect 16716 19796 16772 19806
rect 16716 19702 16772 19740
rect 17724 19684 17780 20638
rect 17836 20580 17892 20590
rect 17836 20486 17892 20524
rect 18060 20188 18116 22990
rect 18172 20916 18228 20926
rect 18172 20822 18228 20860
rect 17948 20132 18116 20188
rect 17724 19618 17780 19628
rect 17836 19794 17892 19806
rect 17836 19742 17838 19794
rect 17890 19742 17892 19794
rect 16604 18622 16606 18674
rect 16658 18622 16660 18674
rect 16604 18610 16660 18622
rect 17052 18844 17444 18900
rect 16268 18398 16270 18450
rect 16322 18398 16324 18450
rect 16268 18386 16324 18398
rect 16380 18450 16436 18462
rect 16380 18398 16382 18450
rect 16434 18398 16436 18450
rect 15820 18162 15876 18172
rect 15708 17938 15764 17948
rect 16380 17892 16436 18398
rect 16492 18452 16548 18462
rect 16492 18358 16548 18396
rect 16828 18450 16884 18462
rect 16828 18398 16830 18450
rect 16882 18398 16884 18450
rect 16380 17826 16436 17836
rect 16828 17780 16884 18398
rect 16828 17714 16884 17724
rect 15372 17602 15428 17612
rect 16492 17668 16548 17678
rect 16548 17612 16772 17668
rect 16492 17602 16548 17612
rect 15260 17388 15652 17444
rect 15484 15988 15540 15998
rect 15596 15988 15652 17388
rect 16716 17106 16772 17612
rect 16716 17054 16718 17106
rect 16770 17054 16772 17106
rect 16716 17042 16772 17054
rect 16828 16884 16884 16894
rect 16268 16770 16324 16782
rect 16268 16718 16270 16770
rect 16322 16718 16324 16770
rect 15820 15988 15876 15998
rect 15596 15986 15876 15988
rect 15596 15934 15822 15986
rect 15874 15934 15876 15986
rect 15596 15932 15876 15934
rect 15484 15894 15540 15932
rect 15820 15922 15876 15932
rect 16156 15988 16212 15998
rect 16268 15988 16324 16718
rect 16828 16098 16884 16828
rect 17052 16548 17108 18844
rect 17276 18676 17332 18686
rect 17164 18620 17276 18676
rect 17164 16660 17220 18620
rect 17276 18610 17332 18620
rect 17388 18674 17444 18844
rect 17388 18622 17390 18674
rect 17442 18622 17444 18674
rect 17388 18610 17444 18622
rect 17612 18676 17668 18686
rect 17612 18582 17668 18620
rect 17500 18564 17556 18574
rect 17388 18004 17444 18014
rect 17388 16996 17444 17948
rect 17500 17556 17556 18508
rect 17724 18562 17780 18574
rect 17724 18510 17726 18562
rect 17778 18510 17780 18562
rect 17724 18116 17780 18510
rect 17836 18340 17892 19742
rect 17836 18274 17892 18284
rect 17836 18116 17892 18126
rect 17724 18060 17836 18116
rect 17836 18050 17892 18060
rect 17500 17500 17892 17556
rect 17836 17106 17892 17500
rect 17836 17054 17838 17106
rect 17890 17054 17892 17106
rect 17836 17042 17892 17054
rect 17724 16996 17780 17006
rect 17388 16994 17780 16996
rect 17388 16942 17726 16994
rect 17778 16942 17780 16994
rect 17388 16940 17780 16942
rect 17724 16930 17780 16940
rect 17164 16604 17444 16660
rect 17052 16492 17332 16548
rect 17164 16212 17220 16222
rect 17164 16118 17220 16156
rect 16828 16046 16830 16098
rect 16882 16046 16884 16098
rect 16828 16034 16884 16046
rect 17276 16100 17332 16492
rect 17276 16006 17332 16044
rect 17388 16098 17444 16604
rect 17388 16046 17390 16098
rect 17442 16046 17444 16098
rect 17388 16034 17444 16046
rect 17836 16210 17892 16222
rect 17836 16158 17838 16210
rect 17890 16158 17892 16210
rect 17836 16100 17892 16158
rect 17836 16034 17892 16044
rect 16156 15986 16324 15988
rect 16156 15934 16158 15986
rect 16210 15934 16324 15986
rect 16156 15932 16324 15934
rect 17612 15988 17668 15998
rect 15148 15876 15204 15886
rect 15148 15782 15204 15820
rect 14252 15362 14308 15372
rect 14476 15316 14532 15326
rect 14532 15260 14756 15316
rect 14476 15250 14532 15260
rect 14140 15204 14196 15214
rect 13916 14478 13918 14530
rect 13970 14478 13972 14530
rect 13916 14466 13972 14478
rect 14028 15148 14140 15204
rect 12796 13918 12798 13970
rect 12850 13918 12852 13970
rect 12796 13906 12852 13918
rect 12460 13806 12462 13858
rect 12514 13806 12516 13858
rect 12460 13794 12516 13806
rect 13916 13860 13972 13870
rect 14028 13860 14084 15148
rect 14140 15138 14196 15148
rect 13916 13858 14084 13860
rect 13916 13806 13918 13858
rect 13970 13806 14084 13858
rect 13916 13804 14084 13806
rect 14140 14644 14196 14654
rect 13916 13794 13972 13804
rect 13244 13746 13300 13758
rect 13244 13694 13246 13746
rect 13298 13694 13300 13746
rect 12124 13412 12180 13422
rect 11900 13076 11956 13086
rect 11900 12982 11956 13020
rect 12124 12962 12180 13356
rect 12124 12910 12126 12962
rect 12178 12910 12180 12962
rect 12124 12898 12180 12910
rect 12348 13412 12404 13422
rect 12348 13076 12404 13356
rect 12348 12850 12404 13020
rect 12460 12964 12516 12974
rect 12796 12964 12852 12974
rect 12516 12962 12852 12964
rect 12516 12910 12798 12962
rect 12850 12910 12852 12962
rect 12516 12908 12852 12910
rect 12460 12870 12516 12908
rect 12796 12898 12852 12908
rect 13244 12964 13300 13694
rect 14028 13412 14084 13422
rect 14028 13074 14084 13356
rect 14028 13022 14030 13074
rect 14082 13022 14084 13074
rect 14028 13010 14084 13022
rect 13244 12898 13300 12908
rect 13804 12962 13860 12974
rect 13804 12910 13806 12962
rect 13858 12910 13860 12962
rect 12348 12798 12350 12850
rect 12402 12798 12404 12850
rect 12348 11618 12404 12798
rect 12908 12852 12964 12862
rect 12908 12758 12964 12796
rect 13692 12852 13748 12862
rect 13468 12740 13524 12750
rect 12348 11566 12350 11618
rect 12402 11566 12404 11618
rect 12236 11508 12292 11518
rect 12348 11508 12404 11566
rect 13020 12738 13524 12740
rect 13020 12686 13470 12738
rect 13522 12686 13524 12738
rect 13020 12684 13524 12686
rect 11788 11506 12068 11508
rect 11788 11454 11790 11506
rect 11842 11454 12068 11506
rect 11788 11452 12068 11454
rect 11788 11442 11844 11452
rect 11564 11218 11620 11228
rect 11004 10882 11060 10892
rect 10892 10724 10948 10734
rect 10892 10722 11060 10724
rect 10892 10670 10894 10722
rect 10946 10670 11060 10722
rect 10892 10668 11060 10670
rect 10892 10658 10948 10668
rect 10780 9174 10836 9212
rect 11004 9604 11060 10668
rect 11788 10722 11844 10734
rect 11788 10670 11790 10722
rect 11842 10670 11844 10722
rect 11228 10612 11284 10622
rect 11228 10518 11284 10556
rect 11564 10388 11620 10398
rect 11452 10386 11620 10388
rect 11452 10334 11566 10386
rect 11618 10334 11620 10386
rect 11452 10332 11620 10334
rect 11004 9042 11060 9548
rect 11004 8990 11006 9042
rect 11058 8990 11060 9042
rect 10444 8932 10500 8942
rect 10220 8818 10276 8830
rect 10220 8766 10222 8818
rect 10274 8766 10276 8818
rect 10220 8258 10276 8766
rect 10220 8206 10222 8258
rect 10274 8206 10276 8258
rect 10220 8194 10276 8206
rect 10108 6514 10164 6524
rect 8988 6020 9044 6030
rect 8988 6018 9156 6020
rect 8988 5966 8990 6018
rect 9042 5966 9156 6018
rect 8988 5964 9156 5966
rect 8988 5954 9044 5964
rect 8764 5122 8820 5134
rect 8764 5070 8766 5122
rect 8818 5070 8820 5122
rect 8764 4116 8820 5070
rect 8876 5012 8932 5740
rect 8988 5124 9044 5134
rect 8988 5030 9044 5068
rect 8876 4946 8932 4956
rect 8764 4050 8820 4060
rect 9100 3892 9156 5964
rect 10444 5908 10500 8876
rect 11004 8930 11060 8990
rect 11340 9940 11396 9950
rect 11340 9044 11396 9884
rect 11452 9268 11508 10332
rect 11564 10322 11620 10332
rect 11788 10052 11844 10670
rect 11900 10388 11956 10398
rect 11900 10294 11956 10332
rect 11900 10052 11956 10062
rect 11788 10050 11956 10052
rect 11788 9998 11902 10050
rect 11954 9998 11956 10050
rect 11788 9996 11956 9998
rect 11564 9940 11620 9950
rect 11564 9846 11620 9884
rect 11676 9604 11732 9614
rect 11564 9268 11620 9278
rect 11452 9266 11620 9268
rect 11452 9214 11566 9266
rect 11618 9214 11620 9266
rect 11452 9212 11620 9214
rect 11564 9202 11620 9212
rect 11676 9266 11732 9548
rect 11676 9214 11678 9266
rect 11730 9214 11732 9266
rect 11676 9202 11732 9214
rect 11452 9044 11508 9054
rect 11340 9042 11508 9044
rect 11340 8990 11454 9042
rect 11506 8990 11508 9042
rect 11340 8988 11508 8990
rect 11452 8978 11508 8988
rect 11004 8878 11006 8930
rect 11058 8878 11060 8930
rect 11004 8866 11060 8878
rect 11788 8820 11844 9996
rect 11900 9986 11956 9996
rect 12012 9380 12068 11452
rect 12236 11506 12404 11508
rect 12236 11454 12238 11506
rect 12290 11454 12404 11506
rect 12236 11452 12404 11454
rect 12236 11442 12292 11452
rect 12236 9826 12292 9838
rect 12236 9774 12238 9826
rect 12290 9774 12292 9826
rect 12236 9604 12292 9774
rect 12236 9538 12292 9548
rect 12012 9314 12068 9324
rect 12236 9268 12292 9278
rect 12348 9268 12404 11452
rect 12796 11508 12852 11518
rect 12572 11284 12628 11294
rect 12572 11190 12628 11228
rect 12796 10498 12852 11452
rect 12908 11396 12964 11406
rect 13020 11396 13076 12684
rect 13468 12674 13524 12684
rect 13692 12066 13748 12796
rect 13692 12014 13694 12066
rect 13746 12014 13748 12066
rect 13692 12002 13748 12014
rect 13804 11508 13860 12910
rect 14140 12628 14196 14588
rect 14700 14642 14756 15260
rect 15036 15314 15092 15484
rect 16156 15428 16212 15932
rect 17052 15874 17108 15886
rect 17052 15822 17054 15874
rect 17106 15822 17108 15874
rect 17052 15652 17108 15822
rect 16716 15596 17108 15652
rect 16716 15538 16772 15596
rect 16716 15486 16718 15538
rect 16770 15486 16772 15538
rect 16716 15474 16772 15486
rect 17276 15540 17332 15550
rect 16604 15428 16660 15438
rect 16156 15426 16660 15428
rect 16156 15374 16606 15426
rect 16658 15374 16660 15426
rect 16156 15372 16660 15374
rect 16604 15362 16660 15372
rect 15036 15262 15038 15314
rect 15090 15262 15092 15314
rect 15036 15250 15092 15262
rect 15484 15316 15540 15326
rect 15484 15314 15652 15316
rect 15484 15262 15486 15314
rect 15538 15262 15652 15314
rect 15484 15260 15652 15262
rect 15484 15250 15540 15260
rect 14700 14590 14702 14642
rect 14754 14590 14756 14642
rect 14700 14578 14756 14590
rect 14140 12562 14196 12572
rect 14364 12964 14420 12974
rect 14140 12068 14196 12078
rect 14140 11974 14196 12012
rect 13804 11442 13860 11452
rect 12908 11394 13076 11396
rect 12908 11342 12910 11394
rect 12962 11342 13076 11394
rect 12908 11340 13076 11342
rect 12908 11330 12964 11340
rect 13692 11284 13748 11294
rect 14364 11284 14420 12908
rect 15148 12852 15204 12862
rect 15148 12850 15540 12852
rect 15148 12798 15150 12850
rect 15202 12798 15540 12850
rect 15148 12796 15540 12798
rect 15148 12786 15204 12796
rect 14476 12180 14532 12190
rect 14476 12086 14532 12124
rect 14812 12178 14868 12190
rect 14812 12126 14814 12178
rect 14866 12126 14868 12178
rect 13692 11282 14420 11284
rect 13692 11230 13694 11282
rect 13746 11230 14420 11282
rect 13692 11228 14420 11230
rect 14588 12066 14644 12078
rect 14588 12014 14590 12066
rect 14642 12014 14644 12066
rect 12796 10446 12798 10498
rect 12850 10446 12852 10498
rect 12460 9940 12516 9950
rect 12460 9846 12516 9884
rect 12796 9828 12852 10446
rect 13020 10610 13076 10622
rect 13020 10558 13022 10610
rect 13074 10558 13076 10610
rect 13020 10500 13076 10558
rect 13020 10434 13076 10444
rect 13580 10612 13636 10622
rect 12908 9828 12964 9838
rect 12796 9772 12908 9828
rect 13580 9828 13636 10556
rect 13692 10500 13748 11228
rect 14588 11172 14644 12014
rect 13804 11116 14644 11172
rect 14700 12068 14756 12078
rect 13804 10722 13860 11116
rect 13804 10670 13806 10722
rect 13858 10670 13860 10722
rect 13804 10658 13860 10670
rect 14476 10948 14532 10958
rect 13692 10434 13748 10444
rect 13916 10612 13972 10622
rect 13692 9828 13748 9838
rect 13580 9826 13748 9828
rect 13580 9774 13694 9826
rect 13746 9774 13748 9826
rect 13580 9772 13748 9774
rect 12908 9734 12964 9772
rect 13692 9492 13748 9772
rect 13916 9604 13972 10556
rect 13692 9426 13748 9436
rect 13804 9602 13972 9604
rect 13804 9550 13918 9602
rect 13970 9550 13972 9602
rect 13804 9548 13972 9550
rect 12236 9266 12404 9268
rect 12236 9214 12238 9266
rect 12290 9214 12404 9266
rect 12236 9212 12404 9214
rect 12236 9202 12292 9212
rect 12908 9156 12964 9166
rect 12796 9154 12964 9156
rect 12796 9102 12910 9154
rect 12962 9102 12964 9154
rect 12796 9100 12964 9102
rect 12572 8930 12628 8942
rect 12572 8878 12574 8930
rect 12626 8878 12628 8930
rect 11340 8764 11844 8820
rect 11900 8820 11956 8830
rect 11340 8484 11396 8764
rect 10780 8428 11396 8484
rect 10780 8258 10836 8428
rect 11340 8370 11396 8428
rect 11340 8318 11342 8370
rect 11394 8318 11396 8370
rect 11340 8306 11396 8318
rect 11676 8372 11732 8382
rect 11676 8278 11732 8316
rect 10780 8206 10782 8258
rect 10834 8206 10836 8258
rect 10780 8194 10836 8206
rect 11116 8258 11172 8270
rect 11116 8206 11118 8258
rect 11170 8206 11172 8258
rect 10668 8148 10724 8158
rect 10668 8054 10724 8092
rect 10556 8034 10612 8046
rect 10556 7982 10558 8034
rect 10610 7982 10612 8034
rect 10556 7812 10612 7982
rect 11116 7812 11172 8206
rect 10556 7756 11172 7812
rect 10556 7362 10612 7374
rect 10556 7310 10558 7362
rect 10610 7310 10612 7362
rect 10556 6804 10612 7310
rect 10556 6738 10612 6748
rect 10892 7028 10948 7038
rect 10444 5842 10500 5852
rect 9996 5796 10052 5806
rect 9996 5124 10052 5740
rect 9772 5122 10052 5124
rect 9772 5070 9998 5122
rect 10050 5070 10052 5122
rect 9772 5068 10052 5070
rect 9436 4898 9492 4910
rect 9436 4846 9438 4898
rect 9490 4846 9492 4898
rect 9436 4004 9492 4846
rect 9436 3938 9492 3948
rect 9548 4898 9604 4910
rect 9548 4846 9550 4898
rect 9602 4846 9604 4898
rect 9100 3826 9156 3836
rect 8652 3714 8708 3724
rect 9548 3778 9604 4846
rect 9660 4900 9716 4910
rect 9660 4806 9716 4844
rect 9660 4340 9716 4350
rect 9772 4340 9828 5068
rect 9996 5058 10052 5068
rect 10780 5012 10836 5022
rect 10780 4918 10836 4956
rect 9660 4338 9828 4340
rect 9660 4286 9662 4338
rect 9714 4286 9828 4338
rect 9660 4284 9828 4286
rect 10444 4900 10500 4910
rect 9660 4274 9716 4284
rect 10332 4228 10388 4238
rect 9884 4226 10388 4228
rect 9884 4174 10334 4226
rect 10386 4174 10388 4226
rect 9884 4172 10388 4174
rect 9548 3726 9550 3778
rect 9602 3726 9604 3778
rect 9548 3714 9604 3726
rect 9772 3892 9828 3902
rect 8764 3556 8820 3566
rect 8204 3444 8260 3454
rect 6972 2706 7028 2716
rect 7420 3330 7476 3342
rect 7420 3278 7422 3330
rect 7474 3278 7476 3330
rect 7420 1762 7476 3278
rect 7868 3332 7924 3342
rect 8204 3332 8260 3388
rect 8316 3332 8372 3342
rect 8204 3330 8372 3332
rect 8204 3278 8318 3330
rect 8370 3278 8372 3330
rect 8204 3276 8372 3278
rect 7868 3238 7924 3276
rect 8316 3266 8372 3276
rect 8764 3330 8820 3500
rect 9772 3442 9828 3836
rect 9884 3778 9940 4172
rect 10332 4162 10388 4172
rect 9884 3726 9886 3778
rect 9938 3726 9940 3778
rect 9884 3714 9940 3726
rect 10220 4004 10276 4014
rect 10220 3666 10276 3948
rect 10444 3778 10500 4844
rect 10892 4676 10948 6972
rect 11116 6804 11172 7756
rect 11676 6804 11732 6814
rect 11116 6802 11732 6804
rect 11116 6750 11678 6802
rect 11730 6750 11732 6802
rect 11116 6748 11732 6750
rect 11676 6738 11732 6748
rect 11788 5012 11844 5022
rect 10892 4610 10948 4620
rect 11228 4900 11284 4910
rect 10444 3726 10446 3778
rect 10498 3726 10500 3778
rect 10444 3714 10500 3726
rect 10780 3780 10836 3790
rect 10780 3686 10836 3724
rect 10220 3614 10222 3666
rect 10274 3614 10276 3666
rect 10220 3602 10276 3614
rect 11228 3666 11284 4844
rect 11676 4564 11732 4574
rect 11340 4452 11396 4462
rect 11340 3778 11396 4396
rect 11340 3726 11342 3778
rect 11394 3726 11396 3778
rect 11340 3714 11396 3726
rect 11676 3892 11732 4508
rect 11228 3614 11230 3666
rect 11282 3614 11284 3666
rect 11228 3602 11284 3614
rect 11676 3554 11732 3836
rect 11788 3666 11844 4956
rect 11900 4116 11956 8764
rect 12572 8818 12628 8878
rect 12572 8766 12574 8818
rect 12626 8766 12628 8818
rect 12572 8754 12628 8766
rect 12124 8316 12404 8372
rect 12012 8258 12068 8270
rect 12012 8206 12014 8258
rect 12066 8206 12068 8258
rect 12012 7588 12068 8206
rect 12012 6802 12068 7532
rect 12012 6750 12014 6802
rect 12066 6750 12068 6802
rect 12012 6738 12068 6750
rect 12124 5796 12180 8316
rect 12348 8258 12404 8316
rect 12348 8206 12350 8258
rect 12402 8206 12404 8258
rect 12348 8194 12404 8206
rect 12684 8260 12740 8270
rect 12684 8166 12740 8204
rect 12236 8146 12292 8158
rect 12236 8094 12238 8146
rect 12290 8094 12292 8146
rect 12236 7588 12292 8094
rect 12796 7812 12852 9100
rect 12908 9090 12964 9100
rect 13692 9154 13748 9166
rect 13692 9102 13694 9154
rect 13746 9102 13748 9154
rect 13132 9044 13188 9054
rect 13580 9044 13636 9054
rect 13132 9042 13636 9044
rect 13132 8990 13134 9042
rect 13186 8990 13582 9042
rect 13634 8990 13636 9042
rect 13132 8988 13636 8990
rect 13132 8372 13188 8988
rect 13580 8978 13636 8988
rect 13132 8306 13188 8316
rect 13020 8148 13076 8158
rect 13020 8054 13076 8092
rect 13020 7924 13076 7934
rect 12796 7746 12852 7756
rect 12908 7868 13020 7924
rect 12236 7532 12852 7588
rect 12236 7364 12292 7374
rect 12236 6690 12292 7308
rect 12684 7364 12740 7402
rect 12684 7298 12740 7308
rect 12236 6638 12238 6690
rect 12290 6638 12292 6690
rect 12236 6626 12292 6638
rect 12348 7252 12404 7262
rect 12348 6690 12404 7196
rect 12348 6638 12350 6690
rect 12402 6638 12404 6690
rect 12348 6626 12404 6638
rect 12684 7140 12740 7150
rect 12684 6690 12740 7084
rect 12684 6638 12686 6690
rect 12738 6638 12740 6690
rect 12684 6626 12740 6638
rect 12124 5730 12180 5740
rect 12796 5236 12852 7532
rect 12908 6692 12964 7868
rect 13020 7858 13076 7868
rect 13692 7812 13748 9102
rect 13244 7756 13748 7812
rect 13020 7700 13076 7710
rect 13020 7140 13076 7644
rect 13244 7698 13300 7756
rect 13244 7646 13246 7698
rect 13298 7646 13300 7698
rect 13020 7074 13076 7084
rect 13132 7362 13188 7374
rect 13132 7310 13134 7362
rect 13186 7310 13188 7362
rect 13020 6692 13076 6702
rect 12908 6690 13076 6692
rect 12908 6638 13022 6690
rect 13074 6638 13076 6690
rect 12908 6636 13076 6638
rect 13020 6626 13076 6636
rect 13132 6692 13188 7310
rect 13244 7364 13300 7646
rect 13244 7298 13300 7308
rect 13468 7588 13524 7598
rect 13804 7588 13860 9548
rect 13916 9538 13972 9548
rect 14364 9268 14420 9278
rect 13916 9042 13972 9054
rect 13916 8990 13918 9042
rect 13970 8990 13972 9042
rect 13916 8370 13972 8990
rect 13916 8318 13918 8370
rect 13970 8318 13972 8370
rect 13916 8306 13972 8318
rect 13468 7586 13860 7588
rect 13468 7534 13470 7586
rect 13522 7534 13860 7586
rect 13468 7532 13860 7534
rect 14140 8258 14196 8270
rect 14140 8206 14142 8258
rect 14194 8206 14196 8258
rect 13132 6626 13188 6636
rect 13356 7140 13412 7150
rect 13356 6690 13412 7084
rect 13356 6638 13358 6690
rect 13410 6638 13412 6690
rect 13356 6626 13412 6638
rect 12908 5236 12964 5246
rect 12796 5234 13188 5236
rect 12796 5182 12910 5234
rect 12962 5182 13188 5234
rect 12796 5180 13188 5182
rect 12908 5170 12964 5180
rect 12908 4564 12964 4574
rect 12908 4470 12964 4508
rect 13132 4562 13188 5180
rect 13356 5124 13412 5134
rect 13132 4510 13134 4562
rect 13186 4510 13188 4562
rect 12460 4226 12516 4238
rect 12460 4174 12462 4226
rect 12514 4174 12516 4226
rect 11900 4050 11956 4060
rect 12124 4116 12180 4126
rect 11788 3614 11790 3666
rect 11842 3614 11844 3666
rect 11788 3602 11844 3614
rect 12012 3780 12068 3790
rect 11676 3502 11678 3554
rect 11730 3502 11732 3554
rect 11676 3490 11732 3502
rect 12012 3554 12068 3724
rect 12012 3502 12014 3554
rect 12066 3502 12068 3554
rect 12012 3490 12068 3502
rect 9772 3390 9774 3442
rect 9826 3390 9828 3442
rect 9772 3378 9828 3390
rect 11900 3444 11956 3454
rect 8764 3278 8766 3330
rect 8818 3278 8820 3330
rect 8764 3266 8820 3278
rect 10108 3332 10164 3342
rect 7420 1710 7422 1762
rect 7474 1710 7476 1762
rect 7420 1698 7476 1710
rect 8316 1762 8372 1774
rect 8316 1710 8318 1762
rect 8370 1710 8372 1762
rect 6524 1596 6692 1652
rect 6524 800 6580 1596
rect 8316 800 8372 1710
rect 10108 800 10164 3276
rect 11900 800 11956 3388
rect 12124 2996 12180 4060
rect 12460 4116 12516 4174
rect 12460 4050 12516 4060
rect 13020 4226 13076 4238
rect 13020 4174 13022 4226
rect 13074 4174 13076 4226
rect 13020 3892 13076 4174
rect 12236 3836 13076 3892
rect 12236 3554 12292 3836
rect 13132 3780 13188 4510
rect 12236 3502 12238 3554
rect 12290 3502 12292 3554
rect 12236 3490 12292 3502
rect 13020 3668 13076 3678
rect 13020 3388 13076 3612
rect 13132 3556 13188 3724
rect 13244 5068 13356 5124
rect 13244 3778 13300 5068
rect 13356 5058 13412 5068
rect 13468 4338 13524 7532
rect 13692 7364 13748 7374
rect 13580 6804 13636 6814
rect 13580 6690 13636 6748
rect 13580 6638 13582 6690
rect 13634 6638 13636 6690
rect 13580 6626 13636 6638
rect 13692 6690 13748 7308
rect 13916 7364 13972 7374
rect 14140 7364 14196 8206
rect 13916 7362 14196 7364
rect 13916 7310 13918 7362
rect 13970 7310 14196 7362
rect 13916 7308 14196 7310
rect 13916 7252 13972 7308
rect 13916 7186 13972 7196
rect 13692 6638 13694 6690
rect 13746 6638 13748 6690
rect 13692 6626 13748 6638
rect 13916 6692 13972 6702
rect 13916 6598 13972 6636
rect 14364 5906 14420 9212
rect 14476 9266 14532 10892
rect 14476 9214 14478 9266
rect 14530 9214 14532 9266
rect 14476 9156 14532 9214
rect 14476 9090 14532 9100
rect 14700 7476 14756 12012
rect 14812 10500 14868 12126
rect 15036 12178 15092 12190
rect 15036 12126 15038 12178
rect 15090 12126 15092 12178
rect 15036 10836 15092 12126
rect 15372 12178 15428 12190
rect 15372 12126 15374 12178
rect 15426 12126 15428 12178
rect 15036 10770 15092 10780
rect 15260 11172 15316 11182
rect 14812 10434 14868 10444
rect 15260 9938 15316 11116
rect 15372 10612 15428 12126
rect 15484 11956 15540 12796
rect 15596 12516 15652 15260
rect 15708 15314 15764 15326
rect 15708 15262 15710 15314
rect 15762 15262 15764 15314
rect 15708 13748 15764 15262
rect 16044 15316 16100 15326
rect 16828 15316 16884 15326
rect 16044 15314 16324 15316
rect 16044 15262 16046 15314
rect 16098 15262 16324 15314
rect 16044 15260 16324 15262
rect 16044 15250 16100 15260
rect 15820 15204 15876 15214
rect 15820 15110 15876 15148
rect 16044 13748 16100 13758
rect 15708 13692 16044 13748
rect 16044 13634 16100 13692
rect 16044 13582 16046 13634
rect 16098 13582 16100 13634
rect 15932 13524 15988 13534
rect 15596 12460 15876 12516
rect 15820 12402 15876 12460
rect 15820 12350 15822 12402
rect 15874 12350 15876 12402
rect 15820 12338 15876 12350
rect 15932 12402 15988 13468
rect 15932 12350 15934 12402
rect 15986 12350 15988 12402
rect 15932 12338 15988 12350
rect 15708 12180 15764 12190
rect 16044 12180 16100 13582
rect 16268 13524 16324 15260
rect 16828 14642 16884 15260
rect 16828 14590 16830 14642
rect 16882 14590 16884 14642
rect 16828 14578 16884 14590
rect 17276 14642 17332 15484
rect 17612 15538 17668 15932
rect 17612 15486 17614 15538
rect 17666 15486 17668 15538
rect 17612 15474 17668 15486
rect 17948 15204 18004 20132
rect 18060 19908 18116 19918
rect 18060 19906 18228 19908
rect 18060 19854 18062 19906
rect 18114 19854 18228 19906
rect 18060 19852 18228 19854
rect 18060 19842 18116 19852
rect 18060 18452 18116 18462
rect 18060 18358 18116 18396
rect 18172 18338 18228 19852
rect 18172 18286 18174 18338
rect 18226 18286 18228 18338
rect 18172 18274 18228 18286
rect 18172 17444 18228 17454
rect 18172 16884 18228 17388
rect 18172 16770 18228 16828
rect 18172 16718 18174 16770
rect 18226 16718 18228 16770
rect 18172 16706 18228 16718
rect 18284 15652 18340 24444
rect 18396 21476 18452 25452
rect 18620 24610 18676 26460
rect 18732 25506 18788 26572
rect 18732 25454 18734 25506
rect 18786 25454 18788 25506
rect 18732 25442 18788 25454
rect 19292 26178 19348 26572
rect 19292 26126 19294 26178
rect 19346 26126 19348 26178
rect 19292 25508 19348 26126
rect 19292 25442 19348 25452
rect 18620 24558 18622 24610
rect 18674 24558 18676 24610
rect 18620 24546 18676 24558
rect 19404 24722 19460 24734
rect 19404 24670 19406 24722
rect 19458 24670 19460 24722
rect 19404 23940 19460 24670
rect 19404 23874 19460 23884
rect 19516 23716 19572 30828
rect 19628 30818 19684 30828
rect 20076 30994 20132 31006
rect 20076 30942 20078 30994
rect 20130 30942 20132 30994
rect 20076 29988 20132 30942
rect 20076 29922 20132 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19852 29092 19908 29102
rect 19628 28644 19684 28654
rect 19628 28082 19684 28588
rect 19852 28642 19908 29036
rect 20188 28756 20244 31388
rect 20524 31332 20580 31612
rect 20636 31444 20692 36990
rect 20748 33570 20804 37102
rect 20972 35586 21028 35598
rect 20972 35534 20974 35586
rect 21026 35534 21028 35586
rect 20972 34916 21028 35534
rect 21308 35028 21364 38612
rect 21644 38164 21700 38782
rect 21756 38834 21812 38846
rect 21756 38782 21758 38834
rect 21810 38782 21812 38834
rect 21756 38274 21812 38782
rect 21756 38222 21758 38274
rect 21810 38222 21812 38274
rect 21756 38210 21812 38222
rect 21980 38834 22036 38846
rect 21980 38782 21982 38834
rect 22034 38782 22036 38834
rect 21644 38098 21700 38108
rect 21868 38052 21924 38062
rect 21868 37958 21924 37996
rect 21756 37828 21812 37838
rect 21756 37734 21812 37772
rect 21868 37266 21924 37278
rect 21868 37214 21870 37266
rect 21922 37214 21924 37266
rect 21868 37044 21924 37214
rect 21868 36978 21924 36988
rect 21980 36596 22036 38782
rect 22092 38722 22148 39004
rect 22652 38946 22708 39340
rect 22876 39060 22932 40236
rect 22988 39060 23044 39070
rect 22876 39058 23044 39060
rect 22876 39006 22990 39058
rect 23042 39006 23044 39058
rect 22876 39004 23044 39006
rect 24332 39060 24388 40572
rect 24444 40402 24500 40414
rect 24444 40350 24446 40402
rect 24498 40350 24500 40402
rect 24444 40292 24500 40350
rect 24444 40226 24500 40236
rect 24556 40178 24612 40190
rect 24556 40126 24558 40178
rect 24610 40126 24612 40178
rect 24556 39730 24612 40126
rect 24556 39678 24558 39730
rect 24610 39678 24612 39730
rect 24556 39666 24612 39678
rect 24668 39956 24724 39966
rect 24332 39004 24500 39060
rect 22988 38994 23044 39004
rect 22652 38894 22654 38946
rect 22706 38894 22708 38946
rect 22652 38882 22708 38894
rect 23772 38948 23828 38958
rect 23772 38854 23828 38892
rect 22092 38670 22094 38722
rect 22146 38670 22148 38722
rect 22092 38658 22148 38670
rect 22204 38834 22260 38846
rect 22204 38782 22206 38834
rect 22258 38782 22260 38834
rect 22204 38724 22260 38782
rect 23324 38836 23380 38846
rect 23324 38742 23380 38780
rect 23884 38836 23940 38846
rect 24332 38836 24388 38846
rect 23940 38834 24388 38836
rect 23940 38782 24334 38834
rect 24386 38782 24388 38834
rect 23940 38780 24388 38782
rect 23884 38742 23940 38780
rect 24332 38770 24388 38780
rect 24444 38836 24500 39004
rect 24668 39058 24724 39900
rect 24668 39006 24670 39058
rect 24722 39006 24724 39058
rect 24668 38994 24724 39006
rect 24444 38770 24500 38780
rect 22540 38724 22596 38734
rect 22204 38722 22596 38724
rect 22204 38670 22542 38722
rect 22594 38670 22596 38722
rect 22204 38668 22596 38670
rect 22204 38388 22260 38668
rect 22540 38658 22596 38668
rect 23996 38612 24052 38622
rect 23996 38518 24052 38556
rect 21980 36530 22036 36540
rect 22092 38332 22260 38388
rect 21868 36372 21924 36382
rect 22092 36372 22148 38332
rect 22764 38164 22820 38174
rect 22764 38070 22820 38108
rect 23324 38162 23380 38174
rect 23324 38110 23326 38162
rect 23378 38110 23380 38162
rect 22204 38050 22260 38062
rect 22204 37998 22206 38050
rect 22258 37998 22260 38050
rect 22204 37828 22260 37998
rect 22204 36708 22260 37772
rect 22428 38052 22484 38062
rect 22428 36932 22484 37996
rect 22540 37940 22596 37950
rect 22540 37266 22596 37884
rect 22540 37214 22542 37266
rect 22594 37214 22596 37266
rect 22540 37202 22596 37214
rect 22652 37826 22708 37838
rect 22652 37774 22654 37826
rect 22706 37774 22708 37826
rect 22540 36932 22596 36942
rect 22428 36876 22540 36932
rect 22540 36866 22596 36876
rect 22204 36642 22260 36652
rect 22316 36596 22372 36606
rect 22316 36482 22372 36540
rect 22316 36430 22318 36482
rect 22370 36430 22372 36482
rect 22316 36418 22372 36430
rect 21868 36370 22148 36372
rect 21868 36318 21870 36370
rect 21922 36318 22148 36370
rect 21868 36316 22148 36318
rect 21868 36306 21924 36316
rect 21644 36260 21700 36270
rect 21644 36166 21700 36204
rect 22652 36260 22708 37774
rect 22876 37828 22932 37838
rect 23324 37828 23380 38110
rect 22876 37826 23380 37828
rect 22876 37774 22878 37826
rect 22930 37774 23380 37826
rect 22876 37772 23380 37774
rect 22876 37762 22932 37772
rect 23100 37268 23156 37278
rect 23100 37174 23156 37212
rect 23324 37268 23380 37772
rect 24668 37940 24724 37950
rect 24668 37490 24724 37884
rect 24668 37438 24670 37490
rect 24722 37438 24724 37490
rect 24668 37426 24724 37438
rect 23324 37202 23380 37212
rect 23884 37268 23940 37278
rect 23324 36932 23380 36942
rect 22428 36036 22484 36046
rect 22428 35924 22484 35980
rect 22204 35922 22484 35924
rect 22204 35870 22430 35922
rect 22482 35870 22484 35922
rect 22204 35868 22484 35870
rect 22092 35812 22148 35822
rect 22092 35718 22148 35756
rect 21308 34962 21364 34972
rect 21420 35698 21476 35710
rect 21420 35646 21422 35698
rect 21474 35646 21476 35698
rect 20972 34850 21028 34860
rect 20860 34244 20916 34254
rect 20860 34130 20916 34188
rect 20860 34078 20862 34130
rect 20914 34078 20916 34130
rect 20860 34066 20916 34078
rect 20748 33518 20750 33570
rect 20802 33518 20804 33570
rect 20748 33506 20804 33518
rect 21420 33460 21476 35646
rect 21532 35698 21588 35710
rect 21532 35646 21534 35698
rect 21586 35646 21588 35698
rect 21532 35252 21588 35646
rect 21644 35700 21700 35710
rect 21644 35606 21700 35644
rect 21532 35186 21588 35196
rect 21644 35364 21700 35374
rect 20860 33404 21476 33460
rect 21532 34244 21588 34254
rect 20860 32786 20916 33404
rect 20860 32734 20862 32786
rect 20914 32734 20916 32786
rect 20860 32452 20916 32734
rect 20860 32386 20916 32396
rect 21196 32562 21252 32574
rect 21196 32510 21198 32562
rect 21250 32510 21252 32562
rect 21196 32004 21252 32510
rect 21532 32562 21588 34188
rect 21644 34242 21700 35308
rect 21644 34190 21646 34242
rect 21698 34190 21700 34242
rect 21644 34178 21700 34190
rect 22092 33460 22148 33470
rect 22204 33460 22260 35868
rect 22428 35858 22484 35868
rect 22652 35922 22708 36204
rect 22652 35870 22654 35922
rect 22706 35870 22708 35922
rect 22652 35858 22708 35870
rect 22876 36708 22932 36718
rect 22876 36482 22932 36652
rect 22876 36430 22878 36482
rect 22930 36430 22932 36482
rect 22876 35924 22932 36430
rect 23324 36482 23380 36876
rect 23324 36430 23326 36482
rect 23378 36430 23380 36482
rect 23324 36418 23380 36430
rect 23884 36370 23940 37212
rect 24556 37156 24612 37166
rect 24556 37062 24612 37100
rect 24668 36932 24724 36942
rect 24668 36594 24724 36876
rect 24668 36542 24670 36594
rect 24722 36542 24724 36594
rect 24668 36530 24724 36542
rect 23884 36318 23886 36370
rect 23938 36318 23940 36370
rect 23884 36306 23940 36318
rect 24108 36260 24164 36270
rect 24556 36260 24612 36270
rect 24164 36204 24388 36260
rect 24108 36166 24164 36204
rect 22876 35830 22932 35868
rect 23996 35924 24052 35934
rect 23996 35830 24052 35868
rect 23324 35810 23380 35822
rect 23324 35758 23326 35810
rect 23378 35758 23380 35810
rect 22540 35700 22596 35710
rect 22540 35606 22596 35644
rect 21532 32510 21534 32562
rect 21586 32510 21588 32562
rect 21532 32498 21588 32510
rect 21980 33458 22260 33460
rect 21980 33406 22094 33458
rect 22146 33406 22260 33458
rect 21980 33404 22260 33406
rect 22316 35476 22372 35486
rect 21196 31938 21252 31948
rect 21868 31780 21924 31790
rect 21868 31686 21924 31724
rect 20636 31378 20692 31388
rect 20748 31666 20804 31678
rect 20748 31614 20750 31666
rect 20802 31614 20804 31666
rect 20748 31556 20804 31614
rect 20524 31266 20580 31276
rect 20748 31218 20804 31500
rect 21532 31554 21588 31566
rect 21532 31502 21534 31554
rect 21586 31502 21588 31554
rect 21532 31444 21588 31502
rect 21532 31378 21588 31388
rect 20748 31166 20750 31218
rect 20802 31166 20804 31218
rect 20748 31154 20804 31166
rect 21532 31220 21588 31230
rect 20300 31108 20356 31118
rect 20300 31014 20356 31052
rect 21308 31108 21364 31118
rect 20636 30884 20692 30894
rect 20300 30882 20692 30884
rect 20300 30830 20638 30882
rect 20690 30830 20692 30882
rect 20300 30828 20692 30830
rect 20300 29314 20356 30828
rect 20636 30818 20692 30828
rect 20300 29262 20302 29314
rect 20354 29262 20356 29314
rect 20300 29250 20356 29262
rect 20636 30210 20692 30222
rect 20636 30158 20638 30210
rect 20690 30158 20692 30210
rect 20636 28980 20692 30158
rect 21196 29988 21252 29998
rect 20748 29428 20804 29438
rect 20748 29426 20916 29428
rect 20748 29374 20750 29426
rect 20802 29374 20916 29426
rect 20748 29372 20916 29374
rect 20748 29362 20804 29372
rect 20636 28924 20804 28980
rect 20188 28700 20356 28756
rect 19852 28590 19854 28642
rect 19906 28590 19908 28642
rect 19852 28420 19908 28590
rect 19852 28354 19908 28364
rect 20188 28530 20244 28542
rect 20188 28478 20190 28530
rect 20242 28478 20244 28530
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 28030 19630 28082
rect 19682 28030 19684 28082
rect 19628 28018 19684 28030
rect 19628 27860 19684 27870
rect 19628 26516 19684 27804
rect 19852 27860 19908 27870
rect 19852 27858 20020 27860
rect 19852 27806 19854 27858
rect 19906 27806 20020 27858
rect 19852 27804 20020 27806
rect 19852 27794 19908 27804
rect 19740 27746 19796 27758
rect 19740 27694 19742 27746
rect 19794 27694 19796 27746
rect 19740 27300 19796 27694
rect 19740 27234 19796 27244
rect 19852 27636 19908 27646
rect 19964 27636 20020 27804
rect 20076 27636 20132 27646
rect 20188 27636 20244 28478
rect 20300 27860 20356 28700
rect 20636 28644 20692 28682
rect 20636 28578 20692 28588
rect 20748 28084 20804 28924
rect 20748 27990 20804 28028
rect 20300 27794 20356 27804
rect 19964 27580 20076 27636
rect 20132 27580 20244 27636
rect 19852 27186 19908 27580
rect 20076 27570 20132 27580
rect 19852 27134 19854 27186
rect 19906 27134 19908 27186
rect 19852 27122 19908 27134
rect 20412 27188 20468 27198
rect 20412 26962 20468 27132
rect 20748 27188 20804 27198
rect 20748 27074 20804 27132
rect 20748 27022 20750 27074
rect 20802 27022 20804 27074
rect 20748 27010 20804 27022
rect 20412 26910 20414 26962
rect 20466 26910 20468 26962
rect 20412 26898 20468 26910
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19740 26516 19796 26526
rect 19628 26514 19796 26516
rect 19628 26462 19742 26514
rect 19794 26462 19796 26514
rect 19628 26460 19796 26462
rect 19740 26450 19796 26460
rect 20524 26516 20580 26526
rect 19628 25508 19684 25518
rect 19628 25414 19684 25452
rect 20412 25508 20468 25518
rect 20412 25414 20468 25452
rect 20524 25506 20580 26460
rect 20524 25454 20526 25506
rect 20578 25454 20580 25506
rect 20524 25442 20580 25454
rect 20748 25508 20804 25518
rect 20748 25414 20804 25452
rect 20076 25394 20132 25406
rect 20076 25342 20078 25394
rect 20130 25342 20132 25394
rect 19740 25284 19796 25294
rect 19628 25282 19796 25284
rect 19628 25230 19742 25282
rect 19794 25230 19796 25282
rect 19628 25228 19796 25230
rect 19628 24612 19684 25228
rect 19740 25218 19796 25228
rect 20076 25284 20132 25342
rect 20076 25218 20132 25228
rect 20300 25284 20356 25294
rect 20300 25190 20356 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20748 24722 20804 24734
rect 20748 24670 20750 24722
rect 20802 24670 20804 24722
rect 19628 24556 20020 24612
rect 19964 24050 20020 24556
rect 20748 24164 20804 24670
rect 20748 24098 20804 24108
rect 19964 23998 19966 24050
rect 20018 23998 20020 24050
rect 19964 23986 20020 23998
rect 20860 24052 20916 29372
rect 21084 28980 21140 28990
rect 21084 28532 21140 28924
rect 21196 28868 21252 29932
rect 21308 29540 21364 31052
rect 21420 30996 21476 31006
rect 21420 30902 21476 30940
rect 21420 29986 21476 29998
rect 21420 29934 21422 29986
rect 21474 29934 21476 29986
rect 21420 29764 21476 29934
rect 21420 29698 21476 29708
rect 21420 29540 21476 29550
rect 21308 29538 21476 29540
rect 21308 29486 21422 29538
rect 21474 29486 21476 29538
rect 21308 29484 21476 29486
rect 21420 29474 21476 29484
rect 21308 28868 21364 28878
rect 21196 28866 21364 28868
rect 21196 28814 21310 28866
rect 21362 28814 21364 28866
rect 21196 28812 21364 28814
rect 21308 28802 21364 28812
rect 21084 28082 21140 28476
rect 21084 28030 21086 28082
rect 21138 28030 21140 28082
rect 21084 28018 21140 28030
rect 21420 27858 21476 27870
rect 21420 27806 21422 27858
rect 21474 27806 21476 27858
rect 21308 27186 21364 27198
rect 21308 27134 21310 27186
rect 21362 27134 21364 27186
rect 21308 26908 21364 27134
rect 21420 27188 21476 27806
rect 21420 27122 21476 27132
rect 21196 26852 21364 26908
rect 21420 26964 21476 26974
rect 20972 26516 21028 26526
rect 20972 26422 21028 26460
rect 21196 25396 21252 26852
rect 21420 26514 21476 26908
rect 21420 26462 21422 26514
rect 21474 26462 21476 26514
rect 21420 26450 21476 26462
rect 21308 26180 21364 26190
rect 21308 26086 21364 26124
rect 21196 25330 21252 25340
rect 21308 25394 21364 25406
rect 21308 25342 21310 25394
rect 21362 25342 21364 25394
rect 21308 24948 21364 25342
rect 21532 25396 21588 31164
rect 21868 30212 21924 30222
rect 21980 30212 22036 33404
rect 22092 33394 22148 33404
rect 22316 33236 22372 35420
rect 23324 35364 23380 35758
rect 23548 35812 23604 35822
rect 23548 35698 23604 35756
rect 24108 35700 24164 35710
rect 23548 35646 23550 35698
rect 23602 35646 23604 35698
rect 23548 35634 23604 35646
rect 23884 35698 24164 35700
rect 23884 35646 24110 35698
rect 24162 35646 24164 35698
rect 23884 35644 24164 35646
rect 23324 35298 23380 35308
rect 23660 35252 23716 35262
rect 22988 34916 23044 34926
rect 22988 33796 23044 34860
rect 23548 34802 23604 34814
rect 23548 34750 23550 34802
rect 23602 34750 23604 34802
rect 23548 34244 23604 34750
rect 23548 34178 23604 34188
rect 22988 33740 23604 33796
rect 22092 33180 22372 33236
rect 23436 33572 23492 33582
rect 22092 31780 22148 33180
rect 22316 32452 22372 32462
rect 22316 32450 22596 32452
rect 22316 32398 22318 32450
rect 22370 32398 22596 32450
rect 22316 32396 22596 32398
rect 22316 32386 22372 32396
rect 22540 32002 22596 32396
rect 22540 31950 22542 32002
rect 22594 31950 22596 32002
rect 22540 31938 22596 31950
rect 22428 31780 22484 31790
rect 22988 31780 23044 31790
rect 22092 31778 22484 31780
rect 22092 31726 22430 31778
rect 22482 31726 22484 31778
rect 22092 31724 22484 31726
rect 22092 31666 22148 31724
rect 22428 31714 22484 31724
rect 22540 31778 23044 31780
rect 22540 31726 22990 31778
rect 23042 31726 23044 31778
rect 22540 31724 23044 31726
rect 22092 31614 22094 31666
rect 22146 31614 22148 31666
rect 22092 31602 22148 31614
rect 22540 31666 22596 31724
rect 22988 31714 23044 31724
rect 23436 31778 23492 33516
rect 23436 31726 23438 31778
rect 23490 31726 23492 31778
rect 23436 31714 23492 31726
rect 22540 31614 22542 31666
rect 22594 31614 22596 31666
rect 22540 31602 22596 31614
rect 22092 30884 22148 30894
rect 22764 30884 22820 30894
rect 22092 30882 22596 30884
rect 22092 30830 22094 30882
rect 22146 30830 22596 30882
rect 22092 30828 22596 30830
rect 22092 30818 22148 30828
rect 21868 30210 22036 30212
rect 21868 30158 21870 30210
rect 21922 30158 22036 30210
rect 21868 30156 22036 30158
rect 21868 30146 21924 30156
rect 21644 29986 21700 29998
rect 21644 29934 21646 29986
rect 21698 29934 21700 29986
rect 21644 29876 21700 29934
rect 21644 28644 21700 29820
rect 21644 28578 21700 28588
rect 21756 29986 21812 29998
rect 21756 29934 21758 29986
rect 21810 29934 21812 29986
rect 21756 28642 21812 29934
rect 22428 29988 22484 29998
rect 22428 29894 22484 29932
rect 22540 28866 22596 30828
rect 22652 30098 22708 30110
rect 22652 30046 22654 30098
rect 22706 30046 22708 30098
rect 22652 29876 22708 30046
rect 22652 29810 22708 29820
rect 22540 28814 22542 28866
rect 22594 28814 22596 28866
rect 22540 28802 22596 28814
rect 21756 28590 21758 28642
rect 21810 28590 21812 28642
rect 21756 28578 21812 28590
rect 21868 28756 21924 28766
rect 21868 28642 21924 28700
rect 21868 28590 21870 28642
rect 21922 28590 21924 28642
rect 21868 28578 21924 28590
rect 21980 28642 22036 28654
rect 21980 28590 21982 28642
rect 22034 28590 22036 28642
rect 21756 27972 21812 27982
rect 21756 27746 21812 27916
rect 21756 27694 21758 27746
rect 21810 27694 21812 27746
rect 21756 27682 21812 27694
rect 21980 27300 22036 28590
rect 22540 28644 22596 28654
rect 22428 28532 22484 28542
rect 22428 28438 22484 28476
rect 22540 28530 22596 28588
rect 22540 28478 22542 28530
rect 22594 28478 22596 28530
rect 22540 28466 22596 28478
rect 22764 28308 22820 30828
rect 23436 30436 23492 30446
rect 23212 30212 23268 30222
rect 22988 30100 23044 30110
rect 23212 30100 23268 30156
rect 22988 30098 23268 30100
rect 22988 30046 22990 30098
rect 23042 30046 23268 30098
rect 22988 30044 23268 30046
rect 22988 30034 23044 30044
rect 22764 28242 22820 28252
rect 22988 28868 23044 28878
rect 21980 27234 22036 27244
rect 22988 26852 23044 28812
rect 23100 28756 23156 28766
rect 23100 28662 23156 28700
rect 23212 28642 23268 30044
rect 23212 28590 23214 28642
rect 23266 28590 23268 28642
rect 23212 28578 23268 28590
rect 23324 30098 23380 30110
rect 23324 30046 23326 30098
rect 23378 30046 23380 30098
rect 23324 28644 23380 30046
rect 23324 28578 23380 28588
rect 23436 28420 23492 30380
rect 23548 30100 23604 33740
rect 23660 33458 23716 35196
rect 23660 33406 23662 33458
rect 23714 33406 23716 33458
rect 23660 33394 23716 33406
rect 23772 34020 23828 34030
rect 23884 34020 23940 35644
rect 24108 35634 24164 35644
rect 23772 34018 23940 34020
rect 23772 33966 23774 34018
rect 23826 33966 23940 34018
rect 23772 33964 23940 33966
rect 24332 34354 24388 36204
rect 24556 36036 24612 36204
rect 24556 35922 24612 35980
rect 24556 35870 24558 35922
rect 24610 35870 24612 35922
rect 24556 35858 24612 35870
rect 24332 34302 24334 34354
rect 24386 34302 24388 34354
rect 23772 33236 23828 33964
rect 24332 33572 24388 34302
rect 24444 34020 24500 34030
rect 24444 34018 24836 34020
rect 24444 33966 24446 34018
rect 24498 33966 24836 34018
rect 24444 33964 24836 33966
rect 24444 33954 24500 33964
rect 24332 33506 24388 33516
rect 24780 33346 24836 33964
rect 24780 33294 24782 33346
rect 24834 33294 24836 33346
rect 24668 33236 24724 33246
rect 23772 33234 24724 33236
rect 23772 33182 24670 33234
rect 24722 33182 24724 33234
rect 23772 33180 24724 33182
rect 24668 33170 24724 33180
rect 24780 33012 24836 33294
rect 24444 32956 24836 33012
rect 24444 32450 24500 32956
rect 24444 32398 24446 32450
rect 24498 32398 24500 32450
rect 24444 32386 24500 32398
rect 23884 32116 23940 32126
rect 23884 31890 23940 32060
rect 23884 31838 23886 31890
rect 23938 31838 23940 31890
rect 23884 31444 23940 31838
rect 23884 31378 23940 31388
rect 24556 31778 24612 31790
rect 24556 31726 24558 31778
rect 24610 31726 24612 31778
rect 24556 30996 24612 31726
rect 24220 30882 24276 30894
rect 24220 30830 24222 30882
rect 24274 30830 24276 30882
rect 24108 30322 24164 30334
rect 24108 30270 24110 30322
rect 24162 30270 24164 30322
rect 23548 30034 23604 30044
rect 23772 30210 23828 30222
rect 23772 30158 23774 30210
rect 23826 30158 23828 30210
rect 23772 29876 23828 30158
rect 24108 29988 24164 30270
rect 24220 30212 24276 30830
rect 24220 30146 24276 30156
rect 24220 29988 24276 29998
rect 24108 29932 24220 29988
rect 24220 29922 24276 29932
rect 23772 29810 23828 29820
rect 23884 29764 23940 29774
rect 23884 29650 23940 29708
rect 23884 29598 23886 29650
rect 23938 29598 23940 29650
rect 23884 29586 23940 29598
rect 23996 29428 24052 29438
rect 23548 29426 24052 29428
rect 23548 29374 23998 29426
rect 24050 29374 24052 29426
rect 23548 29372 24052 29374
rect 23548 29314 23604 29372
rect 23548 29262 23550 29314
rect 23602 29262 23604 29314
rect 23548 29250 23604 29262
rect 23996 28532 24052 29372
rect 24556 28756 24612 30940
rect 24668 30882 24724 30894
rect 24668 30830 24670 30882
rect 24722 30830 24724 30882
rect 24668 30100 24724 30830
rect 25004 30212 25060 46396
rect 27020 46114 27076 47292
rect 29708 47346 29764 47358
rect 29708 47294 29710 47346
rect 29762 47294 29764 47346
rect 29372 47236 29428 47246
rect 29372 47234 29652 47236
rect 29372 47182 29374 47234
rect 29426 47182 29652 47234
rect 29372 47180 29652 47182
rect 29372 47170 29428 47180
rect 29596 46786 29652 47180
rect 29596 46734 29598 46786
rect 29650 46734 29652 46786
rect 29596 46722 29652 46734
rect 28924 46674 28980 46686
rect 28924 46622 28926 46674
rect 28978 46622 28980 46674
rect 27020 46062 27022 46114
rect 27074 46062 27076 46114
rect 27020 46050 27076 46062
rect 28140 46562 28196 46574
rect 28140 46510 28142 46562
rect 28194 46510 28196 46562
rect 28140 46004 28196 46510
rect 28924 46004 28980 46622
rect 29708 46114 29764 47294
rect 31052 47346 31108 47358
rect 31052 47294 31054 47346
rect 31106 47294 31108 47346
rect 29708 46062 29710 46114
rect 29762 46062 29764 46114
rect 29708 46050 29764 46062
rect 30268 46228 30324 46238
rect 30268 46114 30324 46172
rect 30268 46062 30270 46114
rect 30322 46062 30324 46114
rect 30268 46050 30324 46062
rect 28140 45948 28420 46004
rect 26572 45892 26628 45902
rect 26572 45798 26628 45836
rect 27356 45892 27412 45902
rect 27356 45798 27412 45836
rect 27580 45892 27636 45902
rect 26684 45780 26740 45790
rect 26684 45686 26740 45724
rect 26460 45666 26516 45678
rect 26460 45614 26462 45666
rect 26514 45614 26516 45666
rect 26460 45332 26516 45614
rect 26460 45266 26516 45276
rect 26796 45332 26852 45342
rect 25228 45218 25284 45230
rect 25228 45166 25230 45218
rect 25282 45166 25284 45218
rect 25228 44436 25284 45166
rect 25564 45108 25620 45118
rect 25564 45014 25620 45052
rect 25228 44370 25284 44380
rect 26684 44436 26740 44446
rect 26684 44342 26740 44380
rect 25900 44100 25956 44110
rect 25900 43426 25956 44044
rect 26796 43708 26852 45276
rect 26908 45220 26964 45230
rect 26908 45106 26964 45164
rect 26908 45054 26910 45106
rect 26962 45054 26964 45106
rect 26908 45042 26964 45054
rect 27020 45108 27076 45118
rect 27020 44546 27076 45052
rect 27020 44494 27022 44546
rect 27074 44494 27076 44546
rect 27020 44482 27076 44494
rect 27132 45106 27188 45118
rect 27580 45108 27636 45836
rect 27916 45778 27972 45790
rect 27916 45726 27918 45778
rect 27970 45726 27972 45778
rect 27916 45220 27972 45726
rect 28028 45780 28084 45790
rect 28028 45686 28084 45724
rect 28252 45778 28308 45790
rect 28252 45726 28254 45778
rect 28306 45726 28308 45778
rect 28140 45332 28196 45342
rect 28140 45238 28196 45276
rect 27916 45154 27972 45164
rect 27132 45054 27134 45106
rect 27186 45054 27188 45106
rect 27132 44100 27188 45054
rect 27132 44034 27188 44044
rect 27244 45052 27636 45108
rect 27244 43708 27300 45052
rect 27804 44996 27860 45006
rect 27356 44994 27860 44996
rect 27356 44942 27806 44994
rect 27858 44942 27860 44994
rect 27356 44940 27860 44942
rect 27356 44546 27412 44940
rect 27804 44930 27860 44940
rect 27356 44494 27358 44546
rect 27410 44494 27412 44546
rect 27356 44482 27412 44494
rect 27916 44436 27972 44446
rect 27580 44322 27636 44334
rect 27580 44270 27582 44322
rect 27634 44270 27636 44322
rect 27580 43708 27636 44270
rect 27916 44324 27972 44380
rect 27916 44322 28196 44324
rect 27916 44270 27918 44322
rect 27970 44270 28196 44322
rect 27916 44268 28196 44270
rect 27916 44258 27972 44268
rect 26796 43652 27076 43708
rect 25900 43374 25902 43426
rect 25954 43374 25956 43426
rect 25900 43204 25956 43374
rect 26348 43426 26404 43438
rect 26348 43374 26350 43426
rect 26402 43374 26404 43426
rect 26236 43316 26292 43326
rect 25900 43138 25956 43148
rect 26012 43314 26292 43316
rect 26012 43262 26238 43314
rect 26290 43262 26292 43314
rect 26012 43260 26292 43262
rect 25452 42532 25508 42542
rect 25228 41972 25284 41982
rect 25228 41878 25284 41916
rect 25228 41188 25284 41198
rect 25228 39618 25284 41132
rect 25452 41076 25508 42476
rect 26012 42196 26068 43260
rect 26236 43250 26292 43260
rect 25564 42140 26068 42196
rect 25564 41298 25620 42140
rect 25564 41246 25566 41298
rect 25618 41246 25620 41298
rect 25564 41234 25620 41246
rect 25452 41020 25620 41076
rect 25452 40516 25508 40526
rect 25452 40422 25508 40460
rect 25228 39566 25230 39618
rect 25282 39566 25284 39618
rect 25228 39554 25284 39566
rect 25340 38836 25396 38846
rect 25340 38742 25396 38780
rect 25564 38500 25620 41020
rect 25900 40852 25956 40862
rect 25900 40626 25956 40796
rect 25900 40574 25902 40626
rect 25954 40574 25956 40626
rect 25900 40562 25956 40574
rect 26348 40628 26404 43374
rect 26908 43426 26964 43438
rect 26908 43374 26910 43426
rect 26962 43374 26964 43426
rect 26908 43092 26964 43374
rect 26796 43036 26964 43092
rect 26796 42756 26852 43036
rect 26908 42868 26964 42878
rect 26908 42774 26964 42812
rect 26796 42690 26852 42700
rect 26908 42532 26964 42542
rect 26908 40740 26964 42476
rect 26908 40674 26964 40684
rect 26348 40562 26404 40572
rect 25676 40402 25732 40414
rect 25676 40350 25678 40402
rect 25730 40350 25732 40402
rect 25676 39956 25732 40350
rect 26124 40402 26180 40414
rect 26124 40350 26126 40402
rect 26178 40350 26180 40402
rect 25788 40292 25844 40302
rect 25788 40198 25844 40236
rect 25676 39890 25732 39900
rect 25676 39730 25732 39742
rect 25676 39678 25678 39730
rect 25730 39678 25732 39730
rect 25676 39396 25732 39678
rect 25676 39330 25732 39340
rect 26124 39060 26180 40350
rect 26684 40290 26740 40302
rect 26684 40238 26686 40290
rect 26738 40238 26740 40290
rect 26572 39956 26628 39966
rect 26124 38994 26180 39004
rect 26236 39620 26292 39630
rect 25788 38948 25844 38958
rect 25788 38854 25844 38892
rect 25564 38434 25620 38444
rect 26236 38050 26292 39564
rect 26348 39396 26404 39406
rect 26348 38946 26404 39340
rect 26348 38894 26350 38946
rect 26402 38894 26404 38946
rect 26348 38882 26404 38894
rect 26572 39058 26628 39900
rect 26572 39006 26574 39058
rect 26626 39006 26628 39058
rect 26572 38668 26628 39006
rect 26684 39058 26740 40238
rect 26796 40180 26852 40190
rect 26796 40086 26852 40124
rect 26684 39006 26686 39058
rect 26738 39006 26740 39058
rect 26684 38994 26740 39006
rect 26908 39060 26964 39070
rect 26908 38966 26964 39004
rect 26796 38836 26852 38846
rect 26796 38742 26852 38780
rect 26236 37998 26238 38050
rect 26290 37998 26292 38050
rect 26236 37986 26292 37998
rect 26460 38612 26628 38668
rect 25452 37940 25508 37950
rect 25452 37846 25508 37884
rect 26460 37716 26516 38612
rect 25452 37660 26516 37716
rect 25452 37490 25508 37660
rect 25452 37438 25454 37490
rect 25506 37438 25508 37490
rect 25452 37426 25508 37438
rect 26348 37492 26404 37502
rect 25676 37380 25732 37390
rect 25676 37286 25732 37324
rect 25228 37268 25284 37278
rect 25228 37174 25284 37212
rect 25900 37268 25956 37278
rect 25900 37174 25956 37212
rect 26236 37266 26292 37278
rect 26236 37214 26238 37266
rect 26290 37214 26292 37266
rect 25564 37156 25620 37166
rect 25564 37062 25620 37100
rect 26236 36932 26292 37214
rect 26348 37044 26404 37436
rect 26460 37490 26516 37660
rect 26460 37438 26462 37490
rect 26514 37438 26516 37490
rect 26460 37426 26516 37438
rect 26572 37938 26628 37950
rect 26572 37886 26574 37938
rect 26626 37886 26628 37938
rect 26572 37490 26628 37886
rect 26572 37438 26574 37490
rect 26626 37438 26628 37490
rect 26572 37426 26628 37438
rect 26684 37826 26740 37838
rect 26684 37774 26686 37826
rect 26738 37774 26740 37826
rect 26684 37492 26740 37774
rect 26684 37436 26964 37492
rect 26684 37268 26740 37278
rect 26572 37266 26740 37268
rect 26572 37214 26686 37266
rect 26738 37214 26740 37266
rect 26572 37212 26740 37214
rect 26572 37044 26628 37212
rect 26348 36988 26628 37044
rect 26236 36866 26292 36876
rect 26684 36372 26740 37212
rect 26796 37268 26852 37278
rect 26796 37174 26852 37212
rect 26908 37044 26964 37436
rect 26796 36988 26964 37044
rect 26796 36594 26852 36988
rect 26796 36542 26798 36594
rect 26850 36542 26852 36594
rect 26796 36530 26852 36542
rect 27020 36596 27076 43652
rect 27132 43652 27636 43708
rect 27916 44100 27972 44110
rect 27132 39508 27188 43652
rect 27244 43538 27300 43550
rect 27244 43486 27246 43538
rect 27298 43486 27300 43538
rect 27244 42868 27300 43486
rect 27468 43538 27524 43550
rect 27468 43486 27470 43538
rect 27522 43486 27524 43538
rect 27356 43316 27412 43326
rect 27356 42978 27412 43260
rect 27356 42926 27358 42978
rect 27410 42926 27412 42978
rect 27356 42914 27412 42926
rect 27244 42802 27300 42812
rect 27244 42642 27300 42654
rect 27244 42590 27246 42642
rect 27298 42590 27300 42642
rect 27244 42084 27300 42590
rect 27468 42196 27524 43486
rect 27692 43538 27748 43550
rect 27692 43486 27694 43538
rect 27746 43486 27748 43538
rect 27580 43428 27636 43438
rect 27580 43334 27636 43372
rect 27692 43204 27748 43486
rect 27804 43540 27860 43550
rect 27804 43446 27860 43484
rect 27916 43316 27972 44044
rect 28140 43652 28196 44268
rect 28252 44100 28308 45726
rect 28364 45780 28420 45948
rect 28476 45780 28532 45790
rect 28364 45778 28532 45780
rect 28364 45726 28478 45778
rect 28530 45726 28532 45778
rect 28364 45724 28532 45726
rect 28476 45332 28532 45724
rect 28476 45276 28868 45332
rect 28588 45108 28644 45118
rect 28588 45014 28644 45052
rect 28700 45106 28756 45118
rect 28700 45054 28702 45106
rect 28754 45054 28756 45106
rect 28700 44100 28756 45054
rect 28812 45106 28868 45276
rect 28812 45054 28814 45106
rect 28866 45054 28868 45106
rect 28812 44212 28868 45054
rect 28924 44324 28980 45948
rect 29148 45892 29204 45902
rect 29148 45798 29204 45836
rect 29372 45892 29428 45902
rect 30604 45892 30660 45902
rect 29372 45890 30100 45892
rect 29372 45838 29374 45890
rect 29426 45838 30100 45890
rect 29372 45836 30100 45838
rect 29372 45826 29428 45836
rect 30044 45330 30100 45836
rect 30604 45798 30660 45836
rect 30828 45890 30884 45902
rect 30828 45838 30830 45890
rect 30882 45838 30884 45890
rect 30716 45332 30772 45342
rect 30044 45278 30046 45330
rect 30098 45278 30100 45330
rect 30044 45266 30100 45278
rect 30268 45330 30772 45332
rect 30268 45278 30718 45330
rect 30770 45278 30772 45330
rect 30268 45276 30772 45278
rect 29932 45220 29988 45230
rect 29932 45126 29988 45164
rect 30268 45106 30324 45276
rect 30716 45266 30772 45276
rect 30268 45054 30270 45106
rect 30322 45054 30324 45106
rect 30268 45042 30324 45054
rect 30604 45106 30660 45118
rect 30604 45054 30606 45106
rect 30658 45054 30660 45106
rect 30604 44996 30660 45054
rect 30604 44930 30660 44940
rect 30828 44548 30884 45838
rect 30940 45108 30996 45118
rect 30940 45014 30996 45052
rect 29148 44324 29204 44334
rect 28924 44322 29204 44324
rect 28924 44270 29150 44322
rect 29202 44270 29204 44322
rect 28924 44268 29204 44270
rect 29148 44258 29204 44268
rect 28812 44156 28980 44212
rect 28308 44044 28756 44100
rect 28252 44006 28308 44044
rect 28252 43652 28308 43662
rect 28140 43650 28308 43652
rect 28140 43598 28254 43650
rect 28306 43598 28308 43650
rect 28140 43596 28308 43598
rect 28252 43586 28308 43596
rect 27692 42308 27748 43148
rect 27804 43260 27972 43316
rect 28028 43540 28084 43550
rect 27804 42754 27860 43260
rect 27804 42702 27806 42754
rect 27858 42702 27860 42754
rect 27804 42690 27860 42702
rect 27916 42980 27972 42990
rect 27916 42754 27972 42924
rect 27916 42702 27918 42754
rect 27970 42702 27972 42754
rect 27916 42690 27972 42702
rect 27916 42308 27972 42318
rect 27692 42252 27916 42308
rect 27916 42242 27972 42252
rect 27468 42140 27860 42196
rect 27804 42084 27860 42140
rect 27916 42084 27972 42094
rect 27244 42028 27748 42084
rect 27244 41860 27300 41870
rect 27244 41766 27300 41804
rect 27356 40402 27412 42028
rect 27692 41298 27748 42028
rect 27692 41246 27694 41298
rect 27746 41246 27748 41298
rect 27692 41234 27748 41246
rect 27804 42028 27916 42084
rect 27804 41076 27860 42028
rect 27916 42018 27972 42028
rect 27468 41020 27860 41076
rect 27468 40626 27524 41020
rect 27692 40740 27748 40750
rect 27468 40574 27470 40626
rect 27522 40574 27524 40626
rect 27468 40562 27524 40574
rect 27580 40628 27636 40638
rect 27580 40534 27636 40572
rect 27692 40626 27748 40684
rect 27692 40574 27694 40626
rect 27746 40574 27748 40626
rect 27692 40562 27748 40574
rect 27356 40350 27358 40402
rect 27410 40350 27412 40402
rect 27356 40338 27412 40350
rect 27916 40404 27972 40414
rect 28028 40404 28084 43484
rect 28140 43428 28196 43438
rect 28924 43428 28980 44156
rect 29932 44210 29988 44222
rect 29932 44158 29934 44210
rect 29986 44158 29988 44210
rect 29932 43764 29988 44158
rect 30044 43764 30100 43774
rect 29932 43762 30100 43764
rect 29932 43710 30046 43762
rect 30098 43710 30100 43762
rect 29932 43708 30100 43710
rect 30044 43698 30100 43708
rect 30828 43652 30884 44492
rect 30716 43596 30884 43652
rect 29932 43540 29988 43550
rect 29148 43428 29204 43438
rect 28924 43372 29148 43428
rect 28140 42754 28196 43372
rect 29148 43334 29204 43372
rect 28364 43316 28420 43326
rect 28252 43092 28308 43102
rect 28252 42866 28308 43036
rect 28252 42814 28254 42866
rect 28306 42814 28308 42866
rect 28252 42802 28308 42814
rect 28140 42702 28142 42754
rect 28194 42702 28196 42754
rect 28140 42690 28196 42702
rect 28364 42754 28420 43260
rect 28476 43314 28532 43326
rect 28812 43316 28868 43326
rect 28476 43262 28478 43314
rect 28530 43262 28532 43314
rect 28476 42980 28532 43262
rect 28476 42914 28532 42924
rect 28588 43314 28868 43316
rect 28588 43262 28814 43314
rect 28866 43262 28868 43314
rect 28588 43260 28868 43262
rect 28364 42702 28366 42754
rect 28418 42702 28420 42754
rect 28364 42690 28420 42702
rect 28476 41300 28532 41310
rect 28588 41300 28644 43260
rect 28812 43250 28868 43260
rect 29372 43316 29428 43326
rect 29708 43316 29764 43326
rect 29372 43222 29428 43260
rect 29484 43314 29764 43316
rect 29484 43262 29710 43314
rect 29762 43262 29764 43314
rect 29484 43260 29764 43262
rect 28924 43204 28980 43214
rect 28924 41524 28980 43148
rect 28476 41298 28588 41300
rect 28476 41246 28478 41298
rect 28530 41246 28588 41298
rect 28476 41244 28588 41246
rect 28476 41234 28532 41244
rect 28588 41206 28644 41244
rect 28700 41468 28980 41524
rect 29036 43092 29092 43102
rect 28588 41076 28644 41086
rect 28700 41076 28756 41468
rect 29036 41188 29092 43036
rect 29148 42980 29204 42990
rect 29148 42886 29204 42924
rect 29260 42868 29316 42878
rect 29260 42774 29316 42812
rect 29484 41972 29540 43260
rect 29708 43250 29764 43260
rect 29932 42754 29988 43484
rect 30156 43426 30212 43438
rect 30156 43374 30158 43426
rect 30210 43374 30212 43426
rect 30156 42866 30212 43374
rect 30380 43316 30436 43326
rect 30156 42814 30158 42866
rect 30210 42814 30212 42866
rect 30156 42802 30212 42814
rect 30268 43260 30380 43316
rect 29932 42702 29934 42754
rect 29986 42702 29988 42754
rect 29932 42690 29988 42702
rect 29372 41300 29428 41310
rect 29148 41188 29204 41198
rect 29036 41186 29204 41188
rect 29036 41134 29150 41186
rect 29202 41134 29204 41186
rect 29036 41132 29204 41134
rect 29148 41122 29204 41132
rect 29372 41186 29428 41244
rect 29372 41134 29374 41186
rect 29426 41134 29428 41186
rect 29372 41122 29428 41134
rect 29484 41186 29540 41916
rect 30156 42644 30212 42654
rect 30268 42644 30324 43260
rect 30380 43250 30436 43260
rect 30604 42756 30660 42766
rect 30604 42662 30660 42700
rect 30156 42642 30324 42644
rect 30156 42590 30158 42642
rect 30210 42590 30324 42642
rect 30156 42588 30324 42590
rect 30156 41748 30212 42588
rect 30380 42532 30436 42542
rect 30380 42530 30548 42532
rect 30380 42478 30382 42530
rect 30434 42478 30548 42530
rect 30380 42476 30548 42478
rect 30380 42466 30436 42476
rect 30156 41682 30212 41692
rect 30492 42084 30548 42476
rect 29484 41134 29486 41186
rect 29538 41134 29540 41186
rect 29484 41122 29540 41134
rect 30380 41298 30436 41310
rect 30380 41246 30382 41298
rect 30434 41246 30436 41298
rect 28588 41074 28756 41076
rect 28588 41022 28590 41074
rect 28642 41022 28756 41074
rect 28588 41020 28756 41022
rect 28588 41010 28644 41020
rect 28140 40962 28196 40974
rect 29932 40964 29988 40974
rect 28140 40910 28142 40962
rect 28194 40910 28196 40962
rect 28140 40740 28196 40910
rect 28140 40674 28196 40684
rect 29820 40962 29988 40964
rect 29820 40910 29934 40962
rect 29986 40910 29988 40962
rect 29820 40908 29988 40910
rect 29820 40514 29876 40908
rect 29932 40898 29988 40908
rect 29820 40462 29822 40514
rect 29874 40462 29876 40514
rect 29820 40450 29876 40462
rect 30156 40516 30212 40526
rect 27916 40402 28420 40404
rect 27916 40350 27918 40402
rect 27970 40350 28420 40402
rect 27916 40348 28420 40350
rect 27916 40338 27972 40348
rect 27804 40180 27860 40190
rect 27804 39730 27860 40124
rect 27804 39678 27806 39730
rect 27858 39678 27860 39730
rect 27804 39666 27860 39678
rect 27132 39452 27860 39508
rect 27356 39060 27412 39070
rect 27132 38612 27188 38622
rect 27132 38162 27188 38556
rect 27132 38110 27134 38162
rect 27186 38110 27188 38162
rect 27132 37492 27188 38110
rect 27132 37426 27188 37436
rect 27356 37268 27412 39004
rect 27692 38834 27748 38846
rect 27692 38782 27694 38834
rect 27746 38782 27748 38834
rect 27692 38724 27748 38782
rect 27692 37828 27748 38668
rect 27692 37762 27748 37772
rect 27804 37492 27860 39452
rect 28364 39060 28420 40348
rect 30156 40402 30212 40460
rect 30156 40350 30158 40402
rect 30210 40350 30212 40402
rect 30156 40338 30212 40350
rect 28476 40290 28532 40302
rect 28476 40238 28478 40290
rect 28530 40238 28532 40290
rect 28476 39396 28532 40238
rect 28588 40180 28644 40190
rect 28588 40178 28980 40180
rect 28588 40126 28590 40178
rect 28642 40126 28980 40178
rect 28588 40124 28980 40126
rect 28588 40114 28644 40124
rect 28924 39732 28980 40124
rect 28924 39676 29988 39732
rect 28588 39618 28644 39630
rect 28588 39566 28590 39618
rect 28642 39566 28644 39618
rect 28588 39508 28644 39566
rect 28588 39442 28644 39452
rect 29372 39508 29428 39518
rect 28476 39330 28532 39340
rect 28476 39060 28532 39070
rect 28364 39058 28532 39060
rect 28364 39006 28478 39058
rect 28530 39006 28532 39058
rect 28364 39004 28532 39006
rect 28140 38836 28196 38846
rect 28140 38742 28196 38780
rect 28476 38052 28532 39004
rect 28700 38834 28756 38846
rect 28700 38782 28702 38834
rect 28754 38782 28756 38834
rect 28700 38668 28756 38782
rect 29260 38836 29316 38846
rect 29372 38836 29428 39452
rect 29260 38834 29428 38836
rect 29260 38782 29262 38834
rect 29314 38782 29428 38834
rect 29260 38780 29428 38782
rect 29484 39396 29540 39406
rect 29260 38770 29316 38780
rect 28588 38612 28756 38668
rect 28588 38164 28644 38612
rect 28588 38070 28644 38108
rect 28812 38276 28868 38286
rect 28476 37986 28532 37996
rect 28252 37940 28308 37950
rect 27916 37828 27972 37838
rect 27916 37734 27972 37772
rect 28252 37492 28308 37884
rect 27804 37490 28084 37492
rect 27804 37438 27806 37490
rect 27858 37438 28084 37490
rect 27804 37436 28084 37438
rect 27804 37426 27860 37436
rect 27356 37202 27412 37212
rect 27468 37266 27524 37278
rect 27468 37214 27470 37266
rect 27522 37214 27524 37266
rect 27020 36540 27412 36596
rect 26684 36316 26964 36372
rect 26796 35588 26852 35598
rect 26460 35586 26852 35588
rect 26460 35534 26798 35586
rect 26850 35534 26852 35586
rect 26460 35532 26852 35534
rect 25228 34244 25284 34254
rect 25228 34130 25284 34188
rect 25228 34078 25230 34130
rect 25282 34078 25284 34130
rect 25228 34066 25284 34078
rect 26012 34020 26068 34030
rect 25788 34018 26068 34020
rect 25788 33966 26014 34018
rect 26066 33966 26068 34018
rect 25788 33964 26068 33966
rect 25676 33124 25732 33134
rect 25676 32788 25732 33068
rect 25564 32732 25732 32788
rect 25788 32786 25844 33964
rect 26012 33954 26068 33964
rect 26460 33348 26516 35532
rect 26796 35522 26852 35532
rect 26908 33348 26964 36316
rect 27356 35812 27412 36540
rect 27356 35698 27412 35756
rect 27356 35646 27358 35698
rect 27410 35646 27412 35698
rect 27356 35634 27412 35646
rect 27020 35476 27076 35486
rect 27020 35474 27300 35476
rect 27020 35422 27022 35474
rect 27074 35422 27300 35474
rect 27020 35420 27300 35422
rect 27020 35410 27076 35420
rect 27244 35252 27300 35420
rect 27468 35364 27524 37214
rect 27580 37044 27636 37054
rect 27580 36482 27636 36988
rect 28028 36594 28084 37436
rect 28252 37398 28308 37436
rect 28812 37490 28868 38220
rect 29484 38162 29540 39340
rect 29820 38948 29876 38958
rect 29484 38110 29486 38162
rect 29538 38110 29540 38162
rect 29484 38098 29540 38110
rect 29596 38276 29652 38286
rect 29372 38052 29428 38062
rect 29372 37958 29428 37996
rect 29596 38050 29652 38220
rect 29596 37998 29598 38050
rect 29650 37998 29652 38050
rect 29596 37986 29652 37998
rect 29820 38052 29876 38892
rect 29932 38946 29988 39676
rect 29932 38894 29934 38946
rect 29986 38894 29988 38946
rect 29932 38882 29988 38894
rect 30044 39060 30100 39070
rect 29820 37996 29988 38052
rect 28812 37438 28814 37490
rect 28866 37438 28868 37490
rect 28812 37426 28868 37438
rect 29372 37828 29428 37838
rect 29148 37268 29204 37278
rect 28924 37266 29204 37268
rect 28924 37214 29150 37266
rect 29202 37214 29204 37266
rect 28924 37212 29204 37214
rect 28924 36820 28980 37212
rect 29148 37202 29204 37212
rect 28588 36764 28980 36820
rect 28588 36706 28644 36764
rect 28588 36654 28590 36706
rect 28642 36654 28644 36706
rect 28588 36642 28644 36654
rect 28028 36542 28030 36594
rect 28082 36542 28084 36594
rect 28028 36530 28084 36542
rect 29148 36594 29204 36606
rect 29148 36542 29150 36594
rect 29202 36542 29204 36594
rect 28252 36484 28308 36494
rect 27580 36430 27582 36482
rect 27634 36430 27636 36482
rect 27580 36418 27636 36430
rect 28140 36482 28308 36484
rect 28140 36430 28254 36482
rect 28306 36430 28308 36482
rect 28140 36428 28308 36430
rect 28140 36036 28196 36428
rect 28252 36418 28308 36428
rect 27916 35980 28196 36036
rect 27916 35810 27972 35980
rect 27916 35758 27918 35810
rect 27970 35758 27972 35810
rect 27916 35746 27972 35758
rect 28028 35812 28084 35822
rect 27580 35700 27636 35710
rect 27580 35606 27636 35644
rect 28028 35698 28084 35756
rect 28028 35646 28030 35698
rect 28082 35646 28084 35698
rect 28028 35634 28084 35646
rect 28588 35700 28644 35710
rect 28588 35606 28644 35644
rect 29148 35700 29204 36542
rect 29372 35812 29428 37772
rect 29820 37826 29876 37838
rect 29820 37774 29822 37826
rect 29874 37774 29876 37826
rect 29820 37492 29876 37774
rect 29820 37426 29876 37436
rect 29932 37490 29988 37996
rect 30044 38050 30100 39004
rect 30044 37998 30046 38050
rect 30098 37998 30100 38050
rect 30044 37986 30100 37998
rect 30156 38052 30212 38062
rect 29932 37438 29934 37490
rect 29986 37438 29988 37490
rect 29484 37378 29540 37390
rect 29484 37326 29486 37378
rect 29538 37326 29540 37378
rect 29484 36596 29540 37326
rect 29932 37156 29988 37438
rect 29932 37090 29988 37100
rect 30156 37268 30212 37996
rect 30380 37380 30436 41246
rect 30492 37828 30548 42028
rect 30716 42084 30772 43596
rect 30828 43426 30884 43438
rect 30828 43374 30830 43426
rect 30882 43374 30884 43426
rect 30828 43316 30884 43374
rect 30828 43250 30884 43260
rect 31052 42980 31108 47294
rect 32060 46674 32116 46686
rect 32060 46622 32062 46674
rect 32114 46622 32116 46674
rect 31724 46562 31780 46574
rect 31724 46510 31726 46562
rect 31778 46510 31780 46562
rect 31276 45892 31332 45902
rect 31332 45836 31556 45892
rect 31276 45826 31332 45836
rect 31500 45218 31556 45836
rect 31500 45166 31502 45218
rect 31554 45166 31556 45218
rect 31500 45154 31556 45166
rect 31164 45108 31220 45118
rect 31164 45106 31332 45108
rect 31164 45054 31166 45106
rect 31218 45054 31332 45106
rect 31164 45052 31332 45054
rect 31164 45042 31220 45052
rect 31276 44884 31332 45052
rect 31164 43538 31220 43550
rect 31164 43486 31166 43538
rect 31218 43486 31220 43538
rect 31164 43092 31220 43486
rect 31164 43026 31220 43036
rect 30716 42018 30772 42028
rect 30940 42924 31108 42980
rect 30828 41970 30884 41982
rect 30828 41918 30830 41970
rect 30882 41918 30884 41970
rect 30716 41412 30772 41422
rect 30604 41410 30772 41412
rect 30604 41358 30718 41410
rect 30770 41358 30772 41410
rect 30604 41356 30772 41358
rect 30604 38612 30660 41356
rect 30716 41346 30772 41356
rect 30828 41076 30884 41918
rect 30828 39508 30884 41020
rect 30828 39442 30884 39452
rect 30940 38668 30996 42924
rect 31276 42868 31332 44828
rect 31724 44884 31780 46510
rect 32060 46228 32116 46622
rect 32060 46162 32116 46172
rect 32172 46676 32228 47406
rect 32956 47348 33012 47358
rect 32396 47346 33012 47348
rect 32396 47294 32958 47346
rect 33010 47294 33012 47346
rect 32396 47292 33012 47294
rect 32396 46898 32452 47292
rect 32956 47282 33012 47292
rect 32396 46846 32398 46898
rect 32450 46846 32452 46898
rect 32396 46834 32452 46846
rect 33740 46898 33796 47964
rect 33740 46846 33742 46898
rect 33794 46846 33796 46898
rect 33740 46834 33796 46846
rect 34076 48018 34132 48030
rect 34076 47966 34078 48018
rect 34130 47966 34132 48018
rect 31948 46004 32004 46014
rect 32172 46004 32228 46620
rect 32004 45948 32228 46004
rect 31948 45910 32004 45948
rect 32956 45220 33012 45230
rect 32956 45126 33012 45164
rect 33404 45220 33460 45230
rect 31724 44818 31780 44828
rect 32172 45108 32228 45118
rect 32060 44436 32116 44446
rect 31948 44434 32116 44436
rect 31948 44382 32062 44434
rect 32114 44382 32116 44434
rect 31948 44380 32116 44382
rect 32172 44436 32228 45052
rect 33404 45106 33460 45164
rect 33404 45054 33406 45106
rect 33458 45054 33460 45106
rect 33404 45042 33460 45054
rect 33628 45108 33684 45118
rect 32396 44996 32452 45006
rect 32396 44902 32452 44940
rect 32508 44436 32564 44446
rect 33404 44436 33460 44446
rect 32172 44380 32508 44436
rect 31612 43540 31668 43550
rect 31612 43446 31668 43484
rect 31836 43538 31892 43550
rect 31836 43486 31838 43538
rect 31890 43486 31892 43538
rect 31052 42812 31332 42868
rect 31724 43426 31780 43438
rect 31724 43374 31726 43426
rect 31778 43374 31780 43426
rect 31052 42644 31108 42812
rect 31724 42756 31780 43374
rect 31836 43204 31892 43486
rect 31836 43138 31892 43148
rect 31948 43428 32004 44380
rect 32060 44370 32116 44380
rect 32508 44342 32564 44380
rect 32844 44434 33460 44436
rect 32844 44382 33406 44434
rect 33458 44382 33460 44434
rect 32844 44380 33460 44382
rect 32396 44100 32452 44110
rect 31052 42550 31108 42588
rect 31500 42700 31780 42756
rect 31948 42756 32004 43372
rect 31164 42530 31220 42542
rect 31164 42478 31166 42530
rect 31218 42478 31220 42530
rect 31164 42196 31220 42478
rect 31052 40404 31108 40414
rect 31164 40404 31220 42140
rect 31052 40402 31220 40404
rect 31052 40350 31054 40402
rect 31106 40350 31220 40402
rect 31052 40348 31220 40350
rect 31276 42084 31332 42094
rect 31052 40338 31108 40348
rect 31276 38668 31332 42028
rect 31500 42082 31556 42700
rect 31948 42662 32004 42700
rect 32060 44098 32452 44100
rect 32060 44046 32398 44098
rect 32450 44046 32452 44098
rect 32060 44044 32452 44046
rect 32060 42754 32116 44044
rect 32396 44034 32452 44044
rect 32620 43540 32676 43550
rect 32676 43484 32788 43540
rect 32620 43474 32676 43484
rect 32060 42702 32062 42754
rect 32114 42702 32116 42754
rect 32060 42690 32116 42702
rect 32172 43426 32228 43438
rect 32172 43374 32174 43426
rect 32226 43374 32228 43426
rect 31612 42532 31668 42542
rect 31612 42438 31668 42476
rect 31724 42530 31780 42542
rect 31724 42478 31726 42530
rect 31778 42478 31780 42530
rect 31612 42196 31668 42206
rect 31724 42196 31780 42478
rect 31668 42140 31780 42196
rect 31836 42530 31892 42542
rect 31836 42478 31838 42530
rect 31890 42478 31892 42530
rect 31836 42196 31892 42478
rect 31612 42130 31668 42140
rect 31836 42130 31892 42140
rect 32172 42532 32228 43374
rect 32284 43314 32340 43326
rect 32284 43262 32286 43314
rect 32338 43262 32340 43314
rect 32284 43204 32340 43262
rect 32284 43138 32340 43148
rect 32732 42866 32788 43484
rect 32732 42814 32734 42866
rect 32786 42814 32788 42866
rect 32732 42802 32788 42814
rect 32620 42756 32676 42766
rect 32620 42662 32676 42700
rect 31500 42030 31502 42082
rect 31554 42030 31556 42082
rect 31500 42018 31556 42030
rect 31388 41972 31444 41982
rect 31388 41878 31444 41916
rect 31500 41858 31556 41870
rect 31500 41806 31502 41858
rect 31554 41806 31556 41858
rect 31500 41186 31556 41806
rect 31500 41134 31502 41186
rect 31554 41134 31556 41186
rect 31500 41122 31556 41134
rect 31836 41188 31892 41198
rect 31836 40178 31892 41132
rect 31836 40126 31838 40178
rect 31890 40126 31892 40178
rect 31836 40114 31892 40126
rect 32172 40402 32228 42476
rect 32732 42532 32788 42542
rect 32732 42438 32788 42476
rect 32396 42196 32452 42206
rect 32396 42102 32452 42140
rect 32508 41972 32564 41982
rect 32844 41972 32900 44380
rect 33404 44370 33460 44380
rect 33516 44324 33572 44334
rect 33628 44324 33684 45052
rect 33516 44322 33684 44324
rect 33516 44270 33518 44322
rect 33570 44270 33684 44322
rect 33516 44268 33684 44270
rect 33740 45106 33796 45118
rect 33740 45054 33742 45106
rect 33794 45054 33796 45106
rect 33740 44436 33796 45054
rect 33852 45106 33908 45118
rect 33852 45054 33854 45106
rect 33906 45054 33908 45106
rect 33852 44884 33908 45054
rect 33852 44818 33908 44828
rect 33740 44324 33796 44380
rect 33964 44324 34020 44334
rect 34076 44324 34132 47966
rect 35084 48018 35140 48030
rect 35084 47966 35086 48018
rect 35138 47966 35140 48018
rect 35084 47570 35140 47966
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 42364 47684 42420 47694
rect 42252 47628 42364 47684
rect 35084 47518 35086 47570
rect 35138 47518 35140 47570
rect 35084 47506 35140 47518
rect 40572 47572 40628 47582
rect 40572 47478 40628 47516
rect 37772 47460 37828 47470
rect 36316 47346 36372 47358
rect 36316 47294 36318 47346
rect 36370 47294 36372 47346
rect 35196 47236 35252 47246
rect 34188 46900 34244 46910
rect 34188 46806 34244 46844
rect 35196 46786 35252 47180
rect 35980 47236 36036 47246
rect 35980 47142 36036 47180
rect 35196 46734 35198 46786
rect 35250 46734 35252 46786
rect 35196 46722 35252 46734
rect 34412 46676 34468 46686
rect 34412 46582 34468 46620
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 36316 45332 36372 47294
rect 36876 47236 36932 47246
rect 36428 45892 36484 45902
rect 36876 45892 36932 47180
rect 37436 47236 37492 47246
rect 37436 47234 37716 47236
rect 37436 47182 37438 47234
rect 37490 47182 37716 47234
rect 37436 47180 37716 47182
rect 37436 47170 37492 47180
rect 37324 46564 37380 46574
rect 36428 45890 36932 45892
rect 36428 45838 36430 45890
rect 36482 45838 36932 45890
rect 36428 45836 36932 45838
rect 37212 46562 37380 46564
rect 37212 46510 37326 46562
rect 37378 46510 37380 46562
rect 37212 46508 37380 46510
rect 36428 45826 36484 45836
rect 36988 45778 37044 45790
rect 36988 45726 36990 45778
rect 37042 45726 37044 45778
rect 36428 45332 36484 45342
rect 36316 45330 36484 45332
rect 36316 45278 36430 45330
rect 36482 45278 36484 45330
rect 36316 45276 36484 45278
rect 36428 45266 36484 45276
rect 35196 45220 35252 45230
rect 35084 45108 35140 45118
rect 35084 45014 35140 45052
rect 33740 44268 33908 44324
rect 33516 44258 33572 44268
rect 32956 44098 33012 44110
rect 32956 44046 32958 44098
rect 33010 44046 33012 44098
rect 32956 43764 33012 44046
rect 32956 43698 33012 43708
rect 33180 44100 33236 44110
rect 33180 43650 33236 44044
rect 33404 44098 33460 44110
rect 33404 44046 33406 44098
rect 33458 44046 33460 44098
rect 33404 43708 33460 44046
rect 33740 44100 33796 44110
rect 33740 44006 33796 44044
rect 33740 43764 33796 43774
rect 33852 43764 33908 44268
rect 33964 44322 34132 44324
rect 33964 44270 33966 44322
rect 34018 44270 34132 44322
rect 33964 44268 34132 44270
rect 33964 44258 34020 44268
rect 33964 43764 34020 43774
rect 33852 43762 34020 43764
rect 33852 43710 33966 43762
rect 34018 43710 34020 43762
rect 33852 43708 34020 43710
rect 33404 43652 33684 43708
rect 33180 43598 33182 43650
rect 33234 43598 33236 43650
rect 33180 43586 33236 43598
rect 33628 43650 33684 43652
rect 33628 43598 33630 43650
rect 33682 43598 33684 43650
rect 33628 43586 33684 43598
rect 33068 43428 33124 43438
rect 33068 43334 33124 43372
rect 33516 43428 33572 43438
rect 33740 43428 33796 43708
rect 33964 43698 34020 43708
rect 34076 43540 34132 44268
rect 34188 44996 34244 45006
rect 34188 44322 34244 44940
rect 35196 44994 35252 45164
rect 35532 45220 35588 45230
rect 35532 45218 36148 45220
rect 35532 45166 35534 45218
rect 35586 45166 36148 45218
rect 35532 45164 36148 45166
rect 35532 45154 35588 45164
rect 36092 45106 36148 45164
rect 36092 45054 36094 45106
rect 36146 45054 36148 45106
rect 36092 45042 36148 45054
rect 36204 45108 36260 45118
rect 35196 44942 35198 44994
rect 35250 44942 35252 44994
rect 35196 44930 35252 44942
rect 35868 44994 35924 45006
rect 35868 44942 35870 44994
rect 35922 44942 35924 44994
rect 35084 44884 35140 44894
rect 34188 44270 34190 44322
rect 34242 44270 34244 44322
rect 34188 44258 34244 44270
rect 34748 44436 34804 44446
rect 34188 43540 34244 43550
rect 34076 43538 34244 43540
rect 34076 43486 34190 43538
rect 34242 43486 34244 43538
rect 34076 43484 34244 43486
rect 34188 43474 34244 43484
rect 33740 43372 34132 43428
rect 33516 43334 33572 43372
rect 33852 42756 33908 42766
rect 33852 42662 33908 42700
rect 33180 42644 33236 42654
rect 33180 42642 33460 42644
rect 33180 42590 33182 42642
rect 33234 42590 33460 42642
rect 33180 42588 33460 42590
rect 33180 42578 33236 42588
rect 32956 42530 33012 42542
rect 32956 42478 32958 42530
rect 33010 42478 33012 42530
rect 32956 42196 33012 42478
rect 32956 42130 33012 42140
rect 33068 42532 33124 42542
rect 33068 41972 33124 42476
rect 32508 41970 33012 41972
rect 32508 41918 32510 41970
rect 32562 41918 33012 41970
rect 32508 41916 33012 41918
rect 32508 41906 32564 41916
rect 32396 41860 32452 41870
rect 32396 41746 32452 41804
rect 32396 41694 32398 41746
rect 32450 41694 32452 41746
rect 32396 41682 32452 41694
rect 32284 41186 32340 41198
rect 32284 41134 32286 41186
rect 32338 41134 32340 41186
rect 32284 41076 32340 41134
rect 32284 41010 32340 41020
rect 32172 40350 32174 40402
rect 32226 40350 32228 40402
rect 32172 39060 32228 40350
rect 32956 40402 33012 41916
rect 33068 41970 33236 41972
rect 33068 41918 33070 41970
rect 33122 41918 33236 41970
rect 33068 41916 33236 41918
rect 33068 41906 33124 41916
rect 32956 40350 32958 40402
rect 33010 40350 33012 40402
rect 32956 40338 33012 40350
rect 33068 40964 33124 40974
rect 32172 38966 32228 39004
rect 32284 39396 32340 39406
rect 30604 38546 30660 38556
rect 30828 38612 30996 38668
rect 31164 38612 31332 38668
rect 31724 38612 31780 38622
rect 30604 38052 30660 38062
rect 30604 37958 30660 37996
rect 30492 37762 30548 37772
rect 30380 37314 30436 37324
rect 30492 37378 30548 37390
rect 30492 37326 30494 37378
rect 30546 37326 30548 37378
rect 30156 37044 30212 37212
rect 30492 37156 30548 37326
rect 30268 37044 30324 37054
rect 30156 37042 30324 37044
rect 30156 36990 30270 37042
rect 30322 36990 30324 37042
rect 30156 36988 30324 36990
rect 30268 36978 30324 36988
rect 29484 36530 29540 36540
rect 29372 35746 29428 35756
rect 30380 36484 30436 36494
rect 29148 35634 29204 35644
rect 30268 35700 30324 35710
rect 30268 35606 30324 35644
rect 29260 35586 29316 35598
rect 29260 35534 29262 35586
rect 29314 35534 29316 35586
rect 28364 35364 28420 35374
rect 27468 35308 27636 35364
rect 27244 35196 27524 35252
rect 27468 35140 27524 35196
rect 27468 35046 27524 35084
rect 27132 34692 27188 34702
rect 27132 34690 27412 34692
rect 27132 34638 27134 34690
rect 27186 34638 27412 34690
rect 27132 34636 27412 34638
rect 27132 34626 27188 34636
rect 26460 33346 26628 33348
rect 26460 33294 26462 33346
rect 26514 33294 26628 33346
rect 26460 33292 26628 33294
rect 26460 33282 26516 33292
rect 25788 32734 25790 32786
rect 25842 32734 25844 32786
rect 25564 32562 25620 32732
rect 25788 32722 25844 32734
rect 25900 33234 25956 33246
rect 25900 33182 25902 33234
rect 25954 33182 25956 33234
rect 25564 32510 25566 32562
rect 25618 32510 25620 32562
rect 25564 32498 25620 32510
rect 25900 32452 25956 33182
rect 25788 32396 25956 32452
rect 25788 31892 25844 32396
rect 26460 32340 26516 32350
rect 25340 31668 25396 31678
rect 25340 31666 25620 31668
rect 25340 31614 25342 31666
rect 25394 31614 25620 31666
rect 25340 31612 25620 31614
rect 25340 31602 25396 31612
rect 25564 31218 25620 31612
rect 25564 31166 25566 31218
rect 25618 31166 25620 31218
rect 25564 31154 25620 31166
rect 25004 30156 25172 30212
rect 24668 29428 24724 30044
rect 24780 29988 24836 29998
rect 24780 29650 24836 29932
rect 25004 29988 25060 29998
rect 25004 29894 25060 29932
rect 24780 29598 24782 29650
rect 24834 29598 24836 29650
rect 24780 29586 24836 29598
rect 25116 29540 25172 30156
rect 24668 29362 24724 29372
rect 25004 29484 25172 29540
rect 25564 30210 25620 30222
rect 25564 30158 25566 30210
rect 25618 30158 25620 30210
rect 25564 29540 25620 30158
rect 24556 28700 24836 28756
rect 24668 28532 24724 28542
rect 23996 28530 24724 28532
rect 23996 28478 24670 28530
rect 24722 28478 24724 28530
rect 23996 28476 24724 28478
rect 24668 28466 24724 28476
rect 23324 28364 23492 28420
rect 22988 26786 23044 26796
rect 23212 28196 23268 28206
rect 23212 26516 23268 28140
rect 23212 26450 23268 26460
rect 21756 26178 21812 26190
rect 21756 26126 21758 26178
rect 21810 26126 21812 26178
rect 21756 25620 21812 26126
rect 21756 25554 21812 25564
rect 22092 26180 22148 26190
rect 22092 25618 22148 26124
rect 23100 26180 23156 26190
rect 22092 25566 22094 25618
rect 22146 25566 22148 25618
rect 22092 25554 22148 25566
rect 22204 25844 22260 25854
rect 21980 25508 22036 25518
rect 21980 25414 22036 25452
rect 22204 25506 22260 25788
rect 23100 25730 23156 26124
rect 23100 25678 23102 25730
rect 23154 25678 23156 25730
rect 23100 25666 23156 25678
rect 22204 25454 22206 25506
rect 22258 25454 22260 25506
rect 22204 25442 22260 25454
rect 22540 25506 22596 25518
rect 22540 25454 22542 25506
rect 22594 25454 22596 25506
rect 22540 25396 22596 25454
rect 21532 25340 21812 25396
rect 21420 25284 21476 25294
rect 21420 25282 21588 25284
rect 21420 25230 21422 25282
rect 21474 25230 21588 25282
rect 21420 25228 21588 25230
rect 21420 25218 21476 25228
rect 21308 24882 21364 24892
rect 21420 25060 21476 25070
rect 20972 24612 21028 24622
rect 20972 24610 21140 24612
rect 20972 24558 20974 24610
rect 21026 24558 21140 24610
rect 20972 24556 21140 24558
rect 20972 24546 21028 24556
rect 20748 23940 20804 23950
rect 20860 23940 20916 23996
rect 19404 23660 19572 23716
rect 20300 23938 20916 23940
rect 20300 23886 20750 23938
rect 20802 23886 20916 23938
rect 20300 23884 20916 23886
rect 19180 23266 19236 23278
rect 19180 23214 19182 23266
rect 19234 23214 19236 23266
rect 18956 23156 19012 23166
rect 19180 23156 19236 23214
rect 18956 23154 19180 23156
rect 18956 23102 18958 23154
rect 19010 23102 19180 23154
rect 18956 23100 19180 23102
rect 18956 23090 19012 23100
rect 19180 23090 19236 23100
rect 19404 23154 19460 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23268 19684 23278
rect 19404 23102 19406 23154
rect 19458 23102 19460 23154
rect 18508 23044 18564 23054
rect 18508 22950 18564 22988
rect 19068 22932 19124 22942
rect 18956 22930 19124 22932
rect 18956 22878 19070 22930
rect 19122 22878 19124 22930
rect 18956 22876 19124 22878
rect 18956 21812 19012 22876
rect 19068 22866 19124 22876
rect 19404 22932 19460 23102
rect 19404 22866 19460 22876
rect 19516 23266 19684 23268
rect 19516 23214 19630 23266
rect 19682 23214 19684 23266
rect 19516 23212 19684 23214
rect 19516 22484 19572 23212
rect 19628 23202 19684 23212
rect 19180 22428 19572 22484
rect 19964 23154 20020 23166
rect 19964 23102 19966 23154
rect 20018 23102 20020 23154
rect 18956 21746 19012 21756
rect 19068 22260 19124 22270
rect 18396 20802 18452 21420
rect 19068 20916 19124 22204
rect 19180 21140 19236 22428
rect 19404 22258 19460 22270
rect 19404 22206 19406 22258
rect 19458 22206 19460 22258
rect 19404 21700 19460 22206
rect 19404 21634 19460 21644
rect 19516 22148 19572 22158
rect 19964 22148 20020 23102
rect 20188 23154 20244 23166
rect 20188 23102 20190 23154
rect 20242 23102 20244 23154
rect 19516 21698 19572 22092
rect 19516 21646 19518 21698
rect 19570 21646 19572 21698
rect 19516 21634 19572 21646
rect 19628 22092 20020 22148
rect 20076 23042 20132 23054
rect 20076 22990 20078 23042
rect 20130 22990 20132 23042
rect 20076 22148 20132 22990
rect 20188 22708 20244 23102
rect 20188 22642 20244 22652
rect 20188 22372 20244 22382
rect 20300 22372 20356 23884
rect 20748 23874 20804 23884
rect 20636 23156 20692 23166
rect 20636 23154 20916 23156
rect 20636 23102 20638 23154
rect 20690 23102 20916 23154
rect 20636 23100 20916 23102
rect 20636 23090 20692 23100
rect 20636 22708 20692 22718
rect 20636 22482 20692 22652
rect 20636 22430 20638 22482
rect 20690 22430 20692 22482
rect 20636 22418 20692 22430
rect 20188 22370 20356 22372
rect 20188 22318 20190 22370
rect 20242 22318 20356 22370
rect 20188 22316 20356 22318
rect 20188 22306 20244 22316
rect 19628 21476 19684 22092
rect 20076 22082 20132 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20300 21586 20356 22316
rect 20860 22036 20916 23100
rect 20972 23044 21028 23054
rect 20972 22950 21028 22988
rect 21084 22260 21140 24556
rect 21196 23156 21252 23166
rect 21196 22596 21252 23100
rect 21308 23044 21364 23054
rect 21420 23044 21476 25004
rect 21532 24276 21588 25228
rect 21532 24210 21588 24220
rect 21644 25172 21700 25182
rect 21644 24498 21700 25116
rect 21644 24446 21646 24498
rect 21698 24446 21700 24498
rect 21532 24052 21588 24062
rect 21532 23958 21588 23996
rect 21308 23042 21476 23044
rect 21308 22990 21310 23042
rect 21362 22990 21476 23042
rect 21308 22988 21476 22990
rect 21308 22978 21364 22988
rect 21644 22708 21700 24446
rect 21644 22642 21700 22652
rect 21196 22540 21476 22596
rect 21420 22484 21476 22540
rect 21756 22484 21812 25340
rect 22540 25330 22596 25340
rect 22876 25508 22932 25518
rect 23324 25508 23380 28364
rect 24108 28308 24164 28318
rect 23884 27748 23940 27758
rect 23884 27654 23940 27692
rect 23436 26964 23492 27002
rect 23436 26898 23492 26908
rect 24108 26908 24164 28252
rect 24668 27860 24724 27870
rect 24780 27860 24836 28700
rect 24668 27858 24780 27860
rect 24668 27806 24670 27858
rect 24722 27806 24780 27858
rect 24668 27804 24780 27806
rect 24220 27076 24276 27086
rect 24668 27076 24724 27804
rect 24780 27766 24836 27804
rect 24892 27636 24948 27646
rect 24892 27186 24948 27580
rect 24892 27134 24894 27186
rect 24946 27134 24948 27186
rect 24892 27122 24948 27134
rect 24220 27074 24724 27076
rect 24220 27022 24222 27074
rect 24274 27022 24724 27074
rect 24220 27020 24724 27022
rect 24220 27010 24276 27020
rect 24108 26852 24612 26908
rect 23884 26180 23940 26190
rect 23884 26086 23940 26124
rect 23996 26068 24052 26078
rect 23996 25732 24052 26012
rect 23884 25676 24388 25732
rect 22428 25284 22484 25322
rect 22428 25218 22484 25228
rect 22652 25284 22708 25294
rect 22428 25060 22484 25070
rect 22428 24834 22484 25004
rect 22652 24946 22708 25228
rect 22652 24894 22654 24946
rect 22706 24894 22708 24946
rect 22652 24882 22708 24894
rect 22764 24948 22820 24958
rect 22876 24948 22932 25452
rect 23100 25452 23380 25508
rect 23436 25620 23492 25630
rect 23436 25506 23492 25564
rect 23436 25454 23438 25506
rect 23490 25454 23492 25506
rect 22988 25396 23044 25406
rect 22988 25302 23044 25340
rect 22988 24948 23044 24958
rect 22876 24946 23044 24948
rect 22876 24894 22990 24946
rect 23042 24894 23044 24946
rect 22876 24892 23044 24894
rect 22764 24854 22820 24892
rect 22988 24882 23044 24892
rect 22428 24782 22430 24834
rect 22482 24782 22484 24834
rect 22428 24770 22484 24782
rect 22876 24722 22932 24734
rect 22876 24670 22878 24722
rect 22930 24670 22932 24722
rect 22876 23940 22932 24670
rect 22876 23874 22932 23884
rect 21420 22482 21700 22484
rect 21420 22430 21422 22482
rect 21474 22430 21700 22482
rect 21420 22428 21700 22430
rect 21420 22418 21476 22428
rect 21084 22194 21140 22204
rect 20860 21980 21364 22036
rect 20860 21812 20916 21822
rect 21308 21812 21364 21980
rect 21308 21756 21476 21812
rect 20860 21718 20916 21756
rect 21196 21700 21252 21710
rect 21196 21606 21252 21644
rect 21084 21588 21140 21598
rect 20300 21534 20302 21586
rect 20354 21534 20356 21586
rect 20300 21522 20356 21534
rect 20860 21586 21140 21588
rect 20860 21534 21086 21586
rect 21138 21534 21140 21586
rect 20860 21532 21140 21534
rect 19628 21410 19684 21420
rect 20412 21476 20468 21486
rect 19180 21074 19236 21084
rect 19292 20916 19348 20926
rect 19068 20914 19348 20916
rect 19068 20862 19294 20914
rect 19346 20862 19348 20914
rect 19068 20860 19348 20862
rect 19292 20850 19348 20860
rect 18396 20750 18398 20802
rect 18450 20750 18452 20802
rect 18396 20738 18452 20750
rect 18732 20802 18788 20814
rect 18732 20750 18734 20802
rect 18786 20750 18788 20802
rect 18732 20188 18788 20750
rect 18956 20802 19012 20814
rect 18956 20750 18958 20802
rect 19010 20750 19012 20802
rect 18956 20188 19012 20750
rect 19740 20804 19796 20814
rect 19740 20710 19796 20748
rect 19628 20692 19684 20702
rect 19628 20578 19684 20636
rect 20412 20690 20468 21420
rect 20412 20638 20414 20690
rect 20466 20638 20468 20690
rect 20412 20626 20468 20638
rect 20748 20692 20804 20702
rect 20748 20598 20804 20636
rect 19628 20526 19630 20578
rect 19682 20526 19684 20578
rect 19516 20356 19572 20366
rect 18732 20132 18900 20188
rect 18956 20132 19348 20188
rect 18732 19906 18788 19918
rect 18732 19854 18734 19906
rect 18786 19854 18788 19906
rect 18172 15596 18340 15652
rect 18396 19348 18452 19358
rect 18396 17666 18452 19292
rect 18732 19236 18788 19854
rect 18732 19170 18788 19180
rect 18732 18676 18788 18686
rect 18508 18562 18564 18574
rect 18508 18510 18510 18562
rect 18562 18510 18564 18562
rect 18508 18004 18564 18510
rect 18620 18564 18676 18574
rect 18732 18564 18788 18620
rect 18620 18562 18788 18564
rect 18620 18510 18622 18562
rect 18674 18510 18788 18562
rect 18620 18508 18788 18510
rect 18620 18498 18676 18508
rect 18620 18340 18676 18350
rect 18620 18226 18676 18284
rect 18620 18174 18622 18226
rect 18674 18174 18676 18226
rect 18620 18162 18676 18174
rect 18508 17938 18564 17948
rect 18396 17614 18398 17666
rect 18450 17614 18452 17666
rect 18060 15316 18116 15326
rect 18060 15222 18116 15260
rect 17948 15138 18004 15148
rect 17276 14590 17278 14642
rect 17330 14590 17332 14642
rect 17276 14578 17332 14590
rect 17388 15090 17444 15102
rect 17388 15038 17390 15090
rect 17442 15038 17444 15090
rect 17388 14084 17444 15038
rect 18172 15090 18228 15596
rect 18396 15540 18452 17614
rect 18620 16212 18676 16222
rect 18732 16212 18788 18508
rect 18844 18116 18900 20132
rect 19068 19906 19124 19918
rect 19068 19854 19070 19906
rect 19122 19854 19124 19906
rect 19068 19460 19124 19854
rect 19068 18340 19124 19404
rect 19180 18564 19236 18574
rect 19180 18470 19236 18508
rect 19292 18450 19348 20132
rect 19404 18676 19460 18686
rect 19404 18582 19460 18620
rect 19292 18398 19294 18450
rect 19346 18398 19348 18450
rect 19292 18386 19348 18398
rect 19068 18284 19236 18340
rect 19068 18116 19124 18126
rect 18844 18060 19068 18116
rect 19068 17890 19124 18060
rect 19068 17838 19070 17890
rect 19122 17838 19124 17890
rect 19068 17826 19124 17838
rect 19180 17780 19236 18284
rect 19404 17780 19460 17790
rect 19180 17724 19404 17780
rect 19404 17686 19460 17724
rect 18956 17108 19012 17118
rect 18676 16156 18788 16212
rect 18844 16324 18900 16334
rect 18620 16146 18676 16156
rect 18844 15540 18900 16268
rect 18172 15038 18174 15090
rect 18226 15038 18228 15090
rect 18172 15026 18228 15038
rect 18284 15484 18396 15540
rect 17948 14868 18004 14878
rect 17948 14642 18004 14812
rect 17948 14590 17950 14642
rect 18002 14590 18004 14642
rect 17948 14578 18004 14590
rect 16828 14028 17444 14084
rect 18172 14308 18228 14318
rect 16828 13970 16884 14028
rect 16828 13918 16830 13970
rect 16882 13918 16884 13970
rect 16268 13458 16324 13468
rect 16604 13636 16660 13646
rect 15708 12178 16100 12180
rect 15708 12126 15710 12178
rect 15762 12126 16100 12178
rect 15708 12124 16100 12126
rect 16380 12964 16436 12974
rect 16380 12404 16436 12908
rect 16380 12178 16436 12348
rect 16380 12126 16382 12178
rect 16434 12126 16436 12178
rect 15708 12114 15764 12124
rect 16268 11956 16324 11966
rect 15484 11954 16324 11956
rect 15484 11902 16270 11954
rect 16322 11902 16324 11954
rect 15484 11900 16324 11902
rect 16268 11890 16324 11900
rect 16380 11732 16436 12126
rect 16604 12178 16660 13580
rect 16828 12964 16884 13918
rect 17276 13746 17332 13758
rect 17276 13694 17278 13746
rect 17330 13694 17332 13746
rect 17276 13524 17332 13694
rect 17612 13748 17668 13758
rect 17612 13654 17668 13692
rect 17948 13746 18004 13758
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17500 13636 17556 13646
rect 17500 13542 17556 13580
rect 17276 13458 17332 13468
rect 17948 13188 18004 13694
rect 17276 13132 18004 13188
rect 17276 13074 17332 13132
rect 17276 13022 17278 13074
rect 17330 13022 17332 13074
rect 17276 13010 17332 13022
rect 16828 12898 16884 12908
rect 17724 12962 17780 12974
rect 17724 12910 17726 12962
rect 17778 12910 17780 12962
rect 17724 12852 17780 12910
rect 16604 12126 16606 12178
rect 16658 12126 16660 12178
rect 16604 12114 16660 12126
rect 16716 12180 16772 12190
rect 17388 12180 17444 12190
rect 16772 12124 16884 12180
rect 16716 12086 16772 12124
rect 16380 11666 16436 11676
rect 16716 10836 16772 10846
rect 16716 10742 16772 10780
rect 16828 10834 16884 12124
rect 17388 12086 17444 12124
rect 16828 10782 16830 10834
rect 16882 10782 16884 10834
rect 15372 10546 15428 10556
rect 16156 10612 16212 10622
rect 16156 10518 16212 10556
rect 16604 10610 16660 10622
rect 16604 10558 16606 10610
rect 16658 10558 16660 10610
rect 15932 10500 15988 10510
rect 15260 9886 15262 9938
rect 15314 9886 15316 9938
rect 15260 9874 15316 9886
rect 15708 10444 15932 10500
rect 15596 9828 15652 9838
rect 15596 9734 15652 9772
rect 15708 9826 15764 10444
rect 15932 10406 15988 10444
rect 16604 10500 16660 10558
rect 16604 10434 16660 10444
rect 16828 10276 16884 10782
rect 15708 9774 15710 9826
rect 15762 9774 15764 9826
rect 15708 9762 15764 9774
rect 15820 10220 16884 10276
rect 16940 11620 16996 11630
rect 15820 9826 15876 10220
rect 15820 9774 15822 9826
rect 15874 9774 15876 9826
rect 15820 9762 15876 9774
rect 16044 10052 16100 10062
rect 14812 9602 14868 9614
rect 14812 9550 14814 9602
rect 14866 9550 14868 9602
rect 14812 8484 14868 9550
rect 16044 9268 16100 9996
rect 16828 9826 16884 9838
rect 16828 9774 16830 9826
rect 16882 9774 16884 9826
rect 16268 9604 16324 9614
rect 16268 9602 16436 9604
rect 16268 9550 16270 9602
rect 16322 9550 16436 9602
rect 16268 9548 16436 9550
rect 16268 9538 16324 9548
rect 16044 9174 16100 9212
rect 15260 9154 15316 9166
rect 15260 9102 15262 9154
rect 15314 9102 15316 9154
rect 14812 8418 14868 8428
rect 15036 8932 15092 8942
rect 15036 8372 15092 8876
rect 15036 8306 15092 8316
rect 14812 8148 14868 8158
rect 15148 8148 15204 8158
rect 14812 8146 15204 8148
rect 14812 8094 14814 8146
rect 14866 8094 15150 8146
rect 15202 8094 15204 8146
rect 14812 8092 15204 8094
rect 14812 8082 14868 8092
rect 15148 8082 15204 8092
rect 14700 7140 14756 7420
rect 14700 7074 14756 7084
rect 14588 6692 14644 6702
rect 14588 6598 14644 6636
rect 15260 6690 15316 9102
rect 16380 9154 16436 9548
rect 16380 9102 16382 9154
rect 16434 9102 16436 9154
rect 16380 9090 16436 9102
rect 16716 9154 16772 9166
rect 16716 9102 16718 9154
rect 16770 9102 16772 9154
rect 15596 9042 15652 9054
rect 15596 8990 15598 9042
rect 15650 8990 15652 9042
rect 15260 6638 15262 6690
rect 15314 6638 15316 6690
rect 15260 6626 15316 6638
rect 15372 8372 15428 8382
rect 15372 8034 15428 8316
rect 15372 7982 15374 8034
rect 15426 7982 15428 8034
rect 15372 7252 15428 7982
rect 15484 8370 15540 8382
rect 15484 8318 15486 8370
rect 15538 8318 15540 8370
rect 15484 7700 15540 8318
rect 15596 7924 15652 8990
rect 16492 8372 16548 8382
rect 16156 8260 16212 8270
rect 16156 8166 16212 8204
rect 16492 8036 16548 8316
rect 16716 8372 16772 9102
rect 16716 8306 16772 8316
rect 16492 7970 16548 7980
rect 16828 8260 16884 9774
rect 16940 9828 16996 11564
rect 17724 10612 17780 12796
rect 17948 12290 18004 13132
rect 17948 12238 17950 12290
rect 18002 12238 18004 12290
rect 17948 12226 18004 12238
rect 18060 13748 18116 13758
rect 18060 12290 18116 13692
rect 18060 12238 18062 12290
rect 18114 12238 18116 12290
rect 18060 12226 18116 12238
rect 17836 12178 17892 12190
rect 17836 12126 17838 12178
rect 17890 12126 17892 12178
rect 17836 11956 17892 12126
rect 18172 11956 18228 14252
rect 17836 11900 18228 11956
rect 17724 10518 17780 10556
rect 18284 11508 18340 15484
rect 18396 15474 18452 15484
rect 18620 15484 18900 15540
rect 18396 15316 18452 15326
rect 18620 15316 18676 15484
rect 18396 15314 18676 15316
rect 18396 15262 18398 15314
rect 18450 15262 18676 15314
rect 18396 15260 18676 15262
rect 18732 15316 18788 15326
rect 18844 15316 18900 15326
rect 18788 15314 18900 15316
rect 18788 15262 18846 15314
rect 18898 15262 18900 15314
rect 18788 15260 18900 15262
rect 18396 15250 18452 15260
rect 18508 14308 18564 14318
rect 18508 14306 18676 14308
rect 18508 14254 18510 14306
rect 18562 14254 18676 14306
rect 18508 14252 18676 14254
rect 18508 14242 18564 14252
rect 18620 13858 18676 14252
rect 18620 13806 18622 13858
rect 18674 13806 18676 13858
rect 18508 13522 18564 13534
rect 18508 13470 18510 13522
rect 18562 13470 18564 13522
rect 18508 13074 18564 13470
rect 18620 13524 18676 13806
rect 18620 13458 18676 13468
rect 18732 13188 18788 15260
rect 18844 15250 18900 15260
rect 18956 14980 19012 17052
rect 19516 15652 19572 20300
rect 19628 17778 19684 20526
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20860 20188 20916 21532
rect 21084 21522 21140 21532
rect 21308 21586 21364 21598
rect 21308 21534 21310 21586
rect 21362 21534 21364 21586
rect 21308 21476 21364 21534
rect 21308 21410 21364 21420
rect 21420 20914 21476 21756
rect 21420 20862 21422 20914
rect 21474 20862 21476 20914
rect 21420 20850 21476 20862
rect 21532 21364 21588 21374
rect 21532 20802 21588 21308
rect 21532 20750 21534 20802
rect 21586 20750 21588 20802
rect 21532 20738 21588 20750
rect 21308 20580 21364 20590
rect 21644 20580 21700 22428
rect 21756 22390 21812 22428
rect 22876 22820 22932 22830
rect 22764 22260 22820 22270
rect 21756 21588 21812 21598
rect 21756 21494 21812 21532
rect 22428 21474 22484 21486
rect 22428 21422 22430 21474
rect 22482 21422 22484 21474
rect 21756 21140 21812 21150
rect 21756 20802 21812 21084
rect 21756 20750 21758 20802
rect 21810 20750 21812 20802
rect 21756 20738 21812 20750
rect 22316 20916 22372 20926
rect 21308 20578 21700 20580
rect 21308 20526 21310 20578
rect 21362 20526 21700 20578
rect 21308 20524 21700 20526
rect 21308 20188 21364 20524
rect 20412 20132 20916 20188
rect 20972 20132 21364 20188
rect 20076 19236 20132 19246
rect 20076 19142 20132 19180
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19740 18452 19796 18462
rect 19740 18358 19796 18396
rect 20188 18338 20244 18350
rect 20188 18286 20190 18338
rect 20242 18286 20244 18338
rect 20076 18228 20132 18238
rect 20076 18134 20132 18172
rect 20188 18004 20244 18286
rect 20188 17938 20244 17948
rect 20412 18340 20468 20132
rect 19628 17726 19630 17778
rect 19682 17726 19684 17778
rect 19628 17714 19684 17726
rect 20188 17668 20244 17678
rect 20188 17574 20244 17612
rect 20412 17666 20468 18284
rect 20972 18004 21028 20132
rect 21980 20020 22036 20030
rect 21980 19926 22036 19964
rect 21196 19908 21252 19918
rect 21196 19906 21476 19908
rect 21196 19854 21198 19906
rect 21250 19854 21476 19906
rect 21196 19852 21476 19854
rect 21196 19842 21252 19852
rect 21308 19348 21364 19358
rect 21308 19234 21364 19292
rect 21420 19346 21476 19852
rect 21420 19294 21422 19346
rect 21474 19294 21476 19346
rect 21420 19282 21476 19294
rect 21756 19348 21812 19358
rect 21308 19182 21310 19234
rect 21362 19182 21364 19234
rect 21308 19170 21364 19182
rect 21532 19236 21588 19246
rect 21532 18788 21588 19180
rect 21084 18732 21588 18788
rect 21084 18674 21140 18732
rect 21084 18622 21086 18674
rect 21138 18622 21140 18674
rect 21084 18610 21140 18622
rect 20412 17614 20414 17666
rect 20466 17614 20468 17666
rect 20412 17602 20468 17614
rect 20748 17948 21028 18004
rect 21308 18338 21364 18350
rect 21308 18286 21310 18338
rect 21362 18286 21364 18338
rect 21308 18004 21364 18286
rect 20300 17442 20356 17454
rect 20300 17390 20302 17442
rect 20354 17390 20356 17442
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20300 16994 20356 17390
rect 20300 16942 20302 16994
rect 20354 16942 20356 16994
rect 20300 16930 20356 16942
rect 19964 16772 20020 16782
rect 19964 16210 20020 16716
rect 20748 16324 20804 17948
rect 21308 17938 21364 17948
rect 21420 17780 21476 17790
rect 20860 17778 21476 17780
rect 20860 17726 21422 17778
rect 21474 17726 21476 17778
rect 20860 17724 21476 17726
rect 20860 17666 20916 17724
rect 21420 17714 21476 17724
rect 21756 17668 21812 19292
rect 21868 19236 21924 19246
rect 22092 19236 22148 19246
rect 21868 19234 22148 19236
rect 21868 19182 21870 19234
rect 21922 19182 22094 19234
rect 22146 19182 22148 19234
rect 21868 19180 22148 19182
rect 21868 19170 21924 19180
rect 22092 19170 22148 19180
rect 22316 19236 22372 20860
rect 22428 19908 22484 21422
rect 22652 21476 22708 21486
rect 22652 20802 22708 21420
rect 22764 20914 22820 22204
rect 22764 20862 22766 20914
rect 22818 20862 22820 20914
rect 22764 20850 22820 20862
rect 22876 20916 22932 22764
rect 22652 20750 22654 20802
rect 22706 20750 22708 20802
rect 22652 20130 22708 20750
rect 22876 20802 22932 20860
rect 22876 20750 22878 20802
rect 22930 20750 22932 20802
rect 22876 20738 22932 20750
rect 22988 21252 23044 21262
rect 23100 21252 23156 25452
rect 23436 25442 23492 25454
rect 23884 25506 23940 25676
rect 23884 25454 23886 25506
rect 23938 25454 23940 25506
rect 23884 25442 23940 25454
rect 23996 25508 24052 25518
rect 23996 25414 24052 25452
rect 23772 25396 23828 25406
rect 23772 25302 23828 25340
rect 23660 25284 23716 25294
rect 23660 25190 23716 25228
rect 24332 24948 24388 25676
rect 24444 25284 24500 25294
rect 24444 25190 24500 25228
rect 24444 24948 24500 24958
rect 24332 24946 24500 24948
rect 24332 24894 24446 24946
rect 24498 24894 24500 24946
rect 24332 24892 24500 24894
rect 24444 24882 24500 24892
rect 23884 24724 23940 24734
rect 23884 24630 23940 24668
rect 23436 24276 23492 24286
rect 23436 23266 23492 24220
rect 23436 23214 23438 23266
rect 23490 23214 23492 23266
rect 23436 23202 23492 23214
rect 24220 23154 24276 23166
rect 24220 23102 24222 23154
rect 24274 23102 24276 23154
rect 23772 22484 23828 22494
rect 24220 22484 24276 23102
rect 23548 21812 23604 21822
rect 23324 21364 23380 21374
rect 23044 21196 23156 21252
rect 23212 21252 23268 21262
rect 22652 20078 22654 20130
rect 22706 20078 22708 20130
rect 22652 20066 22708 20078
rect 22876 20018 22932 20030
rect 22876 19966 22878 20018
rect 22930 19966 22932 20018
rect 22764 19908 22820 19918
rect 22428 19906 22820 19908
rect 22428 19854 22766 19906
rect 22818 19854 22820 19906
rect 22428 19852 22820 19854
rect 22764 19842 22820 19852
rect 22316 19170 22372 19180
rect 22428 19460 22484 19470
rect 22428 19234 22484 19404
rect 22428 19182 22430 19234
rect 22482 19182 22484 19234
rect 22428 19170 22484 19182
rect 22764 19234 22820 19246
rect 22764 19182 22766 19234
rect 22818 19182 22820 19234
rect 22764 19124 22820 19182
rect 22764 19058 22820 19068
rect 22204 19010 22260 19022
rect 22204 18958 22206 19010
rect 22258 18958 22260 19010
rect 22204 18452 22260 18958
rect 22876 18900 22932 19966
rect 22988 19796 23044 21196
rect 23212 20692 23268 21196
rect 23100 20578 23156 20590
rect 23100 20526 23102 20578
rect 23154 20526 23156 20578
rect 23100 20132 23156 20526
rect 23100 20066 23156 20076
rect 22988 19740 23156 19796
rect 22988 19572 23044 19582
rect 22988 19122 23044 19516
rect 22988 19070 22990 19122
rect 23042 19070 23044 19122
rect 22988 19058 23044 19070
rect 20860 17614 20862 17666
rect 20914 17614 20916 17666
rect 20860 17602 20916 17614
rect 21644 17612 21756 17668
rect 21308 17556 21364 17566
rect 21084 16882 21140 16894
rect 21084 16830 21086 16882
rect 21138 16830 21140 16882
rect 20748 16268 20916 16324
rect 19964 16158 19966 16210
rect 20018 16158 20020 16210
rect 19964 16146 20020 16158
rect 20748 16098 20804 16110
rect 20748 16046 20750 16098
rect 20802 16046 20804 16098
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19516 15596 19684 15652
rect 19836 15642 20100 15652
rect 19404 15540 19460 15550
rect 19628 15540 19684 15596
rect 20076 15540 20132 15550
rect 20524 15540 20580 15550
rect 19628 15538 20468 15540
rect 19628 15486 20078 15538
rect 20130 15486 20468 15538
rect 19628 15484 20468 15486
rect 19404 15446 19460 15484
rect 20076 15474 20132 15484
rect 18956 14914 19012 14924
rect 20412 14980 20468 15484
rect 20524 15446 20580 15484
rect 20748 15092 20804 16046
rect 20748 15026 20804 15036
rect 20860 15538 20916 16268
rect 20860 15486 20862 15538
rect 20914 15486 20916 15538
rect 19852 14532 19908 14542
rect 19404 14530 19908 14532
rect 19404 14478 19854 14530
rect 19906 14478 19908 14530
rect 19404 14476 19908 14478
rect 19292 14306 19348 14318
rect 19292 14254 19294 14306
rect 19346 14254 19348 14306
rect 19292 13748 19348 14254
rect 19404 13748 19460 14476
rect 19852 14466 19908 14476
rect 20076 14530 20132 14542
rect 20076 14478 20078 14530
rect 20130 14478 20132 14530
rect 19516 14308 19572 14318
rect 20076 14308 20132 14478
rect 20412 14530 20468 14924
rect 20412 14478 20414 14530
rect 20466 14478 20468 14530
rect 20412 14466 20468 14478
rect 19516 14214 19572 14252
rect 19628 14252 20132 14308
rect 20748 14306 20804 14318
rect 20748 14254 20750 14306
rect 20802 14254 20804 14306
rect 19628 13972 19684 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13916 19796 13972
rect 19516 13748 19572 13758
rect 19404 13746 19572 13748
rect 19404 13694 19518 13746
rect 19570 13694 19572 13746
rect 19404 13692 19572 13694
rect 19292 13682 19348 13692
rect 18956 13636 19012 13646
rect 18844 13580 18956 13636
rect 18844 13522 18900 13580
rect 18956 13570 19012 13580
rect 18844 13470 18846 13522
rect 18898 13470 18900 13522
rect 18844 13458 18900 13470
rect 18732 13122 18788 13132
rect 18508 13022 18510 13074
rect 18562 13022 18564 13074
rect 18508 13010 18564 13022
rect 19516 12740 19572 13692
rect 19740 13746 19796 13916
rect 19740 13694 19742 13746
rect 19794 13694 19796 13746
rect 19628 13636 19684 13646
rect 19628 13542 19684 13580
rect 19740 13076 19796 13694
rect 19740 13010 19796 13020
rect 20076 13746 20132 13758
rect 20076 13694 20078 13746
rect 20130 13694 20132 13746
rect 20076 12740 20132 13694
rect 20412 13746 20468 13758
rect 20412 13694 20414 13746
rect 20466 13694 20468 13746
rect 20412 12852 20468 13694
rect 20748 13636 20804 14254
rect 20748 13570 20804 13580
rect 20636 13076 20692 13086
rect 20636 12982 20692 13020
rect 20412 12786 20468 12796
rect 20076 12684 20244 12740
rect 19516 12674 19572 12684
rect 20188 12628 20244 12684
rect 19836 12572 20100 12582
rect 20188 12572 20468 12628
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19068 12180 19124 12190
rect 19740 12180 19796 12190
rect 18956 12178 19796 12180
rect 18956 12126 19070 12178
rect 19122 12126 19742 12178
rect 19794 12126 19796 12178
rect 18956 12124 19796 12126
rect 18844 12068 18900 12078
rect 18844 11974 18900 12012
rect 18284 11394 18340 11452
rect 18284 11342 18286 11394
rect 18338 11342 18340 11394
rect 18284 10052 18340 11342
rect 18396 11956 18452 11966
rect 18396 10722 18452 11900
rect 18396 10670 18398 10722
rect 18450 10670 18452 10722
rect 18396 10658 18452 10670
rect 18844 10052 18900 10062
rect 18956 10052 19012 12124
rect 19068 12114 19124 12124
rect 19740 12114 19796 12124
rect 20300 12066 20356 12078
rect 20300 12014 20302 12066
rect 20354 12014 20356 12066
rect 19068 11956 19124 11966
rect 19068 11862 19124 11900
rect 19404 11956 19460 11966
rect 19404 11954 19684 11956
rect 19404 11902 19406 11954
rect 19458 11902 19684 11954
rect 19404 11900 19684 11902
rect 19404 11890 19460 11900
rect 19180 11508 19236 11518
rect 19628 11508 19684 11900
rect 20076 11954 20132 11966
rect 20076 11902 20078 11954
rect 20130 11902 20132 11954
rect 19852 11508 19908 11518
rect 19628 11506 19908 11508
rect 19628 11454 19854 11506
rect 19906 11454 19908 11506
rect 19628 11452 19908 11454
rect 19180 11414 19236 11452
rect 19852 11442 19908 11452
rect 19964 11396 20020 11406
rect 19964 11302 20020 11340
rect 19740 11172 19796 11182
rect 20076 11172 20132 11902
rect 18340 9996 18452 10052
rect 18284 9986 18340 9996
rect 16940 9762 16996 9772
rect 17612 9716 17668 9726
rect 17612 9714 18228 9716
rect 17612 9662 17614 9714
rect 17666 9662 18228 9714
rect 17612 9660 18228 9662
rect 17612 9650 17668 9660
rect 17164 9156 17220 9166
rect 16940 8372 16996 8382
rect 16940 8278 16996 8316
rect 15596 7858 15652 7868
rect 15484 7644 16100 7700
rect 16044 7586 16100 7644
rect 16044 7534 16046 7586
rect 16098 7534 16100 7586
rect 16044 7522 16100 7534
rect 16828 7474 16884 8204
rect 16940 8148 16996 8158
rect 16996 8092 17108 8148
rect 16940 8082 16996 8092
rect 16828 7422 16830 7474
rect 16882 7422 16884 7474
rect 16828 7364 16884 7422
rect 15484 7252 15540 7262
rect 15372 7196 15484 7252
rect 15372 6468 15428 7196
rect 15484 7186 15540 7196
rect 14364 5854 14366 5906
rect 14418 5854 14420 5906
rect 14364 5842 14420 5854
rect 15148 6412 15428 6468
rect 15596 7140 15652 7150
rect 13916 5796 13972 5806
rect 13692 5124 13748 5134
rect 13692 5030 13748 5068
rect 13916 5122 13972 5740
rect 13916 5070 13918 5122
rect 13970 5070 13972 5122
rect 13468 4286 13470 4338
rect 13522 4286 13524 4338
rect 13468 4274 13524 4286
rect 13916 4226 13972 5070
rect 14588 5124 14644 5134
rect 14924 5124 14980 5134
rect 14588 5122 14980 5124
rect 14588 5070 14590 5122
rect 14642 5070 14926 5122
rect 14978 5070 14980 5122
rect 14588 5068 14980 5070
rect 14588 5058 14644 5068
rect 14924 5058 14980 5068
rect 15148 5010 15204 6412
rect 15596 6132 15652 7084
rect 15596 6066 15652 6076
rect 16268 7140 16324 7150
rect 16156 6020 16212 6030
rect 16156 5906 16212 5964
rect 16156 5854 16158 5906
rect 16210 5854 16212 5906
rect 16156 5842 16212 5854
rect 16268 5794 16324 7084
rect 16268 5742 16270 5794
rect 16322 5742 16324 5794
rect 16268 5730 16324 5742
rect 16828 6692 16884 7308
rect 16716 5682 16772 5694
rect 16716 5630 16718 5682
rect 16770 5630 16772 5682
rect 15260 5236 15316 5246
rect 15260 5234 15540 5236
rect 15260 5182 15262 5234
rect 15314 5182 15540 5234
rect 15260 5180 15540 5182
rect 15260 5170 15316 5180
rect 15148 4958 15150 5010
rect 15202 4958 15204 5010
rect 15148 4946 15204 4958
rect 15484 4676 15540 5180
rect 15596 5234 15652 5246
rect 15596 5182 15598 5234
rect 15650 5182 15652 5234
rect 15596 4900 15652 5182
rect 15596 4834 15652 4844
rect 15484 4620 16100 4676
rect 16044 4450 16100 4620
rect 16044 4398 16046 4450
rect 16098 4398 16100 4450
rect 16044 4386 16100 4398
rect 16716 4340 16772 5630
rect 16716 4274 16772 4284
rect 16828 4338 16884 6636
rect 16940 5908 16996 5918
rect 16940 5814 16996 5852
rect 16828 4286 16830 4338
rect 16882 4286 16884 4338
rect 16828 4274 16884 4286
rect 13916 4174 13918 4226
rect 13970 4174 13972 4226
rect 13916 4162 13972 4174
rect 13244 3726 13246 3778
rect 13298 3726 13300 3778
rect 13244 3714 13300 3726
rect 13692 3556 13748 3566
rect 13132 3500 13300 3556
rect 13244 3442 13300 3500
rect 13132 3388 13188 3398
rect 13020 3386 13188 3388
rect 13020 3334 13134 3386
rect 13186 3334 13188 3386
rect 13244 3390 13246 3442
rect 13298 3390 13300 3442
rect 13244 3378 13300 3390
rect 13020 3332 13188 3334
rect 13132 3322 13188 3332
rect 12236 2996 12292 3006
rect 12124 2940 12236 2996
rect 12236 2930 12292 2940
rect 13692 800 13748 3500
rect 16380 3556 16436 3566
rect 16380 3462 16436 3500
rect 17052 3554 17108 8092
rect 17164 5796 17220 9100
rect 17500 8930 17556 8942
rect 17500 8878 17502 8930
rect 17554 8878 17556 8930
rect 17388 8818 17444 8830
rect 17388 8766 17390 8818
rect 17442 8766 17444 8818
rect 17388 7140 17444 8766
rect 17388 7074 17444 7084
rect 17388 6804 17444 6814
rect 17500 6804 17556 8878
rect 18172 8930 18228 9660
rect 18284 9604 18340 9614
rect 18284 9266 18340 9548
rect 18284 9214 18286 9266
rect 18338 9214 18340 9266
rect 18284 9202 18340 9214
rect 18172 8878 18174 8930
rect 18226 8878 18228 8930
rect 18172 8866 18228 8878
rect 18396 8596 18452 9996
rect 18900 9996 19012 10052
rect 19516 11170 20132 11172
rect 19516 11118 19742 11170
rect 19794 11118 20132 11170
rect 19516 11116 20132 11118
rect 20300 11396 20356 12014
rect 18844 9266 18900 9996
rect 19516 9716 19572 11116
rect 19740 11106 19796 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20300 10500 20356 11340
rect 20412 11844 20468 12572
rect 20412 11394 20468 11788
rect 20860 11732 20916 15486
rect 21084 15092 21140 16830
rect 21196 16212 21252 16222
rect 21196 15538 21252 16156
rect 21308 16098 21364 17500
rect 21532 17444 21588 17454
rect 21532 17350 21588 17388
rect 21420 17108 21476 17118
rect 21644 17108 21700 17612
rect 21756 17602 21812 17612
rect 21980 18396 22260 18452
rect 22316 18844 22932 18900
rect 21756 17442 21812 17454
rect 21756 17390 21758 17442
rect 21810 17390 21812 17442
rect 21756 17332 21812 17390
rect 21980 17332 22036 18396
rect 22316 18116 22372 18844
rect 22204 17780 22260 17790
rect 22204 17686 22260 17724
rect 22092 17668 22148 17678
rect 22092 17574 22148 17612
rect 22316 17666 22372 18060
rect 22316 17614 22318 17666
rect 22370 17614 22372 17666
rect 22316 17602 22372 17614
rect 22652 17668 22708 17678
rect 22876 17668 22932 17678
rect 22652 17666 22932 17668
rect 22652 17614 22654 17666
rect 22706 17614 22878 17666
rect 22930 17614 22932 17666
rect 22652 17612 22932 17614
rect 22652 17602 22708 17612
rect 22876 17602 22932 17612
rect 21756 17276 22036 17332
rect 21420 17106 21700 17108
rect 21420 17054 21422 17106
rect 21474 17054 21700 17106
rect 21420 17052 21700 17054
rect 21980 17108 22036 17276
rect 22988 17442 23044 17454
rect 22988 17390 22990 17442
rect 23042 17390 23044 17442
rect 22316 17108 22372 17118
rect 22988 17108 23044 17390
rect 21980 17106 23044 17108
rect 21980 17054 22318 17106
rect 22370 17054 23044 17106
rect 21980 17052 23044 17054
rect 21420 17042 21476 17052
rect 21868 16996 21924 17006
rect 21756 16994 21924 16996
rect 21756 16942 21870 16994
rect 21922 16942 21924 16994
rect 21756 16940 21924 16942
rect 21644 16884 21700 16894
rect 21644 16790 21700 16828
rect 21532 16772 21588 16782
rect 21532 16678 21588 16716
rect 21756 16210 21812 16940
rect 21868 16930 21924 16940
rect 21756 16158 21758 16210
rect 21810 16158 21812 16210
rect 21756 16146 21812 16158
rect 21308 16046 21310 16098
rect 21362 16046 21364 16098
rect 21308 16034 21364 16046
rect 21532 16100 21588 16110
rect 21532 16006 21588 16044
rect 21756 15988 21812 15998
rect 21980 15988 22036 17052
rect 22316 17042 22372 17052
rect 22540 16882 22596 16894
rect 22540 16830 22542 16882
rect 22594 16830 22596 16882
rect 22540 16212 22596 16830
rect 22596 16156 22708 16212
rect 22540 16146 22596 16156
rect 21756 15986 22036 15988
rect 21756 15934 21758 15986
rect 21810 15934 22036 15986
rect 21756 15932 22036 15934
rect 22540 15988 22596 15998
rect 21756 15922 21812 15932
rect 22540 15894 22596 15932
rect 21196 15486 21198 15538
rect 21250 15486 21252 15538
rect 21196 15474 21252 15486
rect 22204 15876 22260 15886
rect 21084 15026 21140 15036
rect 21644 15314 21700 15326
rect 21644 15262 21646 15314
rect 21698 15262 21700 15314
rect 21644 15092 21700 15262
rect 22204 15204 22260 15820
rect 22316 15316 22372 15326
rect 22316 15222 22372 15260
rect 22204 15138 22260 15148
rect 21644 14420 21700 15036
rect 21644 14354 21700 14364
rect 22652 13972 22708 16156
rect 23100 16098 23156 19740
rect 23212 19234 23268 20636
rect 23324 20018 23380 21308
rect 23324 19966 23326 20018
rect 23378 19966 23380 20018
rect 23324 19954 23380 19966
rect 23436 21140 23492 21150
rect 23436 20018 23492 21084
rect 23436 19966 23438 20018
rect 23490 19966 23492 20018
rect 23436 19908 23492 19966
rect 23436 19572 23492 19852
rect 23436 19506 23492 19516
rect 23548 19348 23604 21756
rect 23660 20132 23716 20142
rect 23660 19906 23716 20076
rect 23772 20130 23828 22428
rect 23996 22428 24220 22484
rect 23884 22260 23940 22270
rect 23884 22166 23940 22204
rect 23996 21588 24052 22428
rect 24220 22418 24276 22428
rect 23772 20078 23774 20130
rect 23826 20078 23828 20130
rect 23772 20066 23828 20078
rect 23884 20804 23940 20814
rect 23996 20804 24052 21532
rect 24556 21588 24612 26852
rect 24668 26290 24724 27020
rect 24668 26238 24670 26290
rect 24722 26238 24724 26290
rect 24668 26226 24724 26238
rect 24780 25732 24836 25742
rect 24780 25506 24836 25676
rect 24780 25454 24782 25506
rect 24834 25454 24836 25506
rect 24780 25442 24836 25454
rect 24780 23940 24836 23950
rect 24668 23044 24724 23054
rect 24780 23044 24836 23884
rect 24668 23042 24836 23044
rect 24668 22990 24670 23042
rect 24722 22990 24836 23042
rect 24668 22988 24836 22990
rect 24668 22978 24724 22988
rect 24668 22484 24724 22494
rect 24668 22370 24724 22428
rect 24668 22318 24670 22370
rect 24722 22318 24724 22370
rect 24668 22306 24724 22318
rect 24780 21924 24836 22988
rect 24892 21924 24948 21934
rect 24780 21868 24892 21924
rect 24892 21858 24948 21868
rect 24556 21474 24612 21532
rect 24556 21422 24558 21474
rect 24610 21422 24612 21474
rect 24556 21410 24612 21422
rect 24556 20916 24612 20926
rect 24556 20822 24612 20860
rect 23884 20802 24052 20804
rect 23884 20750 23886 20802
rect 23938 20750 24052 20802
rect 23884 20748 24052 20750
rect 23660 19854 23662 19906
rect 23714 19854 23716 19906
rect 23660 19842 23716 19854
rect 23884 20020 23940 20748
rect 23996 20244 24052 20282
rect 23996 20178 24052 20188
rect 25004 20188 25060 29484
rect 25228 29428 25284 29438
rect 25228 29334 25284 29372
rect 25452 28868 25508 28878
rect 25564 28868 25620 29484
rect 25508 28812 25620 28868
rect 25452 28802 25508 28812
rect 25340 28644 25396 28654
rect 25340 27970 25396 28588
rect 25788 28532 25844 31836
rect 25900 32338 26516 32340
rect 25900 32286 26462 32338
rect 26514 32286 26516 32338
rect 25900 32284 26516 32286
rect 25900 31106 25956 32284
rect 26460 32274 26516 32284
rect 25900 31054 25902 31106
rect 25954 31054 25956 31106
rect 25900 31042 25956 31054
rect 26124 31220 26180 31230
rect 26572 31220 26628 33292
rect 26684 33292 26964 33348
rect 27244 34132 27300 34142
rect 27244 33346 27300 34076
rect 27244 33294 27246 33346
rect 27298 33294 27300 33346
rect 26684 32452 26740 33292
rect 27244 33282 27300 33294
rect 27356 33346 27412 34636
rect 27356 33294 27358 33346
rect 27410 33294 27412 33346
rect 27356 33282 27412 33294
rect 27580 33572 27636 35308
rect 28364 34916 28420 35308
rect 29260 35364 29316 35534
rect 29708 35586 29764 35598
rect 29708 35534 29710 35586
rect 29762 35534 29764 35586
rect 29260 35298 29316 35308
rect 29372 35474 29428 35486
rect 29372 35422 29374 35474
rect 29426 35422 29428 35474
rect 29148 35252 29204 35262
rect 28140 34914 28420 34916
rect 28140 34862 28366 34914
rect 28418 34862 28420 34914
rect 28140 34860 28420 34862
rect 27692 34804 27748 34814
rect 28028 34804 28084 34814
rect 27692 34802 28084 34804
rect 27692 34750 27694 34802
rect 27746 34750 28030 34802
rect 28082 34750 28084 34802
rect 27692 34748 28084 34750
rect 27692 34738 27748 34748
rect 28028 34356 28084 34748
rect 27580 33346 27636 33516
rect 27580 33294 27582 33346
rect 27634 33294 27636 33346
rect 26796 33124 26852 33134
rect 26796 33030 26852 33068
rect 27468 32788 27524 32798
rect 27020 32786 27524 32788
rect 27020 32734 27470 32786
rect 27522 32734 27524 32786
rect 27020 32732 27524 32734
rect 26908 32676 26964 32686
rect 26908 32582 26964 32620
rect 27020 32674 27076 32732
rect 27468 32722 27524 32732
rect 27020 32622 27022 32674
rect 27074 32622 27076 32674
rect 27020 32610 27076 32622
rect 27132 32564 27188 32574
rect 26684 32396 26964 32452
rect 26684 31220 26740 31230
rect 25788 28530 26068 28532
rect 25788 28478 25790 28530
rect 25842 28478 26068 28530
rect 25788 28476 26068 28478
rect 25788 28466 25844 28476
rect 26012 28082 26068 28476
rect 26012 28030 26014 28082
rect 26066 28030 26068 28082
rect 26012 28018 26068 28030
rect 25340 27918 25342 27970
rect 25394 27918 25396 27970
rect 25340 27906 25396 27918
rect 25228 27748 25284 27758
rect 25228 27654 25284 27692
rect 25452 27748 25508 27758
rect 25452 26908 25508 27692
rect 26124 27524 26180 31164
rect 26348 31218 26740 31220
rect 26348 31166 26686 31218
rect 26738 31166 26740 31218
rect 26348 31164 26740 31166
rect 26236 30212 26292 30222
rect 26236 30118 26292 30156
rect 26348 28756 26404 31164
rect 26684 31154 26740 31164
rect 26908 30212 26964 32396
rect 27132 31220 27188 32508
rect 27244 32564 27300 32574
rect 27580 32564 27636 33294
rect 27804 34132 27860 34142
rect 27244 32562 27636 32564
rect 27244 32510 27246 32562
rect 27298 32510 27636 32562
rect 27244 32508 27636 32510
rect 27692 32674 27748 32686
rect 27692 32622 27694 32674
rect 27746 32622 27748 32674
rect 27244 32498 27300 32508
rect 27468 32004 27524 32014
rect 27468 31890 27524 31948
rect 27468 31838 27470 31890
rect 27522 31838 27524 31890
rect 27468 31826 27524 31838
rect 27692 31668 27748 32622
rect 27804 32674 27860 34076
rect 28028 33348 28084 34300
rect 28140 34018 28196 34860
rect 28364 34850 28420 34860
rect 28700 35140 28756 35150
rect 28588 34356 28644 34366
rect 28588 34262 28644 34300
rect 28700 34242 28756 35084
rect 29148 34804 29204 35196
rect 28700 34190 28702 34242
rect 28754 34190 28756 34242
rect 28364 34132 28420 34142
rect 28700 34132 28756 34190
rect 28364 34038 28420 34076
rect 28476 34076 28756 34132
rect 28812 34802 29204 34804
rect 28812 34750 29150 34802
rect 29202 34750 29204 34802
rect 28812 34748 29204 34750
rect 28140 33966 28142 34018
rect 28194 33966 28196 34018
rect 28140 33954 28196 33966
rect 28252 33572 28308 33582
rect 28252 33570 28420 33572
rect 28252 33518 28254 33570
rect 28306 33518 28420 33570
rect 28252 33516 28420 33518
rect 28252 33506 28308 33516
rect 28140 33348 28196 33358
rect 28028 33346 28308 33348
rect 28028 33294 28142 33346
rect 28194 33294 28308 33346
rect 28028 33292 28308 33294
rect 28140 33282 28196 33292
rect 27916 33122 27972 33134
rect 27916 33070 27918 33122
rect 27970 33070 27972 33122
rect 27916 32788 27972 33070
rect 27972 32732 28084 32788
rect 27916 32722 27972 32732
rect 27804 32622 27806 32674
rect 27858 32622 27860 32674
rect 27804 32610 27860 32622
rect 28028 32004 28084 32732
rect 28252 32674 28308 33292
rect 28252 32622 28254 32674
rect 28306 32622 28308 32674
rect 28252 32610 28308 32622
rect 28364 32676 28420 33516
rect 28476 33346 28532 34076
rect 28476 33294 28478 33346
rect 28530 33294 28532 33346
rect 28476 33282 28532 33294
rect 28700 32788 28756 32798
rect 28700 32694 28756 32732
rect 28028 31890 28084 31948
rect 28028 31838 28030 31890
rect 28082 31838 28084 31890
rect 28028 31826 28084 31838
rect 27916 31668 27972 31678
rect 27692 31612 27916 31668
rect 27916 31574 27972 31612
rect 27132 31218 27524 31220
rect 27132 31166 27134 31218
rect 27186 31166 27524 31218
rect 27132 31164 27524 31166
rect 27132 31154 27188 31164
rect 27468 30324 27524 31164
rect 27692 30882 27748 30894
rect 28140 30884 28196 30894
rect 27692 30830 27694 30882
rect 27746 30830 27748 30882
rect 27692 30436 27748 30830
rect 27692 30370 27748 30380
rect 27804 30882 28196 30884
rect 27804 30830 28142 30882
rect 28194 30830 28196 30882
rect 27804 30828 28196 30830
rect 27468 30258 27524 30268
rect 27356 30212 27412 30222
rect 26908 30156 27356 30212
rect 27356 30118 27412 30156
rect 27692 30212 27748 30222
rect 27804 30212 27860 30828
rect 28140 30818 28196 30828
rect 28140 30436 28196 30446
rect 28140 30342 28196 30380
rect 27692 30210 27860 30212
rect 27692 30158 27694 30210
rect 27746 30158 27860 30210
rect 27692 30156 27860 30158
rect 27916 30210 27972 30222
rect 27916 30158 27918 30210
rect 27970 30158 27972 30210
rect 26796 30100 26852 30110
rect 26796 30098 26964 30100
rect 26796 30046 26798 30098
rect 26850 30046 26964 30098
rect 26796 30044 26964 30046
rect 26796 30034 26852 30044
rect 26348 28642 26404 28700
rect 26348 28590 26350 28642
rect 26402 28590 26404 28642
rect 26348 28578 26404 28590
rect 26460 29986 26516 29998
rect 26460 29934 26462 29986
rect 26514 29934 26516 29986
rect 26348 27858 26404 27870
rect 26348 27806 26350 27858
rect 26402 27806 26404 27858
rect 26348 27636 26404 27806
rect 26348 27570 26404 27580
rect 25340 26852 25508 26908
rect 25900 27468 26180 27524
rect 25228 26178 25284 26190
rect 25228 26126 25230 26178
rect 25282 26126 25284 26178
rect 25228 25956 25284 26126
rect 25228 25890 25284 25900
rect 25116 25508 25172 25518
rect 25116 25394 25172 25452
rect 25116 25342 25118 25394
rect 25170 25342 25172 25394
rect 25116 25330 25172 25342
rect 25228 24724 25284 24734
rect 25228 24630 25284 24668
rect 25340 23380 25396 26852
rect 25452 26292 25508 26302
rect 25452 25506 25508 26236
rect 25452 25454 25454 25506
rect 25506 25454 25508 25506
rect 25452 25442 25508 25454
rect 25788 26180 25844 26190
rect 25228 23378 25396 23380
rect 25228 23326 25342 23378
rect 25394 23326 25396 23378
rect 25228 23324 25396 23326
rect 25228 21588 25284 23324
rect 25340 23314 25396 23324
rect 25452 23938 25508 23950
rect 25452 23886 25454 23938
rect 25506 23886 25508 23938
rect 25340 22484 25396 22494
rect 25340 22370 25396 22428
rect 25340 22318 25342 22370
rect 25394 22318 25396 22370
rect 25340 22306 25396 22318
rect 25340 21588 25396 21598
rect 25228 21586 25396 21588
rect 25228 21534 25342 21586
rect 25394 21534 25396 21586
rect 25228 21532 25396 21534
rect 25228 20580 25284 20590
rect 24220 20132 24276 20142
rect 23548 19292 23828 19348
rect 23212 19182 23214 19234
rect 23266 19182 23268 19234
rect 23212 19170 23268 19182
rect 23548 19124 23604 19134
rect 23660 19124 23716 19134
rect 23604 19122 23716 19124
rect 23604 19070 23662 19122
rect 23714 19070 23716 19122
rect 23604 19068 23716 19070
rect 23436 18340 23492 18350
rect 23324 18338 23492 18340
rect 23324 18286 23438 18338
rect 23490 18286 23492 18338
rect 23324 18284 23492 18286
rect 23212 18004 23268 18014
rect 23212 17666 23268 17948
rect 23324 17780 23380 18284
rect 23436 18274 23492 18284
rect 23548 18116 23604 19068
rect 23660 19058 23716 19068
rect 23324 17714 23380 17724
rect 23436 18060 23604 18116
rect 23660 18788 23716 18798
rect 23212 17614 23214 17666
rect 23266 17614 23268 17666
rect 23212 17602 23268 17614
rect 23436 17556 23492 18060
rect 23436 17462 23492 17500
rect 23436 17108 23492 17118
rect 23660 17108 23716 18732
rect 23436 17106 23716 17108
rect 23436 17054 23438 17106
rect 23490 17054 23716 17106
rect 23436 17052 23716 17054
rect 23436 17042 23492 17052
rect 23772 16996 23828 19292
rect 23884 18228 23940 19964
rect 24108 20076 24220 20132
rect 23996 19236 24052 19246
rect 24108 19236 24164 20076
rect 24220 20066 24276 20076
rect 24332 20130 24388 20142
rect 24332 20078 24334 20130
rect 24386 20078 24388 20130
rect 24332 19348 24388 20078
rect 24668 20132 24724 20142
rect 25004 20132 25172 20188
rect 24668 20038 24724 20076
rect 24332 19282 24388 19292
rect 25004 19460 25060 19470
rect 25004 19346 25060 19404
rect 25004 19294 25006 19346
rect 25058 19294 25060 19346
rect 25004 19282 25060 19294
rect 23996 19234 24164 19236
rect 23996 19182 23998 19234
rect 24050 19182 24164 19234
rect 23996 19180 24164 19182
rect 23996 19170 24052 19180
rect 24444 19012 24500 19022
rect 24444 18918 24500 18956
rect 24332 18900 24388 18910
rect 24220 18450 24276 18462
rect 24220 18398 24222 18450
rect 24274 18398 24276 18450
rect 24220 18228 24276 18398
rect 23884 18172 24220 18228
rect 23884 17892 23940 17902
rect 23884 17106 23940 17836
rect 24108 17668 24164 18172
rect 24220 18162 24276 18172
rect 23884 17054 23886 17106
rect 23938 17054 23940 17106
rect 23884 17042 23940 17054
rect 23996 17666 24164 17668
rect 23996 17614 24110 17666
rect 24162 17614 24164 17666
rect 23996 17612 24164 17614
rect 23100 16046 23102 16098
rect 23154 16046 23156 16098
rect 23100 14196 23156 16046
rect 23548 16940 23828 16996
rect 23548 16210 23604 16940
rect 23548 16158 23550 16210
rect 23602 16158 23604 16210
rect 23548 15988 23604 16158
rect 23996 16098 24052 17612
rect 24108 17602 24164 17612
rect 24332 17106 24388 18844
rect 24668 18340 24724 18350
rect 24556 18338 24724 18340
rect 24556 18286 24670 18338
rect 24722 18286 24724 18338
rect 24556 18284 24724 18286
rect 24556 18004 24612 18284
rect 24668 18274 24724 18284
rect 24332 17054 24334 17106
rect 24386 17054 24388 17106
rect 24332 17042 24388 17054
rect 24444 17108 24500 17118
rect 24556 17108 24612 17948
rect 24892 17780 24948 17790
rect 24780 17668 24836 17678
rect 24780 17574 24836 17612
rect 24500 17052 24612 17108
rect 24668 17108 24724 17118
rect 24444 17042 24500 17052
rect 24668 16210 24724 17052
rect 24780 17108 24836 17118
rect 24892 17108 24948 17724
rect 24780 17106 24948 17108
rect 24780 17054 24782 17106
rect 24834 17054 24948 17106
rect 24780 17052 24948 17054
rect 24780 17042 24836 17052
rect 24668 16158 24670 16210
rect 24722 16158 24724 16210
rect 24668 16146 24724 16158
rect 23996 16046 23998 16098
rect 24050 16046 24052 16098
rect 23996 16034 24052 16046
rect 24556 16100 24612 16110
rect 23548 15922 23604 15932
rect 24556 15538 24612 16044
rect 24556 15486 24558 15538
rect 24610 15486 24612 15538
rect 24556 15474 24612 15486
rect 23660 14420 23716 14430
rect 23100 14140 23492 14196
rect 21196 13636 21252 13646
rect 21756 13636 21812 13646
rect 21196 13634 21700 13636
rect 21196 13582 21198 13634
rect 21250 13582 21700 13634
rect 21196 13580 21700 13582
rect 21196 13570 21252 13580
rect 21084 13300 21140 13310
rect 21084 12516 21140 13244
rect 21644 13186 21700 13580
rect 21644 13134 21646 13186
rect 21698 13134 21700 13186
rect 21644 13122 21700 13134
rect 21644 12962 21700 12974
rect 21644 12910 21646 12962
rect 21698 12910 21700 12962
rect 21644 12740 21700 12910
rect 21644 12674 21700 12684
rect 21084 12402 21140 12460
rect 21084 12350 21086 12402
rect 21138 12350 21140 12402
rect 21084 12338 21140 12350
rect 20860 11666 20916 11676
rect 21420 12290 21476 12302
rect 21420 12238 21422 12290
rect 21474 12238 21476 12290
rect 20412 11342 20414 11394
rect 20466 11342 20468 11394
rect 20412 11330 20468 11342
rect 20860 11284 20916 11294
rect 20860 11190 20916 11228
rect 20972 10836 21028 10846
rect 20524 10500 20580 10510
rect 20300 10498 20580 10500
rect 20300 10446 20526 10498
rect 20578 10446 20580 10498
rect 20300 10444 20580 10446
rect 20524 10434 20580 10444
rect 20300 10052 20356 10062
rect 20300 9958 20356 9996
rect 19740 9940 19796 9950
rect 20076 9940 20132 9950
rect 19516 9650 19572 9660
rect 19628 9938 20132 9940
rect 19628 9886 19742 9938
rect 19794 9886 20078 9938
rect 20130 9886 20132 9938
rect 19628 9884 20132 9886
rect 18844 9214 18846 9266
rect 18898 9214 18900 9266
rect 18844 9202 18900 9214
rect 19068 9268 19124 9278
rect 19628 9268 19684 9884
rect 19740 9874 19796 9884
rect 20076 9874 20132 9884
rect 20636 9604 20692 9614
rect 20636 9510 20692 9548
rect 20188 9492 20244 9502
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9268 20244 9436
rect 19068 9266 19684 9268
rect 19068 9214 19070 9266
rect 19122 9214 19684 9266
rect 19068 9212 19684 9214
rect 19964 9212 20244 9268
rect 19068 9202 19124 9212
rect 19516 9044 19572 9054
rect 19964 9044 20020 9212
rect 20636 9156 20692 9166
rect 20636 9062 20692 9100
rect 20524 9044 20580 9054
rect 19516 9042 20020 9044
rect 19516 8990 19518 9042
rect 19570 8990 20020 9042
rect 19516 8988 20020 8990
rect 20412 9042 20580 9044
rect 20412 8990 20526 9042
rect 20578 8990 20580 9042
rect 20412 8988 20580 8990
rect 19516 8978 19572 8988
rect 18956 8930 19012 8942
rect 18956 8878 18958 8930
rect 19010 8878 19012 8930
rect 18508 8820 18564 8830
rect 18956 8820 19012 8878
rect 20076 8932 20132 8942
rect 20076 8838 20132 8876
rect 18508 8818 19012 8820
rect 18508 8766 18510 8818
rect 18562 8766 19012 8818
rect 18508 8764 19012 8766
rect 20188 8818 20244 8830
rect 20188 8766 20190 8818
rect 20242 8766 20244 8818
rect 18508 8754 18564 8764
rect 18396 8540 19236 8596
rect 19068 8372 19124 8382
rect 18844 8370 19124 8372
rect 18844 8318 19070 8370
rect 19122 8318 19124 8370
rect 18844 8316 19124 8318
rect 17948 8148 18004 8158
rect 17388 6802 17556 6804
rect 17388 6750 17390 6802
rect 17442 6750 17556 6802
rect 17388 6748 17556 6750
rect 17724 7364 17780 7374
rect 17388 6738 17444 6748
rect 17724 6690 17780 7308
rect 17724 6638 17726 6690
rect 17778 6638 17780 6690
rect 17724 6356 17780 6638
rect 17724 6290 17780 6300
rect 17836 6580 17892 6590
rect 17724 6132 17780 6142
rect 17724 6038 17780 6076
rect 17836 6130 17892 6524
rect 17836 6078 17838 6130
rect 17890 6078 17892 6130
rect 17836 6066 17892 6078
rect 17948 6018 18004 8092
rect 18508 6580 18564 6618
rect 18508 6514 18564 6524
rect 17948 5966 17950 6018
rect 18002 5966 18004 6018
rect 17948 5954 18004 5966
rect 18508 6356 18564 6366
rect 17164 5730 17220 5740
rect 18508 5122 18564 6300
rect 18508 5070 18510 5122
rect 18562 5070 18564 5122
rect 18508 5058 18564 5070
rect 18620 5908 18676 5918
rect 18620 5124 18676 5852
rect 18844 5236 18900 8316
rect 19068 8306 19124 8316
rect 19180 7476 19236 8540
rect 20188 8372 20244 8766
rect 20188 8306 20244 8316
rect 19180 7410 19236 7420
rect 19404 8258 19460 8270
rect 19404 8206 19406 8258
rect 19458 8206 19460 8258
rect 18956 6020 19012 6030
rect 18956 5906 19012 5964
rect 19404 6020 19460 8206
rect 19852 8258 19908 8270
rect 19852 8206 19854 8258
rect 19906 8206 19908 8258
rect 19852 8036 19908 8206
rect 19852 7970 19908 7980
rect 20412 8036 20468 8988
rect 20524 8978 20580 8988
rect 20748 8932 20804 8942
rect 20636 8818 20692 8830
rect 20636 8766 20638 8818
rect 20690 8766 20692 8818
rect 20524 8596 20580 8606
rect 20524 8146 20580 8540
rect 20636 8260 20692 8766
rect 20748 8370 20804 8876
rect 20748 8318 20750 8370
rect 20802 8318 20804 8370
rect 20748 8306 20804 8318
rect 20636 8194 20692 8204
rect 20524 8094 20526 8146
rect 20578 8094 20580 8146
rect 20524 8082 20580 8094
rect 20412 7970 20468 7980
rect 20636 8036 20692 8046
rect 20636 8034 20804 8036
rect 20636 7982 20638 8034
rect 20690 7982 20804 8034
rect 20636 7980 20804 7982
rect 20636 7970 20692 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20636 6804 20692 6814
rect 20636 6710 20692 6748
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19404 5954 19460 5964
rect 19628 6018 19684 6030
rect 19628 5966 19630 6018
rect 19682 5966 19684 6018
rect 18956 5854 18958 5906
rect 19010 5854 19012 5906
rect 18956 5842 19012 5854
rect 19068 5794 19124 5806
rect 19068 5742 19070 5794
rect 19122 5742 19124 5794
rect 19068 5346 19124 5742
rect 19068 5294 19070 5346
rect 19122 5294 19124 5346
rect 19068 5282 19124 5294
rect 18956 5236 19012 5246
rect 18844 5234 19012 5236
rect 18844 5182 18958 5234
rect 19010 5182 19012 5234
rect 18844 5180 19012 5182
rect 18956 5170 19012 5180
rect 18620 5058 18676 5068
rect 17724 5012 17780 5022
rect 17052 3502 17054 3554
rect 17106 3502 17108 3554
rect 17052 3490 17108 3502
rect 17276 5010 17780 5012
rect 17276 4958 17726 5010
rect 17778 4958 17780 5010
rect 17276 4956 17780 4958
rect 17276 3442 17332 4956
rect 17724 4946 17780 4956
rect 17500 4340 17556 4350
rect 17500 4246 17556 4284
rect 17276 3390 17278 3442
rect 17330 3390 17332 3442
rect 17276 3378 17332 3390
rect 17500 4116 17556 4126
rect 15372 3332 15428 3342
rect 15372 3330 15540 3332
rect 15372 3278 15374 3330
rect 15426 3278 15540 3330
rect 15372 3276 15540 3278
rect 15372 3266 15428 3276
rect 15484 800 15540 3276
rect 17500 980 17556 4060
rect 18508 4116 18564 4126
rect 18508 4022 18564 4060
rect 19628 3556 19684 5966
rect 20188 6020 20244 6030
rect 20076 5908 20132 5918
rect 20076 5814 20132 5852
rect 19740 5124 19796 5134
rect 19740 5030 19796 5068
rect 20188 5122 20244 5964
rect 20748 6018 20804 7980
rect 20972 7924 21028 10780
rect 21308 10612 21364 10622
rect 21308 10518 21364 10556
rect 21420 10164 21476 12238
rect 21756 12290 21812 13580
rect 22652 13076 22708 13916
rect 22428 13020 22708 13076
rect 22764 13748 22820 13758
rect 21980 12852 22036 12862
rect 21980 12758 22036 12796
rect 22428 12402 22484 13020
rect 22764 12964 22820 13692
rect 23324 13636 23380 13646
rect 22540 12908 22764 12964
rect 22540 12850 22596 12908
rect 22764 12898 22820 12908
rect 22988 13634 23380 13636
rect 22988 13582 23326 13634
rect 23378 13582 23380 13634
rect 22988 13580 23380 13582
rect 22988 12962 23044 13580
rect 22988 12910 22990 12962
rect 23042 12910 23044 12962
rect 22988 12898 23044 12910
rect 22540 12798 22542 12850
rect 22594 12798 22596 12850
rect 22540 12786 22596 12798
rect 22876 12852 22932 12862
rect 22876 12758 22932 12796
rect 23212 12852 23268 12862
rect 22428 12350 22430 12402
rect 22482 12350 22484 12402
rect 22428 12338 22484 12350
rect 22652 12740 22708 12750
rect 22652 12404 22708 12684
rect 22764 12738 22820 12750
rect 22764 12686 22766 12738
rect 22818 12686 22820 12738
rect 22764 12628 22820 12686
rect 23212 12738 23268 12796
rect 23212 12686 23214 12738
rect 23266 12686 23268 12738
rect 23100 12628 23156 12638
rect 22764 12572 23100 12628
rect 22764 12404 22820 12414
rect 22652 12402 22820 12404
rect 22652 12350 22766 12402
rect 22818 12350 22820 12402
rect 22652 12348 22820 12350
rect 22764 12338 22820 12348
rect 21756 12238 21758 12290
rect 21810 12238 21812 12290
rect 21756 12226 21812 12238
rect 22092 12290 22148 12302
rect 22092 12238 22094 12290
rect 22146 12238 22148 12290
rect 22092 11844 22148 12238
rect 23100 12178 23156 12572
rect 23100 12126 23102 12178
rect 23154 12126 23156 12178
rect 23100 12114 23156 12126
rect 21644 11284 21700 11294
rect 21644 11190 21700 11228
rect 21980 11170 22036 11182
rect 21980 11118 21982 11170
rect 22034 11118 22036 11170
rect 21980 11060 22036 11118
rect 21980 10994 22036 11004
rect 22092 10948 22148 11788
rect 22428 12068 22484 12078
rect 22428 11508 22484 12012
rect 22428 11506 22596 11508
rect 22428 11454 22430 11506
rect 22482 11454 22596 11506
rect 22428 11452 22596 11454
rect 22428 11442 22484 11452
rect 22092 10892 22484 10948
rect 22092 10500 22148 10510
rect 21308 10108 21476 10164
rect 21756 10498 22148 10500
rect 21756 10446 22094 10498
rect 22146 10446 22148 10498
rect 21756 10444 22148 10446
rect 21308 9268 21364 10108
rect 21756 9938 21812 10444
rect 22092 10434 22148 10444
rect 21756 9886 21758 9938
rect 21810 9886 21812 9938
rect 21756 9874 21812 9886
rect 21644 9826 21700 9838
rect 21644 9774 21646 9826
rect 21698 9774 21700 9826
rect 21644 9716 21700 9774
rect 21980 9828 22036 9838
rect 21980 9734 22036 9772
rect 21644 9650 21700 9660
rect 22428 9602 22484 10892
rect 22428 9550 22430 9602
rect 22482 9550 22484 9602
rect 22428 9492 22484 9550
rect 22428 9426 22484 9436
rect 21308 9202 21364 9212
rect 22316 9268 22372 9278
rect 22540 9268 22596 11452
rect 22988 11284 23044 11294
rect 22988 11170 23044 11228
rect 22988 11118 22990 11170
rect 23042 11118 23044 11170
rect 22652 9828 22708 9838
rect 22876 9828 22932 9838
rect 22708 9772 22820 9828
rect 22652 9762 22708 9772
rect 22764 9714 22820 9772
rect 22876 9734 22932 9772
rect 22764 9662 22766 9714
rect 22818 9662 22820 9714
rect 22764 9650 22820 9662
rect 22652 9604 22708 9614
rect 22652 9510 22708 9548
rect 22316 9174 22372 9212
rect 22428 9212 22596 9268
rect 22876 9380 22932 9390
rect 22988 9380 23044 11118
rect 23212 10948 23268 12686
rect 23324 12178 23380 13580
rect 23324 12126 23326 12178
rect 23378 12126 23380 12178
rect 23324 12114 23380 12126
rect 23324 11732 23380 11742
rect 23324 11506 23380 11676
rect 23324 11454 23326 11506
rect 23378 11454 23380 11506
rect 23324 11442 23380 11454
rect 23212 10892 23380 10948
rect 23212 9716 23268 9726
rect 23212 9622 23268 9660
rect 22932 9324 23044 9380
rect 21420 9154 21476 9166
rect 21420 9102 21422 9154
rect 21474 9102 21476 9154
rect 21420 8596 21476 9102
rect 21420 8530 21476 8540
rect 21644 9042 21700 9054
rect 21644 8990 21646 9042
rect 21698 8990 21700 9042
rect 21420 8260 21476 8270
rect 21420 8166 21476 8204
rect 21308 8148 21364 8158
rect 21308 8054 21364 8092
rect 21644 8036 21700 8990
rect 21980 8708 22036 8718
rect 21644 7970 21700 7980
rect 21756 8258 21812 8270
rect 21756 8206 21758 8258
rect 21810 8206 21812 8258
rect 20972 6580 21028 7868
rect 21756 7588 21812 8206
rect 21756 6804 21812 7532
rect 21756 6738 21812 6748
rect 20972 6514 21028 6524
rect 21420 6690 21476 6702
rect 21420 6638 21422 6690
rect 21474 6638 21476 6690
rect 20748 5966 20750 6018
rect 20802 5966 20804 6018
rect 20748 5954 20804 5966
rect 21420 6020 21476 6638
rect 21868 6690 21924 6702
rect 21868 6638 21870 6690
rect 21922 6638 21924 6690
rect 21420 5954 21476 5964
rect 21756 6578 21812 6590
rect 21756 6526 21758 6578
rect 21810 6526 21812 6578
rect 20188 5070 20190 5122
rect 20242 5070 20244 5122
rect 20188 5058 20244 5070
rect 20412 5234 20468 5246
rect 20412 5182 20414 5234
rect 20466 5182 20468 5234
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20412 4562 20468 5182
rect 21532 5236 21588 5246
rect 21308 5124 21364 5134
rect 20748 5122 21364 5124
rect 20748 5070 21310 5122
rect 21362 5070 21364 5122
rect 20748 5068 21364 5070
rect 20748 5010 20804 5068
rect 21308 5058 21364 5068
rect 20748 4958 20750 5010
rect 20802 4958 20804 5010
rect 20748 4946 20804 4958
rect 20412 4510 20414 4562
rect 20466 4510 20468 4562
rect 20412 4498 20468 4510
rect 21196 4340 21252 4350
rect 20524 4228 20580 4238
rect 20524 4226 20916 4228
rect 20524 4174 20526 4226
rect 20578 4174 20916 4226
rect 20524 4172 20916 4174
rect 20524 4162 20580 4172
rect 20860 3666 20916 4172
rect 21196 4226 21252 4284
rect 21196 4174 21198 4226
rect 21250 4174 21252 4226
rect 21196 4162 21252 4174
rect 20860 3614 20862 3666
rect 20914 3614 20916 3666
rect 20860 3602 20916 3614
rect 19740 3556 19796 3566
rect 19628 3554 19796 3556
rect 19628 3502 19742 3554
rect 19794 3502 19796 3554
rect 19628 3500 19796 3502
rect 19740 3490 19796 3500
rect 19180 3332 19236 3342
rect 17276 924 17556 980
rect 19068 3330 19236 3332
rect 19068 3278 19182 3330
rect 19234 3278 19236 3330
rect 19068 3276 19236 3278
rect 17276 800 17332 924
rect 19068 800 19124 3276
rect 19180 3266 19236 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 924 21140 980
rect 20860 800 20916 924
rect 21084 868 21140 924
rect 21084 812 21252 868
rect 1120 0 1232 800
rect 2912 0 3024 800
rect 4704 0 4816 800
rect 6496 0 6608 800
rect 8288 0 8400 800
rect 10080 0 10192 800
rect 11872 0 11984 800
rect 13664 0 13776 800
rect 15456 0 15568 800
rect 17248 0 17360 800
rect 19040 0 19152 800
rect 20832 0 20944 800
rect 21196 756 21252 812
rect 21532 756 21588 5180
rect 21756 3556 21812 6526
rect 21868 4452 21924 6638
rect 21980 6356 22036 8652
rect 22428 8428 22484 9212
rect 22204 8372 22484 8428
rect 22540 9044 22596 9054
rect 22204 8148 22260 8372
rect 22204 7700 22260 8092
rect 22204 7634 22260 7644
rect 21980 5460 22036 6300
rect 21980 5394 22036 5404
rect 22428 6690 22484 6702
rect 22428 6638 22430 6690
rect 22482 6638 22484 6690
rect 22428 5684 22484 6638
rect 22316 5236 22372 5246
rect 22316 5142 22372 5180
rect 22428 5124 22484 5628
rect 22428 5058 22484 5068
rect 21868 4386 21924 4396
rect 21756 3490 21812 3500
rect 22540 2212 22596 8988
rect 22876 9042 22932 9324
rect 23324 9266 23380 10892
rect 23324 9214 23326 9266
rect 23378 9214 23380 9266
rect 23324 9202 23380 9214
rect 22876 8990 22878 9042
rect 22930 8990 22932 9042
rect 22652 8820 22708 8830
rect 22652 7700 22708 8764
rect 22876 8484 22932 8990
rect 22876 8418 22932 8428
rect 23212 9156 23268 9166
rect 23212 8484 23268 9100
rect 23324 8708 23380 8718
rect 23436 8708 23492 14140
rect 23660 12962 23716 14364
rect 23996 13972 24052 13982
rect 24332 13972 24388 13982
rect 24052 13970 24388 13972
rect 24052 13918 24334 13970
rect 24386 13918 24388 13970
rect 24052 13916 24388 13918
rect 23996 13878 24052 13916
rect 24332 13906 24388 13916
rect 24444 13972 24500 13982
rect 23772 13748 23828 13758
rect 23772 13654 23828 13692
rect 24444 13074 24500 13916
rect 24444 13022 24446 13074
rect 24498 13022 24500 13074
rect 24444 13010 24500 13022
rect 24668 13858 24724 13870
rect 24668 13806 24670 13858
rect 24722 13806 24724 13858
rect 23660 12910 23662 12962
rect 23714 12910 23716 12962
rect 23660 11396 23716 12910
rect 24668 12852 24724 13806
rect 24444 12628 24500 12638
rect 24444 12402 24500 12572
rect 24444 12350 24446 12402
rect 24498 12350 24500 12402
rect 24444 12338 24500 12350
rect 24668 12292 24724 12796
rect 24668 12226 24724 12236
rect 23996 12066 24052 12078
rect 23996 12014 23998 12066
rect 24050 12014 24052 12066
rect 23996 11732 24052 12014
rect 23996 11666 24052 11676
rect 24444 12066 24500 12078
rect 24444 12014 24446 12066
rect 24498 12014 24500 12066
rect 24444 11506 24500 12014
rect 24668 12068 24724 12078
rect 24668 11974 24724 12012
rect 24444 11454 24446 11506
rect 24498 11454 24500 11506
rect 24444 11442 24500 11454
rect 23548 11394 23716 11396
rect 23548 11342 23662 11394
rect 23714 11342 23716 11394
rect 23548 11340 23716 11342
rect 23548 10612 23604 11340
rect 23660 11330 23716 11340
rect 25116 10836 25172 20132
rect 25228 19124 25284 20524
rect 25340 19460 25396 21532
rect 25452 20188 25508 23886
rect 25676 23154 25732 23166
rect 25676 23102 25678 23154
rect 25730 23102 25732 23154
rect 25676 22484 25732 23102
rect 25676 22418 25732 22428
rect 25788 21812 25844 26124
rect 25900 25844 25956 27468
rect 26460 26908 26516 29934
rect 26908 29988 26964 30044
rect 26908 29922 26964 29932
rect 27132 29540 27188 29550
rect 26796 28530 26852 28542
rect 26796 28478 26798 28530
rect 26850 28478 26852 28530
rect 26572 28420 26628 28430
rect 26572 28082 26628 28364
rect 26572 28030 26574 28082
rect 26626 28030 26628 28082
rect 26572 28018 26628 28030
rect 26684 28084 26740 28094
rect 26796 28084 26852 28478
rect 26908 28420 26964 28430
rect 26908 28418 27076 28420
rect 26908 28366 26910 28418
rect 26962 28366 27076 28418
rect 26908 28364 27076 28366
rect 26908 28354 26964 28364
rect 26684 28082 26852 28084
rect 26684 28030 26686 28082
rect 26738 28030 26852 28082
rect 26684 28028 26852 28030
rect 26908 28084 26964 28094
rect 26684 28018 26740 28028
rect 26908 27990 26964 28028
rect 25900 25618 25956 25788
rect 25900 25566 25902 25618
rect 25954 25566 25956 25618
rect 25900 25554 25956 25566
rect 26124 26852 26516 26908
rect 26796 27858 26852 27870
rect 26796 27806 26798 27858
rect 26850 27806 26852 27858
rect 26796 26852 26852 27806
rect 27020 27186 27076 28364
rect 27020 27134 27022 27186
rect 27074 27134 27076 27186
rect 27020 27122 27076 27134
rect 27132 26908 27188 29484
rect 27692 29540 27748 30156
rect 27916 29876 27972 30158
rect 28364 30210 28420 32620
rect 28476 32562 28532 32574
rect 28476 32510 28478 32562
rect 28530 32510 28532 32562
rect 28476 32340 28532 32510
rect 28812 32450 28868 34748
rect 29148 34738 29204 34748
rect 29260 34690 29316 34702
rect 29260 34638 29262 34690
rect 29314 34638 29316 34690
rect 29260 34356 29316 34638
rect 29260 34290 29316 34300
rect 29260 34130 29316 34142
rect 29260 34078 29262 34130
rect 29314 34078 29316 34130
rect 29260 33348 29316 34078
rect 29260 33282 29316 33292
rect 29372 33346 29428 35422
rect 29708 35252 29764 35534
rect 29820 35476 29876 35486
rect 29820 35474 29988 35476
rect 29820 35422 29822 35474
rect 29874 35422 29988 35474
rect 29820 35420 29988 35422
rect 29820 35410 29876 35420
rect 29708 35186 29764 35196
rect 29932 35140 29988 35420
rect 29932 35074 29988 35084
rect 30156 35474 30212 35486
rect 30156 35422 30158 35474
rect 30210 35422 30212 35474
rect 29484 34916 29540 34926
rect 29484 34822 29540 34860
rect 30044 34916 30100 34954
rect 30044 34850 30100 34860
rect 29820 34802 29876 34814
rect 29820 34750 29822 34802
rect 29874 34750 29876 34802
rect 29820 34580 29876 34750
rect 29596 34524 29876 34580
rect 29484 34356 29540 34366
rect 29484 34262 29540 34300
rect 29484 34132 29540 34142
rect 29484 33458 29540 34076
rect 29596 34018 29652 34524
rect 29820 34356 29876 34366
rect 29596 33966 29598 34018
rect 29650 33966 29652 34018
rect 29596 33954 29652 33966
rect 29708 34130 29764 34142
rect 29708 34078 29710 34130
rect 29762 34078 29764 34130
rect 29484 33406 29486 33458
rect 29538 33406 29540 33458
rect 29484 33394 29540 33406
rect 29708 33460 29764 34078
rect 29708 33394 29764 33404
rect 29372 33294 29374 33346
rect 29426 33294 29428 33346
rect 29372 33282 29428 33294
rect 29596 33348 29652 33358
rect 29596 33254 29652 33292
rect 29820 33346 29876 34300
rect 30156 34356 30212 35422
rect 30268 35140 30324 35150
rect 30268 34356 30324 35084
rect 30380 35138 30436 36428
rect 30380 35086 30382 35138
rect 30434 35086 30436 35138
rect 30380 35074 30436 35086
rect 30380 34356 30436 34366
rect 30268 34354 30436 34356
rect 30268 34302 30382 34354
rect 30434 34302 30436 34354
rect 30268 34300 30436 34302
rect 30156 34290 30212 34300
rect 30380 34290 30436 34300
rect 30492 34356 30548 37100
rect 30716 37380 30772 37390
rect 30604 37042 30660 37054
rect 30604 36990 30606 37042
rect 30658 36990 30660 37042
rect 30604 36932 30660 36990
rect 30604 36866 30660 36876
rect 30492 34290 30548 34300
rect 30604 34244 30660 34254
rect 30604 34150 30660 34188
rect 29820 33294 29822 33346
rect 29874 33294 29876 33346
rect 29820 33282 29876 33294
rect 29932 34132 29988 34142
rect 29260 33122 29316 33134
rect 29260 33070 29262 33122
rect 29314 33070 29316 33122
rect 28924 32676 28980 32686
rect 29260 32676 29316 33070
rect 29372 32676 29428 32686
rect 28924 32562 28980 32620
rect 28924 32510 28926 32562
rect 28978 32510 28980 32562
rect 28924 32498 28980 32510
rect 29036 32674 29428 32676
rect 29036 32622 29374 32674
rect 29426 32622 29428 32674
rect 29036 32620 29428 32622
rect 28812 32398 28814 32450
rect 28866 32398 28868 32450
rect 28812 32386 28868 32398
rect 28476 32274 28532 32284
rect 28364 30158 28366 30210
rect 28418 30158 28420 30210
rect 28364 30146 28420 30158
rect 28476 31892 28532 31902
rect 28476 31554 28532 31836
rect 28476 31502 28478 31554
rect 28530 31502 28532 31554
rect 28476 30100 28532 31502
rect 28476 30034 28532 30044
rect 28588 30882 28644 30894
rect 28588 30830 28590 30882
rect 28642 30830 28644 30882
rect 27916 29810 27972 29820
rect 28140 29986 28196 29998
rect 28140 29934 28142 29986
rect 28194 29934 28196 29986
rect 27692 29474 27748 29484
rect 27468 29314 27524 29326
rect 27468 29262 27470 29314
rect 27522 29262 27524 29314
rect 27356 28530 27412 28542
rect 27356 28478 27358 28530
rect 27410 28478 27412 28530
rect 27356 27972 27412 28478
rect 27356 27906 27412 27916
rect 27468 27860 27524 29262
rect 27692 28644 27748 28654
rect 27692 28550 27748 28588
rect 27468 27766 27524 27804
rect 27580 28420 27636 28430
rect 27580 26964 27636 28364
rect 27804 28420 27860 28430
rect 27804 28326 27860 28364
rect 27916 28418 27972 28430
rect 27916 28366 27918 28418
rect 27970 28366 27972 28418
rect 27916 28084 27972 28366
rect 27132 26852 27524 26908
rect 26124 22484 26180 26852
rect 26796 26786 26852 26796
rect 27356 26180 27412 26190
rect 26796 26178 27412 26180
rect 26796 26126 27358 26178
rect 27410 26126 27412 26178
rect 26796 26124 27412 26126
rect 26796 25730 26852 26124
rect 27356 26114 27412 26124
rect 26796 25678 26798 25730
rect 26850 25678 26852 25730
rect 26796 25666 26852 25678
rect 27356 25956 27412 25966
rect 27356 25506 27412 25900
rect 27356 25454 27358 25506
rect 27410 25454 27412 25506
rect 27356 25442 27412 25454
rect 26684 25396 26740 25406
rect 26684 25302 26740 25340
rect 26460 25282 26516 25294
rect 26460 25230 26462 25282
rect 26514 25230 26516 25282
rect 26460 23940 26516 25230
rect 27468 24164 27524 26852
rect 27580 25506 27636 26908
rect 27692 28028 27916 28084
rect 27692 26068 27748 28028
rect 27916 28018 27972 28028
rect 28140 27970 28196 29934
rect 28588 29988 28644 30830
rect 28700 30772 28756 30782
rect 28700 30210 28756 30716
rect 28700 30158 28702 30210
rect 28754 30158 28756 30210
rect 28700 30146 28756 30158
rect 28588 28868 28644 29932
rect 28140 27918 28142 27970
rect 28194 27918 28196 27970
rect 28140 27906 28196 27918
rect 28364 28812 28644 28868
rect 27804 27074 27860 27086
rect 27804 27022 27806 27074
rect 27858 27022 27860 27074
rect 27804 26292 27860 27022
rect 28252 26852 28308 26862
rect 28252 26758 28308 26796
rect 28252 26404 28308 26414
rect 28140 26292 28196 26302
rect 27804 26290 28196 26292
rect 27804 26238 28142 26290
rect 28194 26238 28196 26290
rect 27804 26236 28196 26238
rect 28028 26068 28084 26078
rect 27692 26012 28028 26068
rect 27580 25454 27582 25506
rect 27634 25454 27636 25506
rect 27580 25442 27636 25454
rect 27804 25620 27860 25630
rect 27804 25506 27860 25564
rect 27804 25454 27806 25506
rect 27858 25454 27860 25506
rect 27804 25442 27860 25454
rect 28028 25506 28084 26012
rect 28028 25454 28030 25506
rect 28082 25454 28084 25506
rect 28028 25442 28084 25454
rect 28140 25508 28196 26236
rect 28140 25442 28196 25452
rect 27692 25396 27748 25406
rect 27692 25302 27748 25340
rect 27804 25284 27860 25294
rect 27860 25228 27972 25284
rect 27804 25218 27860 25228
rect 27356 24108 27524 24164
rect 27020 23940 27076 23950
rect 26460 23874 26516 23884
rect 26908 23884 27020 23940
rect 26908 23716 26964 23884
rect 27020 23874 27076 23884
rect 26348 23714 26964 23716
rect 26348 23662 26910 23714
rect 26962 23662 26964 23714
rect 26348 23660 26964 23662
rect 25900 22428 26180 22484
rect 26236 23604 26292 23614
rect 25900 21812 25956 22428
rect 26012 22260 26068 22270
rect 26012 22166 26068 22204
rect 25900 21756 26180 21812
rect 25788 21746 25844 21756
rect 25788 21586 25844 21598
rect 25788 21534 25790 21586
rect 25842 21534 25844 21586
rect 25788 21028 25844 21534
rect 26012 21586 26068 21598
rect 26012 21534 26014 21586
rect 26066 21534 26068 21586
rect 25788 20962 25844 20972
rect 25900 21474 25956 21486
rect 25900 21422 25902 21474
rect 25954 21422 25956 21474
rect 25900 20916 25956 21422
rect 25900 20850 25956 20860
rect 26012 20188 26068 21534
rect 26124 21476 26180 21756
rect 26124 20804 26180 21420
rect 26124 20738 26180 20748
rect 25452 20132 25620 20188
rect 25564 20018 25620 20132
rect 25564 19966 25566 20018
rect 25618 19966 25620 20018
rect 25340 19404 25508 19460
rect 25452 19348 25508 19404
rect 25452 19282 25508 19292
rect 25340 19124 25396 19134
rect 25228 19122 25396 19124
rect 25228 19070 25342 19122
rect 25394 19070 25396 19122
rect 25228 19068 25396 19070
rect 25340 19058 25396 19068
rect 25452 19124 25508 19134
rect 25340 18452 25396 18462
rect 25340 18358 25396 18396
rect 25228 18226 25284 18238
rect 25228 18174 25230 18226
rect 25282 18174 25284 18226
rect 25228 17668 25284 18174
rect 25228 17602 25284 17612
rect 25452 17106 25508 19068
rect 25452 17054 25454 17106
rect 25506 17054 25508 17106
rect 25452 17042 25508 17054
rect 25564 19012 25620 19966
rect 25676 20132 26068 20188
rect 26124 20580 26180 20590
rect 25676 19458 25732 20132
rect 25676 19406 25678 19458
rect 25730 19406 25732 19458
rect 25676 19394 25732 19406
rect 25900 19348 25956 19358
rect 25564 14530 25620 18956
rect 25788 19012 25844 19022
rect 25788 18450 25844 18956
rect 25788 18398 25790 18450
rect 25842 18398 25844 18450
rect 25788 18386 25844 18398
rect 25676 18226 25732 18238
rect 25676 18174 25678 18226
rect 25730 18174 25732 18226
rect 25676 17108 25732 18174
rect 25676 17042 25732 17052
rect 25788 16548 25844 16558
rect 25788 15538 25844 16492
rect 25788 15486 25790 15538
rect 25842 15486 25844 15538
rect 25788 15474 25844 15486
rect 25564 14478 25566 14530
rect 25618 14478 25620 14530
rect 25564 14466 25620 14478
rect 25900 14308 25956 19292
rect 26124 19234 26180 20524
rect 26236 20188 26292 23548
rect 26348 21810 26404 23660
rect 26908 23650 26964 23660
rect 27020 23714 27076 23726
rect 27020 23662 27022 23714
rect 27074 23662 27076 23714
rect 27020 23548 27076 23662
rect 27132 23716 27188 23726
rect 27132 23714 27300 23716
rect 27132 23662 27134 23714
rect 27186 23662 27300 23714
rect 27132 23660 27300 23662
rect 27132 23650 27188 23660
rect 26460 23492 27076 23548
rect 26460 23266 26516 23492
rect 26460 23214 26462 23266
rect 26514 23214 26516 23266
rect 26460 23202 26516 23214
rect 26348 21758 26350 21810
rect 26402 21758 26404 21810
rect 26348 21746 26404 21758
rect 26460 22260 26516 22270
rect 26460 21810 26516 22204
rect 27244 22036 27300 23660
rect 27356 22484 27412 24108
rect 27468 23940 27524 23950
rect 27692 23940 27748 23950
rect 27468 23938 27748 23940
rect 27468 23886 27470 23938
rect 27522 23886 27694 23938
rect 27746 23886 27748 23938
rect 27468 23884 27748 23886
rect 27468 23874 27524 23884
rect 27692 23874 27748 23884
rect 27356 22418 27412 22428
rect 27804 23714 27860 23726
rect 27804 23662 27806 23714
rect 27858 23662 27860 23714
rect 27804 23268 27860 23662
rect 27244 21980 27636 22036
rect 26460 21758 26462 21810
rect 26514 21758 26516 21810
rect 26460 21746 26516 21758
rect 27468 21812 27524 21822
rect 26572 21586 26628 21598
rect 26572 21534 26574 21586
rect 26626 21534 26628 21586
rect 26236 20132 26404 20188
rect 26124 19182 26126 19234
rect 26178 19182 26180 19234
rect 26012 19124 26068 19134
rect 26124 19124 26180 19182
rect 26236 19460 26292 19470
rect 26236 19234 26292 19404
rect 26236 19182 26238 19234
rect 26290 19182 26292 19234
rect 26236 19170 26292 19182
rect 26068 19068 26180 19124
rect 26012 19058 26068 19068
rect 26236 17220 26292 17230
rect 26236 17106 26292 17164
rect 26236 17054 26238 17106
rect 26290 17054 26292 17106
rect 26236 17042 26292 17054
rect 26348 16884 26404 20132
rect 26572 19348 26628 21534
rect 27020 21586 27076 21598
rect 27020 21534 27022 21586
rect 27074 21534 27076 21586
rect 26852 21476 26908 21486
rect 27020 21476 27076 21534
rect 26908 21420 26964 21476
rect 26852 21410 26964 21420
rect 27020 21410 27076 21420
rect 27132 21586 27188 21598
rect 27132 21534 27134 21586
rect 27186 21534 27188 21586
rect 26908 21140 26964 21410
rect 26908 21074 26964 21084
rect 26684 20914 26740 20926
rect 26684 20862 26686 20914
rect 26738 20862 26740 20914
rect 26684 20692 26740 20862
rect 27020 20692 27076 20702
rect 26684 20690 27076 20692
rect 26684 20638 27022 20690
rect 27074 20638 27076 20690
rect 26684 20636 27076 20638
rect 26684 20188 26740 20636
rect 27020 20626 27076 20636
rect 26684 20132 26852 20188
rect 26572 19292 26740 19348
rect 26460 19236 26516 19246
rect 26460 19142 26516 19180
rect 26460 18338 26516 18350
rect 26460 18286 26462 18338
rect 26514 18286 26516 18338
rect 26460 18004 26516 18286
rect 26572 18340 26628 18350
rect 26684 18340 26740 19292
rect 26796 19236 26852 20132
rect 27132 19908 27188 21534
rect 27468 21588 27524 21756
rect 27468 21522 27524 21532
rect 27356 21364 27412 21374
rect 27356 21270 27412 21308
rect 27356 21028 27412 21038
rect 27244 20804 27300 20814
rect 27244 20710 27300 20748
rect 27356 20578 27412 20972
rect 27580 20916 27636 21980
rect 27356 20526 27358 20578
rect 27410 20526 27412 20578
rect 27356 20514 27412 20526
rect 27468 20860 27636 20916
rect 27692 21700 27748 21710
rect 27804 21700 27860 23212
rect 27916 21810 27972 25228
rect 28028 23940 28084 23978
rect 28028 23874 28084 23884
rect 27916 21758 27918 21810
rect 27970 21758 27972 21810
rect 27916 21746 27972 21758
rect 28028 23716 28084 23726
rect 27692 21698 27860 21700
rect 27692 21646 27694 21698
rect 27746 21646 27860 21698
rect 27692 21644 27860 21646
rect 27132 19842 27188 19852
rect 27244 20356 27300 20366
rect 27244 19684 27300 20300
rect 27132 19628 27300 19684
rect 27356 19906 27412 19918
rect 27356 19854 27358 19906
rect 27410 19854 27412 19906
rect 26796 19142 26852 19180
rect 27020 19236 27076 19246
rect 27020 18676 27076 19180
rect 26628 18284 26740 18340
rect 26796 18620 27076 18676
rect 26572 18246 26628 18284
rect 26460 17938 26516 17948
rect 26572 16884 26628 16894
rect 26348 16882 26628 16884
rect 26348 16830 26574 16882
rect 26626 16830 26628 16882
rect 26348 16828 26628 16830
rect 26124 16324 26180 16334
rect 26124 15540 26180 16268
rect 26124 15446 26180 15484
rect 26348 14868 26404 16828
rect 26572 16818 26628 16828
rect 26684 16772 26740 16782
rect 26460 15988 26516 15998
rect 26460 15538 26516 15932
rect 26460 15486 26462 15538
rect 26514 15486 26516 15538
rect 26460 15474 26516 15486
rect 26684 15540 26740 16716
rect 26796 16210 26852 18620
rect 27020 18228 27076 18238
rect 26908 17778 26964 17790
rect 26908 17726 26910 17778
rect 26962 17726 26964 17778
rect 26908 17556 26964 17726
rect 26908 17490 26964 17500
rect 27020 16882 27076 18172
rect 27020 16830 27022 16882
rect 27074 16830 27076 16882
rect 27020 16818 27076 16830
rect 27132 16660 27188 19628
rect 27244 19236 27300 19246
rect 27244 19142 27300 19180
rect 27356 18450 27412 19854
rect 27356 18398 27358 18450
rect 27410 18398 27412 18450
rect 27356 18228 27412 18398
rect 27356 18162 27412 18172
rect 27468 17780 27524 20860
rect 27580 20692 27636 20702
rect 27580 20598 27636 20636
rect 27692 20244 27748 21644
rect 28028 21588 28084 23660
rect 28140 23492 28196 23502
rect 28140 22482 28196 23436
rect 28140 22430 28142 22482
rect 28194 22430 28196 22482
rect 28140 22418 28196 22430
rect 28252 21812 28308 26348
rect 28364 26292 28420 28812
rect 28588 28644 28644 28654
rect 28588 28550 28644 28588
rect 28476 28532 28532 28542
rect 28476 28438 28532 28476
rect 28700 28420 28756 28430
rect 28476 26964 28532 26974
rect 28476 26514 28532 26908
rect 28476 26462 28478 26514
rect 28530 26462 28532 26514
rect 28476 26450 28532 26462
rect 28588 26292 28644 26302
rect 28364 26236 28532 26292
rect 28364 23938 28420 23950
rect 28364 23886 28366 23938
rect 28418 23886 28420 23938
rect 28364 23828 28420 23886
rect 28364 23762 28420 23772
rect 28476 23716 28532 26236
rect 28588 25844 28644 26236
rect 28588 25778 28644 25788
rect 28588 25620 28644 25630
rect 28588 25282 28644 25564
rect 28588 25230 28590 25282
rect 28642 25230 28644 25282
rect 28588 24836 28644 25230
rect 28588 24770 28644 24780
rect 28476 23650 28532 23660
rect 28588 24500 28644 24510
rect 28588 23940 28644 24444
rect 28588 23042 28644 23884
rect 28588 22990 28590 23042
rect 28642 22990 28644 23042
rect 28588 22978 28644 22990
rect 27692 20178 27748 20188
rect 27804 21532 28084 21588
rect 28140 21756 28308 21812
rect 28476 22484 28532 22494
rect 27244 17724 27524 17780
rect 27580 18564 27636 18574
rect 27244 16772 27300 17724
rect 27580 17666 27636 18508
rect 27692 18452 27748 18462
rect 27692 17778 27748 18396
rect 27804 18004 27860 21532
rect 27916 21362 27972 21374
rect 27916 21310 27918 21362
rect 27970 21310 27972 21362
rect 27916 20692 27972 21310
rect 27916 20626 27972 20636
rect 28028 20916 28084 20926
rect 28028 20802 28084 20860
rect 28028 20750 28030 20802
rect 28082 20750 28084 20802
rect 27916 20356 27972 20366
rect 28028 20356 28084 20750
rect 27972 20300 28084 20356
rect 27916 20290 27972 20300
rect 28028 19460 28084 19470
rect 27804 17938 27860 17948
rect 27916 19234 27972 19246
rect 27916 19182 27918 19234
rect 27970 19182 27972 19234
rect 27692 17726 27694 17778
rect 27746 17726 27748 17778
rect 27692 17714 27748 17726
rect 27580 17614 27582 17666
rect 27634 17614 27636 17666
rect 27580 17602 27636 17614
rect 27356 17556 27412 17566
rect 27356 17462 27412 17500
rect 27804 17444 27860 17454
rect 27804 17350 27860 17388
rect 27692 16996 27748 17006
rect 27692 16902 27748 16940
rect 27244 16706 27300 16716
rect 26796 16158 26798 16210
rect 26850 16158 26852 16210
rect 26796 16146 26852 16158
rect 27020 16604 27188 16660
rect 26684 15538 26964 15540
rect 26684 15486 26686 15538
rect 26738 15486 26964 15538
rect 26684 15484 26964 15486
rect 26684 15474 26740 15484
rect 26348 14802 26404 14812
rect 26572 15202 26628 15214
rect 26572 15150 26574 15202
rect 26626 15150 26628 15202
rect 25340 14252 25956 14308
rect 25116 10770 25172 10780
rect 25228 11732 25284 11742
rect 23548 10546 23604 10556
rect 24220 10498 24276 10510
rect 24220 10446 24222 10498
rect 24274 10446 24276 10498
rect 23548 9826 23604 9838
rect 23548 9774 23550 9826
rect 23602 9774 23604 9826
rect 23548 9716 23604 9774
rect 23548 9650 23604 9660
rect 23772 9828 23828 9838
rect 24220 9828 24276 10446
rect 24668 10498 24724 10510
rect 24668 10446 24670 10498
rect 24722 10446 24724 10498
rect 24668 10164 24724 10446
rect 24668 10098 24724 10108
rect 23772 9826 24276 9828
rect 23772 9774 23774 9826
rect 23826 9774 24276 9826
rect 23772 9772 24276 9774
rect 23772 9604 23828 9772
rect 24444 9714 24500 9726
rect 24444 9662 24446 9714
rect 24498 9662 24500 9714
rect 24220 9604 24276 9614
rect 23772 9538 23828 9548
rect 23996 9602 24276 9604
rect 23996 9550 24222 9602
rect 24274 9550 24276 9602
rect 23996 9548 24276 9550
rect 23548 9042 23604 9054
rect 23548 8990 23550 9042
rect 23602 8990 23604 9042
rect 23548 8820 23604 8990
rect 23772 9044 23828 9054
rect 23996 9044 24052 9548
rect 24220 9538 24276 9548
rect 24332 9602 24388 9614
rect 24332 9550 24334 9602
rect 24386 9550 24388 9602
rect 23772 9042 24052 9044
rect 23772 8990 23774 9042
rect 23826 8990 24052 9042
rect 23772 8988 24052 8990
rect 24108 9380 24164 9390
rect 24108 9042 24164 9324
rect 24108 8990 24110 9042
rect 24162 8990 24164 9042
rect 23772 8978 23828 8988
rect 23660 8932 23716 8942
rect 23660 8838 23716 8876
rect 23548 8754 23604 8764
rect 23380 8652 23492 8708
rect 23324 8642 23380 8652
rect 23100 8260 23156 8270
rect 23100 8166 23156 8204
rect 22764 8146 22820 8158
rect 22764 8094 22766 8146
rect 22818 8094 22820 8146
rect 22764 7924 22820 8094
rect 22988 8148 23044 8158
rect 22764 7858 22820 7868
rect 22876 8034 22932 8046
rect 22876 7982 22878 8034
rect 22930 7982 22932 8034
rect 22876 7812 22932 7982
rect 22876 7746 22932 7756
rect 22652 7644 22820 7700
rect 22652 7476 22708 7486
rect 22652 6802 22708 7420
rect 22652 6750 22654 6802
rect 22706 6750 22708 6802
rect 22652 6738 22708 6750
rect 22764 5796 22820 7644
rect 22988 7474 23044 8092
rect 22988 7422 22990 7474
rect 23042 7422 23044 7474
rect 22988 7410 23044 7422
rect 23100 7700 23156 7710
rect 22988 6020 23044 6030
rect 22876 5796 22932 5806
rect 22764 5794 22932 5796
rect 22764 5742 22878 5794
rect 22930 5742 22932 5794
rect 22764 5740 22932 5742
rect 22876 5730 22932 5740
rect 22988 3666 23044 5964
rect 23100 4340 23156 7644
rect 23212 7586 23268 8428
rect 23772 8596 23828 8606
rect 23436 8258 23492 8270
rect 23436 8206 23438 8258
rect 23490 8206 23492 8258
rect 23212 7534 23214 7586
rect 23266 7534 23268 7586
rect 23212 7522 23268 7534
rect 23324 7588 23380 7598
rect 23324 7494 23380 7532
rect 23324 6802 23380 6814
rect 23324 6750 23326 6802
rect 23378 6750 23380 6802
rect 23324 6690 23380 6750
rect 23324 6638 23326 6690
rect 23378 6638 23380 6690
rect 23324 6626 23380 6638
rect 23436 6692 23492 8206
rect 23436 5908 23492 6636
rect 23772 7474 23828 8540
rect 23884 8148 23940 8988
rect 24108 8978 24164 8990
rect 24332 8708 24388 9550
rect 24444 9268 24500 9662
rect 24444 9202 24500 9212
rect 24780 9602 24836 9614
rect 24780 9550 24782 9602
rect 24834 9550 24836 9602
rect 24444 9042 24500 9054
rect 24444 8990 24446 9042
rect 24498 8990 24500 9042
rect 24444 8820 24500 8990
rect 24444 8754 24500 8764
rect 24556 9042 24612 9054
rect 24556 8990 24558 9042
rect 24610 8990 24612 9042
rect 24108 8652 24388 8708
rect 24108 8370 24164 8652
rect 24108 8318 24110 8370
rect 24162 8318 24164 8370
rect 24108 8306 24164 8318
rect 23884 8092 24500 8148
rect 24332 7812 24388 7822
rect 24332 7698 24388 7756
rect 24332 7646 24334 7698
rect 24386 7646 24388 7698
rect 24332 7634 24388 7646
rect 24444 7698 24500 8092
rect 24444 7646 24446 7698
rect 24498 7646 24500 7698
rect 24444 7634 24500 7646
rect 23772 7422 23774 7474
rect 23826 7422 23828 7474
rect 23660 6580 23716 6590
rect 23436 5842 23492 5852
rect 23548 6018 23604 6030
rect 23548 5966 23550 6018
rect 23602 5966 23604 6018
rect 23212 5794 23268 5806
rect 23212 5742 23214 5794
rect 23266 5742 23268 5794
rect 23212 5684 23268 5742
rect 23548 5796 23604 5966
rect 23660 5906 23716 6524
rect 23660 5854 23662 5906
rect 23714 5854 23716 5906
rect 23660 5842 23716 5854
rect 23548 5730 23604 5740
rect 23212 5618 23268 5628
rect 23772 5236 23828 7422
rect 24556 7476 24612 8990
rect 24668 9042 24724 9054
rect 24668 8990 24670 9042
rect 24722 8990 24724 9042
rect 24668 8596 24724 8990
rect 24780 9044 24836 9550
rect 25228 9268 25284 11676
rect 25340 11620 25396 14252
rect 26572 13972 26628 15150
rect 26908 14642 26964 15484
rect 26908 14590 26910 14642
rect 26962 14590 26964 14642
rect 26908 14578 26964 14590
rect 27020 14084 27076 16604
rect 27916 16436 27972 19182
rect 28028 18450 28084 19404
rect 28140 18900 28196 21756
rect 28252 21586 28308 21598
rect 28252 21534 28254 21586
rect 28306 21534 28308 21586
rect 28252 21364 28308 21534
rect 28476 21586 28532 22428
rect 28588 22146 28644 22158
rect 28588 22094 28590 22146
rect 28642 22094 28644 22146
rect 28588 21812 28644 22094
rect 28700 21812 28756 28364
rect 29036 26964 29092 32620
rect 29372 32610 29428 32620
rect 29708 32676 29764 32686
rect 29708 32582 29764 32620
rect 29820 32450 29876 32462
rect 29820 32398 29822 32450
rect 29874 32398 29876 32450
rect 29260 32340 29316 32350
rect 29260 32246 29316 32284
rect 29820 31780 29876 32398
rect 29932 31890 29988 34076
rect 30492 34018 30548 34030
rect 30492 33966 30494 34018
rect 30546 33966 30548 34018
rect 30380 33572 30436 33582
rect 30492 33572 30548 33966
rect 30380 33570 30548 33572
rect 30380 33518 30382 33570
rect 30434 33518 30548 33570
rect 30380 33516 30548 33518
rect 30716 33570 30772 37324
rect 30716 33518 30718 33570
rect 30770 33518 30772 33570
rect 30380 33506 30436 33516
rect 30716 33506 30772 33518
rect 29932 31838 29934 31890
rect 29986 31838 29988 31890
rect 29932 31826 29988 31838
rect 30156 33460 30212 33470
rect 30156 33346 30212 33404
rect 30156 33294 30158 33346
rect 30210 33294 30212 33346
rect 30156 31892 30212 33294
rect 30716 33012 30772 33022
rect 30716 32452 30772 32956
rect 30604 32450 30772 32452
rect 30604 32398 30718 32450
rect 30770 32398 30772 32450
rect 30604 32396 30772 32398
rect 30380 31892 30436 31902
rect 30156 31890 30436 31892
rect 30156 31838 30382 31890
rect 30434 31838 30436 31890
rect 30156 31836 30436 31838
rect 30380 31826 30436 31836
rect 29596 31724 29876 31780
rect 30044 31778 30100 31790
rect 30044 31726 30046 31778
rect 30098 31726 30100 31778
rect 29372 31668 29428 31678
rect 29372 31574 29428 31612
rect 29596 31554 29652 31724
rect 30044 31668 30100 31726
rect 30044 31602 30100 31612
rect 29596 31502 29598 31554
rect 29650 31502 29652 31554
rect 29148 30884 29204 30894
rect 29148 30790 29204 30828
rect 29596 30324 29652 31502
rect 29820 31556 29876 31566
rect 29708 30882 29764 30894
rect 29708 30830 29710 30882
rect 29762 30830 29764 30882
rect 29708 30436 29764 30830
rect 29820 30772 29876 31500
rect 30492 31108 30548 31118
rect 30044 30884 30100 30894
rect 30044 30882 30212 30884
rect 30044 30830 30046 30882
rect 30098 30830 30212 30882
rect 30044 30828 30212 30830
rect 30044 30818 30100 30828
rect 29932 30772 29988 30782
rect 29820 30716 29932 30772
rect 29932 30678 29988 30716
rect 29708 30380 29988 30436
rect 29596 30268 29876 30324
rect 29372 29986 29428 29998
rect 29372 29934 29374 29986
rect 29426 29934 29428 29986
rect 29148 29092 29204 29102
rect 29148 28754 29204 29036
rect 29148 28702 29150 28754
rect 29202 28702 29204 28754
rect 29148 27074 29204 28702
rect 29372 28420 29428 29934
rect 29708 29988 29764 29998
rect 29708 29894 29764 29932
rect 29372 28354 29428 28364
rect 29484 28532 29540 28542
rect 29484 27186 29540 28476
rect 29484 27134 29486 27186
rect 29538 27134 29540 27186
rect 29484 27122 29540 27134
rect 29148 27022 29150 27074
rect 29202 27022 29204 27074
rect 29148 27010 29204 27022
rect 28924 26908 29092 26964
rect 29372 26964 29428 27002
rect 28812 26292 28868 26302
rect 28812 25732 28868 26236
rect 28812 25666 28868 25676
rect 28812 24836 28868 24846
rect 28812 22260 28868 24780
rect 28924 23548 28980 26908
rect 29372 26898 29428 26908
rect 29596 26964 29652 27002
rect 29596 26898 29652 26908
rect 29708 26850 29764 26862
rect 29708 26798 29710 26850
rect 29762 26798 29764 26850
rect 29708 26516 29764 26798
rect 29372 26460 29764 26516
rect 29148 26404 29204 26414
rect 29372 26404 29428 26460
rect 29148 26402 29428 26404
rect 29148 26350 29150 26402
rect 29202 26350 29428 26402
rect 29148 26348 29428 26350
rect 29148 26068 29204 26348
rect 29148 26002 29204 26012
rect 29484 26290 29540 26302
rect 29484 26238 29486 26290
rect 29538 26238 29540 26290
rect 29372 25844 29428 25854
rect 29484 25844 29540 26238
rect 29428 25788 29540 25844
rect 29372 25778 29428 25788
rect 29820 25732 29876 30268
rect 29932 28756 29988 30380
rect 30156 29316 30212 30828
rect 30268 30212 30324 30222
rect 30268 29986 30324 30156
rect 30268 29934 30270 29986
rect 30322 29934 30324 29986
rect 30268 29540 30324 29934
rect 30492 29988 30548 31052
rect 30492 29922 30548 29932
rect 30268 29474 30324 29484
rect 30156 29260 30324 29316
rect 29932 28690 29988 28700
rect 30268 27746 30324 29260
rect 30604 28644 30660 32396
rect 30716 32386 30772 32396
rect 30716 31778 30772 31790
rect 30716 31726 30718 31778
rect 30770 31726 30772 31778
rect 30716 31668 30772 31726
rect 30716 30324 30772 31612
rect 30828 30660 30884 38612
rect 30940 38050 30996 38062
rect 30940 37998 30942 38050
rect 30994 37998 30996 38050
rect 30940 37044 30996 37998
rect 31052 37492 31108 37502
rect 31052 37398 31108 37436
rect 31052 37044 31108 37054
rect 30940 36988 31052 37044
rect 31052 36978 31108 36988
rect 31164 35700 31220 38612
rect 31780 38556 31892 38612
rect 31724 38546 31780 38556
rect 31724 37938 31780 37950
rect 31724 37886 31726 37938
rect 31778 37886 31780 37938
rect 31724 37492 31780 37886
rect 31724 37426 31780 37436
rect 31276 37268 31332 37278
rect 31724 37268 31780 37278
rect 31276 37266 31780 37268
rect 31276 37214 31278 37266
rect 31330 37214 31726 37266
rect 31778 37214 31780 37266
rect 31276 37212 31780 37214
rect 31276 36932 31332 37212
rect 31724 37202 31780 37212
rect 31276 36866 31332 36876
rect 31276 36596 31332 36606
rect 31276 36502 31332 36540
rect 31724 35924 31780 35934
rect 31164 35634 31220 35644
rect 31500 35922 31780 35924
rect 31500 35870 31726 35922
rect 31778 35870 31780 35922
rect 31500 35868 31780 35870
rect 31500 34242 31556 35868
rect 31724 35858 31780 35868
rect 31612 35700 31668 35710
rect 31612 35606 31668 35644
rect 31724 35474 31780 35486
rect 31724 35422 31726 35474
rect 31778 35422 31780 35474
rect 31724 35028 31780 35422
rect 31724 34962 31780 34972
rect 31836 34356 31892 38556
rect 32284 37940 32340 39340
rect 33068 38946 33124 40908
rect 33180 40404 33236 41916
rect 33292 41748 33348 41758
rect 33292 40628 33348 41692
rect 33404 40628 33460 42588
rect 33740 42532 33796 42542
rect 33740 42438 33796 42476
rect 33516 41860 33572 41870
rect 33516 41766 33572 41804
rect 33964 41746 34020 41758
rect 33964 41694 33966 41746
rect 34018 41694 34020 41746
rect 33964 41298 34020 41694
rect 33964 41246 33966 41298
rect 34018 41246 34020 41298
rect 33964 41234 34020 41246
rect 34076 41300 34132 43372
rect 34748 43426 34804 44380
rect 34860 44322 34916 44334
rect 34860 44270 34862 44322
rect 34914 44270 34916 44322
rect 34860 43652 34916 44270
rect 35084 44324 35140 44828
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35868 44548 35924 44942
rect 36204 44884 36260 45052
rect 36092 44828 36260 44884
rect 35924 44492 36036 44548
rect 35868 44482 35924 44492
rect 35084 44322 35252 44324
rect 35084 44270 35086 44322
rect 35138 44270 35252 44322
rect 35084 44268 35252 44270
rect 35084 44258 35140 44268
rect 34860 43586 34916 43596
rect 35196 43540 35252 44268
rect 35868 44210 35924 44222
rect 35868 44158 35870 44210
rect 35922 44158 35924 44210
rect 35420 43652 35476 43662
rect 35476 43596 35588 43652
rect 35420 43586 35476 43596
rect 35196 43446 35252 43484
rect 34748 43374 34750 43426
rect 34802 43374 34804 43426
rect 34748 42868 34804 43374
rect 34748 42802 34804 42812
rect 35084 43428 35140 43438
rect 34860 42754 34916 42766
rect 35084 42756 35140 43372
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35308 42866 35364 42878
rect 35308 42814 35310 42866
rect 35362 42814 35364 42866
rect 35196 42756 35252 42766
rect 34860 42702 34862 42754
rect 34914 42702 34916 42754
rect 34188 42642 34244 42654
rect 34188 42590 34190 42642
rect 34242 42590 34244 42642
rect 34188 41748 34244 42590
rect 34412 42532 34468 42542
rect 34188 41682 34244 41692
rect 34300 42530 34468 42532
rect 34300 42478 34414 42530
rect 34466 42478 34468 42530
rect 34300 42476 34468 42478
rect 34300 41412 34356 42476
rect 34412 42466 34468 42476
rect 34524 42530 34580 42542
rect 34524 42478 34526 42530
rect 34578 42478 34580 42530
rect 34412 42196 34468 42206
rect 34412 42082 34468 42140
rect 34412 42030 34414 42082
rect 34466 42030 34468 42082
rect 34412 42018 34468 42030
rect 34300 41346 34356 41356
rect 34076 41234 34132 41244
rect 33628 41188 33684 41198
rect 33628 41094 33684 41132
rect 34524 41076 34580 42478
rect 34636 42532 34692 42542
rect 34636 42530 34804 42532
rect 34636 42478 34638 42530
rect 34690 42478 34804 42530
rect 34636 42476 34804 42478
rect 34636 42466 34692 42476
rect 34748 41860 34804 42476
rect 34748 41766 34804 41804
rect 34860 41748 34916 42702
rect 34860 41682 34916 41692
rect 34972 42754 35252 42756
rect 34972 42702 35198 42754
rect 35250 42702 35252 42754
rect 34972 42700 35252 42702
rect 33740 41020 34580 41076
rect 34860 41188 34916 41198
rect 33628 40628 33684 40638
rect 33740 40628 33796 41020
rect 33404 40572 33572 40628
rect 33292 40562 33348 40572
rect 33404 40404 33460 40414
rect 33180 40402 33460 40404
rect 33180 40350 33406 40402
rect 33458 40350 33460 40402
rect 33180 40348 33460 40350
rect 33404 40338 33460 40348
rect 33516 40290 33572 40572
rect 33628 40626 33796 40628
rect 33628 40574 33630 40626
rect 33682 40574 33796 40626
rect 33628 40572 33796 40574
rect 33852 40852 33908 40862
rect 33628 40562 33684 40572
rect 33516 40238 33518 40290
rect 33570 40238 33572 40290
rect 33516 40226 33572 40238
rect 33068 38894 33070 38946
rect 33122 38894 33124 38946
rect 33068 38882 33124 38894
rect 32956 38836 33012 38846
rect 32284 37874 32340 37884
rect 32732 37940 32788 37950
rect 32508 37828 32564 37838
rect 32060 37716 32116 37726
rect 32060 37490 32116 37660
rect 32060 37438 32062 37490
rect 32114 37438 32116 37490
rect 32060 37426 32116 37438
rect 32396 37492 32452 37502
rect 32396 37398 32452 37436
rect 32508 37378 32564 37772
rect 32508 37326 32510 37378
rect 32562 37326 32564 37378
rect 32508 37314 32564 37326
rect 32284 37156 32340 37166
rect 31948 37044 32004 37054
rect 31948 36482 32004 36988
rect 31948 36430 31950 36482
rect 32002 36430 32004 36482
rect 31948 34914 32004 36430
rect 32284 35698 32340 37100
rect 32732 36594 32788 37884
rect 32732 36542 32734 36594
rect 32786 36542 32788 36594
rect 32732 36530 32788 36542
rect 32508 36372 32564 36382
rect 32508 35922 32564 36316
rect 32508 35870 32510 35922
rect 32562 35870 32564 35922
rect 32508 35858 32564 35870
rect 32620 36260 32676 36270
rect 32284 35646 32286 35698
rect 32338 35646 32340 35698
rect 32284 35634 32340 35646
rect 32620 35476 32676 36204
rect 32620 35410 32676 35420
rect 32844 36258 32900 36270
rect 32844 36206 32846 36258
rect 32898 36206 32900 36258
rect 32284 35364 32340 35374
rect 31948 34862 31950 34914
rect 32002 34862 32004 34914
rect 31948 34850 32004 34862
rect 32172 35140 32228 35150
rect 31500 34190 31502 34242
rect 31554 34190 31556 34242
rect 31500 34178 31556 34190
rect 31612 34300 31892 34356
rect 30940 34132 30996 34142
rect 30940 34038 30996 34076
rect 31164 33124 31220 33134
rect 31164 33030 31220 33068
rect 31500 32564 31556 32574
rect 31500 32470 31556 32508
rect 31276 32450 31332 32462
rect 31276 32398 31278 32450
rect 31330 32398 31332 32450
rect 31276 32004 31332 32398
rect 31276 31948 31556 32004
rect 31388 31780 31444 31790
rect 31388 31686 31444 31724
rect 30940 31666 30996 31678
rect 30940 31614 30942 31666
rect 30994 31614 30996 31666
rect 30940 31556 30996 31614
rect 30940 31490 30996 31500
rect 31276 31666 31332 31678
rect 31276 31614 31278 31666
rect 31330 31614 31332 31666
rect 30940 31332 30996 31342
rect 30940 31218 30996 31276
rect 31164 31332 31220 31342
rect 31276 31332 31332 31614
rect 31220 31276 31332 31332
rect 31500 31668 31556 31948
rect 31612 31892 31668 34300
rect 31836 34132 31892 34142
rect 31836 33348 31892 34076
rect 32172 34130 32228 35084
rect 32172 34078 32174 34130
rect 32226 34078 32228 34130
rect 32172 34066 32228 34078
rect 31612 31826 31668 31836
rect 31724 33346 31892 33348
rect 31724 33294 31838 33346
rect 31890 33294 31892 33346
rect 31724 33292 31892 33294
rect 31164 31266 31220 31276
rect 30940 31166 30942 31218
rect 30994 31166 30996 31218
rect 30940 31154 30996 31166
rect 31500 30994 31556 31612
rect 31500 30942 31502 30994
rect 31554 30942 31556 30994
rect 30828 30604 30996 30660
rect 30716 30258 30772 30268
rect 30716 30100 30772 30110
rect 30716 29986 30772 30044
rect 30716 29934 30718 29986
rect 30770 29934 30772 29986
rect 30716 29204 30772 29934
rect 30716 29138 30772 29148
rect 30828 29988 30884 29998
rect 30828 29314 30884 29932
rect 30828 29262 30830 29314
rect 30882 29262 30884 29314
rect 30828 28868 30884 29262
rect 30828 28802 30884 28812
rect 30604 28588 30884 28644
rect 30268 27694 30270 27746
rect 30322 27694 30324 27746
rect 30268 27682 30324 27694
rect 30716 27748 30772 27758
rect 30716 27654 30772 27692
rect 30156 27188 30212 27198
rect 30156 26908 30212 27132
rect 30380 26964 30436 27002
rect 30156 26852 30324 26908
rect 30380 26898 30436 26908
rect 29820 25666 29876 25676
rect 30156 26516 30212 26526
rect 30156 26402 30212 26460
rect 30268 26514 30324 26852
rect 30268 26462 30270 26514
rect 30322 26462 30324 26514
rect 30268 26450 30324 26462
rect 30604 26852 30660 26862
rect 30156 26350 30158 26402
rect 30210 26350 30212 26402
rect 29260 25508 29316 25518
rect 29260 25172 29316 25452
rect 29932 25396 29988 25406
rect 29260 25106 29316 25116
rect 29372 25394 29988 25396
rect 29372 25342 29934 25394
rect 29986 25342 29988 25394
rect 29372 25340 29988 25342
rect 29260 24052 29316 24062
rect 29372 24052 29428 25340
rect 29932 25330 29988 25340
rect 30156 25396 30212 26350
rect 30492 26404 30548 26414
rect 30492 26310 30548 26348
rect 30604 26290 30660 26796
rect 30716 26850 30772 26862
rect 30716 26798 30718 26850
rect 30770 26798 30772 26850
rect 30716 26516 30772 26798
rect 30716 26450 30772 26460
rect 30828 26404 30884 28588
rect 30940 26628 30996 30604
rect 31052 30212 31108 30250
rect 31052 30146 31108 30156
rect 31388 29428 31444 29438
rect 31388 29334 31444 29372
rect 31052 29204 31108 29214
rect 31052 29110 31108 29148
rect 31276 28644 31332 28654
rect 31276 28550 31332 28588
rect 31164 27860 31220 27870
rect 31164 27766 31220 27804
rect 31500 27412 31556 30942
rect 31612 31666 31668 31678
rect 31612 31614 31614 31666
rect 31666 31614 31668 31666
rect 31612 30100 31668 31614
rect 31724 31218 31780 33292
rect 31836 33282 31892 33292
rect 31948 34018 32004 34030
rect 31948 33966 31950 34018
rect 32002 33966 32004 34018
rect 31836 33124 31892 33134
rect 31948 33124 32004 33966
rect 32060 33572 32116 33582
rect 32060 33234 32116 33516
rect 32060 33182 32062 33234
rect 32114 33182 32116 33234
rect 32060 33170 32116 33182
rect 31892 33068 32004 33124
rect 31836 33058 31892 33068
rect 32284 33012 32340 35308
rect 32844 35140 32900 36206
rect 32844 35074 32900 35084
rect 32620 35028 32676 35038
rect 32620 34934 32676 34972
rect 32956 33460 33012 38780
rect 33852 38836 33908 40796
rect 34860 40852 34916 41132
rect 34860 40786 34916 40796
rect 34524 40628 34580 40638
rect 34972 40628 35028 42700
rect 35196 42690 35252 42700
rect 35308 42756 35364 42814
rect 35308 42690 35364 42700
rect 35420 42756 35476 42766
rect 35532 42756 35588 43596
rect 35756 43540 35812 43550
rect 35644 43428 35700 43438
rect 35644 43334 35700 43372
rect 35420 42754 35588 42756
rect 35420 42702 35422 42754
rect 35474 42702 35588 42754
rect 35420 42700 35588 42702
rect 35756 42756 35812 43484
rect 35868 42980 35924 44158
rect 35980 43988 36036 44492
rect 35980 43922 36036 43932
rect 35980 43652 36036 43662
rect 35980 43558 36036 43596
rect 36092 43650 36148 44828
rect 36988 44436 37044 45726
rect 37100 45666 37156 45678
rect 37100 45614 37102 45666
rect 37154 45614 37156 45666
rect 37100 45220 37156 45614
rect 37100 45154 37156 45164
rect 37212 45108 37268 46508
rect 37324 46498 37380 46508
rect 37660 46116 37716 47180
rect 37772 47234 37828 47404
rect 40012 47460 40068 47470
rect 40012 47366 40068 47404
rect 41244 47460 41300 47470
rect 38780 47348 38836 47358
rect 38780 47254 38836 47292
rect 37772 47182 37774 47234
rect 37826 47182 37828 47234
rect 37772 46900 37828 47182
rect 38332 47236 38388 47246
rect 39228 47236 39284 47246
rect 38332 47234 38612 47236
rect 38332 47182 38334 47234
rect 38386 47182 38612 47234
rect 38332 47180 38612 47182
rect 38332 47170 38388 47180
rect 38556 47124 38612 47180
rect 38892 47234 39284 47236
rect 38892 47182 39230 47234
rect 39282 47182 39284 47234
rect 38892 47180 39284 47182
rect 38556 47068 38724 47124
rect 37772 46834 37828 46844
rect 37884 46562 37940 46574
rect 37884 46510 37886 46562
rect 37938 46510 37940 46562
rect 37660 46060 37828 46116
rect 37212 45042 37268 45052
rect 37324 45890 37380 45902
rect 37660 45892 37716 45902
rect 37324 45838 37326 45890
rect 37378 45838 37380 45890
rect 37100 44994 37156 45006
rect 37100 44942 37102 44994
rect 37154 44942 37156 44994
rect 37100 44660 37156 44942
rect 37324 44884 37380 45838
rect 37436 45890 37716 45892
rect 37436 45838 37662 45890
rect 37714 45838 37716 45890
rect 37436 45836 37716 45838
rect 37436 45108 37492 45836
rect 37660 45826 37716 45836
rect 37436 45106 37604 45108
rect 37436 45054 37438 45106
rect 37490 45054 37604 45106
rect 37436 45052 37604 45054
rect 37436 45042 37492 45052
rect 37324 44818 37380 44828
rect 37100 44604 37492 44660
rect 36988 44370 37044 44380
rect 37212 44436 37268 44446
rect 37212 44342 37268 44380
rect 37100 44212 37156 44222
rect 36764 44210 37156 44212
rect 36764 44158 37102 44210
rect 37154 44158 37156 44210
rect 36764 44156 37156 44158
rect 36092 43598 36094 43650
rect 36146 43598 36148 43650
rect 36092 43586 36148 43598
rect 36204 44098 36260 44110
rect 36204 44046 36206 44098
rect 36258 44046 36260 44098
rect 35868 42914 35924 42924
rect 35756 42754 35924 42756
rect 35756 42702 35758 42754
rect 35810 42702 35924 42754
rect 35756 42700 35924 42702
rect 35420 42690 35476 42700
rect 35756 42690 35812 42700
rect 35644 42532 35700 42542
rect 35644 42530 35812 42532
rect 35644 42478 35646 42530
rect 35698 42478 35812 42530
rect 35644 42476 35812 42478
rect 35644 42466 35700 42476
rect 35084 41860 35140 41870
rect 35196 41860 35252 41870
rect 35140 41858 35252 41860
rect 35140 41806 35198 41858
rect 35250 41806 35252 41858
rect 35140 41804 35252 41806
rect 35084 40852 35140 41804
rect 35196 41794 35252 41804
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 41186 35252 41198
rect 35196 41134 35198 41186
rect 35250 41134 35252 41186
rect 35196 41076 35252 41134
rect 35532 41188 35588 41198
rect 35532 41094 35588 41132
rect 35196 41010 35252 41020
rect 35756 41076 35812 42476
rect 35868 42196 35924 42700
rect 35868 42130 35924 42140
rect 36204 42084 36260 44046
rect 36764 43650 36820 44156
rect 37100 44146 37156 44156
rect 36764 43598 36766 43650
rect 36818 43598 36820 43650
rect 36764 43586 36820 43598
rect 36988 43988 37044 43998
rect 36540 43540 36596 43550
rect 36540 43446 36596 43484
rect 36652 43538 36708 43550
rect 36652 43486 36654 43538
rect 36706 43486 36708 43538
rect 36652 43316 36708 43486
rect 36652 43250 36708 43260
rect 36876 43538 36932 43550
rect 36876 43486 36878 43538
rect 36930 43486 36932 43538
rect 36428 42532 36484 42542
rect 36428 42438 36484 42476
rect 36876 42196 36932 43486
rect 36988 42866 37044 43932
rect 37100 43876 37156 43886
rect 37100 43650 37156 43820
rect 37100 43598 37102 43650
rect 37154 43598 37156 43650
rect 37100 43586 37156 43598
rect 37212 43428 37268 43438
rect 36988 42814 36990 42866
rect 37042 42814 37044 42866
rect 36988 42802 37044 42814
rect 37100 43316 37156 43326
rect 36876 42130 36932 42140
rect 36204 42018 36260 42028
rect 37100 41972 37156 43260
rect 37212 42978 37268 43372
rect 37212 42926 37214 42978
rect 37266 42926 37268 42978
rect 37212 42914 37268 42926
rect 37436 42308 37492 44604
rect 37548 44322 37604 45052
rect 37548 44270 37550 44322
rect 37602 44270 37604 44322
rect 37548 43538 37604 44270
rect 37548 43486 37550 43538
rect 37602 43486 37604 43538
rect 37548 43204 37604 43486
rect 37772 43316 37828 46060
rect 37772 43250 37828 43260
rect 37548 43138 37604 43148
rect 37548 42980 37604 42990
rect 37548 42886 37604 42924
rect 37436 42252 37604 42308
rect 37436 42084 37492 42094
rect 37100 41916 37268 41972
rect 37100 41748 37156 41758
rect 36204 41412 36260 41422
rect 36204 41318 36260 41356
rect 37100 41410 37156 41692
rect 37100 41358 37102 41410
rect 37154 41358 37156 41410
rect 35756 41010 35812 41020
rect 36316 41074 36372 41086
rect 36316 41022 36318 41074
rect 36370 41022 36372 41074
rect 35308 40962 35364 40974
rect 35308 40910 35310 40962
rect 35362 40910 35364 40962
rect 35196 40852 35252 40862
rect 35084 40796 35196 40852
rect 35196 40786 35252 40796
rect 34972 40572 35252 40628
rect 34524 40534 34580 40572
rect 34412 40404 34468 40414
rect 34412 40310 34468 40348
rect 34636 40402 34692 40414
rect 34636 40350 34638 40402
rect 34690 40350 34692 40402
rect 33964 40292 34020 40302
rect 34188 40292 34244 40302
rect 33964 40198 34020 40236
rect 34076 40290 34244 40292
rect 34076 40238 34190 40290
rect 34242 40238 34244 40290
rect 34076 40236 34244 40238
rect 33852 38770 33908 38780
rect 33740 38722 33796 38734
rect 33740 38670 33742 38722
rect 33794 38670 33796 38722
rect 33180 38612 33236 38622
rect 33180 38518 33236 38556
rect 33068 37266 33124 37278
rect 33068 37214 33070 37266
rect 33122 37214 33124 37266
rect 33068 37044 33124 37214
rect 33068 36978 33124 36988
rect 33628 36932 33684 36942
rect 33292 36484 33348 36494
rect 33292 36390 33348 36428
rect 33628 36482 33684 36876
rect 33628 36430 33630 36482
rect 33682 36430 33684 36482
rect 33628 35812 33684 36430
rect 33516 35810 33684 35812
rect 33516 35758 33630 35810
rect 33682 35758 33684 35810
rect 33516 35756 33684 35758
rect 33404 35700 33460 35710
rect 33404 34354 33460 35644
rect 33404 34302 33406 34354
rect 33458 34302 33460 34354
rect 33404 34290 33460 34302
rect 33068 34132 33124 34142
rect 33068 34038 33124 34076
rect 33180 33460 33236 33470
rect 32956 33458 33236 33460
rect 32956 33406 33182 33458
rect 33234 33406 33236 33458
rect 32956 33404 33236 33406
rect 32284 32946 32340 32956
rect 32396 33348 32452 33358
rect 32284 32788 32340 32798
rect 32172 32732 32284 32788
rect 32060 32562 32116 32574
rect 32060 32510 32062 32562
rect 32114 32510 32116 32562
rect 31948 31892 32004 31902
rect 31836 31668 31892 31678
rect 31836 31574 31892 31612
rect 31724 31166 31726 31218
rect 31778 31166 31780 31218
rect 31724 31154 31780 31166
rect 31948 31108 32004 31836
rect 31724 30996 31780 31006
rect 31724 30902 31780 30940
rect 31836 30324 31892 30334
rect 31724 30100 31780 30110
rect 31612 30098 31724 30100
rect 31612 30046 31614 30098
rect 31666 30046 31724 30098
rect 31612 30044 31724 30046
rect 31612 30034 31668 30044
rect 31724 29538 31780 30044
rect 31724 29486 31726 29538
rect 31778 29486 31780 29538
rect 31724 29474 31780 29486
rect 31724 28868 31780 28878
rect 31724 28082 31780 28812
rect 31724 28030 31726 28082
rect 31778 28030 31780 28082
rect 31724 28018 31780 28030
rect 31500 27346 31556 27356
rect 31724 26964 31780 26974
rect 30940 26562 30996 26572
rect 31612 26852 31668 26862
rect 31612 26514 31668 26796
rect 31612 26462 31614 26514
rect 31666 26462 31668 26514
rect 31612 26450 31668 26462
rect 30828 26348 30996 26404
rect 30604 26238 30606 26290
rect 30658 26238 30660 26290
rect 30604 26226 30660 26238
rect 30156 25330 30212 25340
rect 30156 25172 30212 25182
rect 29596 25060 29652 25070
rect 29260 24050 29428 24052
rect 29260 23998 29262 24050
rect 29314 23998 29428 24050
rect 29260 23996 29428 23998
rect 29484 24724 29540 24734
rect 29260 23986 29316 23996
rect 29484 23828 29540 24668
rect 29148 23716 29204 23726
rect 29148 23714 29316 23716
rect 29148 23662 29150 23714
rect 29202 23662 29316 23714
rect 29148 23660 29316 23662
rect 29148 23650 29204 23660
rect 29260 23604 29316 23660
rect 28924 23492 29204 23548
rect 29260 23538 29316 23548
rect 29372 23714 29428 23726
rect 29372 23662 29374 23714
rect 29426 23662 29428 23714
rect 28924 23426 28980 23436
rect 29148 23378 29204 23492
rect 29148 23326 29150 23378
rect 29202 23326 29204 23378
rect 29148 23314 29204 23326
rect 28924 23268 28980 23306
rect 28924 23202 28980 23212
rect 29372 23156 29428 23662
rect 29148 23100 29428 23156
rect 29484 23156 29540 23772
rect 29596 23548 29652 25004
rect 30044 24612 30100 24622
rect 30044 24518 30100 24556
rect 29820 24500 29876 24510
rect 29820 23938 29876 24444
rect 29820 23886 29822 23938
rect 29874 23886 29876 23938
rect 29820 23874 29876 23886
rect 30156 23938 30212 25116
rect 30828 24948 30884 24958
rect 30828 24834 30884 24892
rect 30828 24782 30830 24834
rect 30882 24782 30884 24834
rect 30716 24500 30772 24510
rect 30716 24406 30772 24444
rect 30828 24276 30884 24782
rect 30156 23886 30158 23938
rect 30210 23886 30212 23938
rect 30156 23874 30212 23886
rect 30716 24220 30884 24276
rect 30380 23828 30436 23838
rect 29820 23660 30212 23716
rect 29820 23548 29876 23660
rect 29596 23492 29876 23548
rect 29820 23380 29876 23492
rect 29708 23378 29876 23380
rect 29708 23326 29822 23378
rect 29874 23326 29876 23378
rect 29708 23324 29876 23326
rect 29484 23154 29652 23156
rect 29484 23102 29486 23154
rect 29538 23102 29652 23154
rect 29484 23100 29652 23102
rect 28812 22204 28980 22260
rect 28700 21756 28868 21812
rect 28588 21746 28644 21756
rect 28476 21534 28478 21586
rect 28530 21534 28532 21586
rect 28476 21522 28532 21534
rect 28700 21586 28756 21598
rect 28700 21534 28702 21586
rect 28754 21534 28756 21586
rect 28252 21298 28308 21308
rect 28364 21474 28420 21486
rect 28364 21422 28366 21474
rect 28418 21422 28420 21474
rect 28252 20578 28308 20590
rect 28252 20526 28254 20578
rect 28306 20526 28308 20578
rect 28252 20244 28308 20526
rect 28364 20580 28420 21422
rect 28700 21028 28756 21534
rect 28700 20962 28756 20972
rect 28364 20514 28420 20524
rect 28252 20178 28308 20188
rect 28252 19348 28308 19358
rect 28252 19254 28308 19292
rect 28588 19348 28644 19358
rect 28140 18834 28196 18844
rect 28252 19122 28308 19134
rect 28252 19070 28254 19122
rect 28306 19070 28308 19122
rect 28028 18398 28030 18450
rect 28082 18398 28084 18450
rect 28028 18386 28084 18398
rect 28028 18228 28084 18238
rect 28028 17666 28084 18172
rect 28028 17614 28030 17666
rect 28082 17614 28084 17666
rect 28028 17602 28084 17614
rect 28140 17780 28196 17790
rect 28140 17444 28196 17724
rect 28252 17668 28308 19070
rect 28588 19012 28644 19292
rect 28588 18946 28644 18956
rect 28700 18788 28756 18798
rect 28812 18788 28868 21756
rect 28756 18732 28868 18788
rect 28700 18722 28756 18732
rect 28924 18452 28980 22204
rect 29148 21588 29204 23100
rect 29484 23090 29540 23100
rect 29260 22932 29316 22942
rect 29260 22930 29540 22932
rect 29260 22878 29262 22930
rect 29314 22878 29540 22930
rect 29260 22876 29540 22878
rect 29260 22866 29316 22876
rect 29260 22484 29316 22494
rect 29260 22390 29316 22428
rect 28924 18386 28980 18396
rect 29036 21532 29204 21588
rect 29372 21924 29428 21934
rect 29036 18340 29092 21532
rect 29148 21364 29204 21374
rect 29148 21362 29316 21364
rect 29148 21310 29150 21362
rect 29202 21310 29316 21362
rect 29148 21308 29316 21310
rect 29148 21298 29204 21308
rect 29260 20916 29316 21308
rect 29372 21028 29428 21868
rect 29484 21588 29540 22876
rect 29596 22258 29652 23100
rect 29596 22206 29598 22258
rect 29650 22206 29652 22258
rect 29596 22194 29652 22206
rect 29708 22036 29764 23324
rect 29820 23314 29876 23324
rect 29932 23492 29988 23502
rect 29932 22370 29988 23436
rect 30156 23044 30212 23660
rect 30268 23380 30324 23390
rect 30268 23286 30324 23324
rect 30380 23378 30436 23772
rect 30380 23326 30382 23378
rect 30434 23326 30436 23378
rect 30380 23314 30436 23326
rect 30492 23268 30548 23278
rect 30156 22988 30436 23044
rect 30380 22482 30436 22988
rect 30492 22820 30548 23212
rect 30492 22754 30548 22764
rect 30380 22430 30382 22482
rect 30434 22430 30436 22482
rect 30380 22418 30436 22430
rect 29932 22318 29934 22370
rect 29986 22318 29988 22370
rect 29932 22306 29988 22318
rect 29484 21522 29540 21532
rect 29596 21980 29764 22036
rect 29596 21698 29652 21980
rect 29596 21646 29598 21698
rect 29650 21646 29652 21698
rect 29596 21364 29652 21646
rect 29596 21298 29652 21308
rect 29708 21812 29764 21822
rect 29708 21698 29764 21756
rect 29708 21646 29710 21698
rect 29762 21646 29764 21698
rect 29708 21140 29764 21646
rect 30604 21812 30660 21822
rect 30716 21812 30772 24220
rect 30828 23828 30884 23838
rect 30828 23734 30884 23772
rect 30940 23548 30996 26348
rect 31052 26180 31108 26190
rect 31052 26086 31108 26124
rect 31052 25732 31108 25742
rect 31052 24946 31108 25676
rect 31612 25284 31668 25294
rect 31724 25284 31780 26908
rect 31668 25228 31780 25284
rect 31612 25218 31668 25228
rect 31052 24894 31054 24946
rect 31106 24894 31108 24946
rect 31052 24882 31108 24894
rect 31612 24948 31668 24958
rect 31612 24854 31668 24892
rect 31836 24948 31892 30268
rect 31836 24854 31892 24892
rect 31388 24724 31444 24734
rect 31388 24630 31444 24668
rect 31500 24500 31556 24510
rect 30828 23492 30996 23548
rect 31276 24498 31556 24500
rect 31276 24446 31502 24498
rect 31554 24446 31556 24498
rect 31276 24444 31556 24446
rect 30828 22372 30884 23492
rect 31164 23380 31220 23390
rect 31164 23286 31220 23324
rect 30940 23156 30996 23166
rect 31276 23156 31332 24444
rect 31500 24434 31556 24444
rect 31612 24500 31668 24510
rect 31500 23492 31556 23502
rect 31500 23378 31556 23436
rect 31500 23326 31502 23378
rect 31554 23326 31556 23378
rect 31500 23314 31556 23326
rect 31612 23156 31668 24444
rect 30940 23154 31332 23156
rect 30940 23102 30942 23154
rect 30994 23102 31332 23154
rect 30940 23100 31332 23102
rect 31500 23100 31668 23156
rect 31724 24388 31780 24398
rect 30940 23090 30996 23100
rect 30940 22372 30996 22382
rect 30828 22316 30940 22372
rect 30940 22306 30996 22316
rect 31388 22258 31444 22270
rect 31388 22206 31390 22258
rect 31442 22206 31444 22258
rect 30604 21810 30772 21812
rect 30604 21758 30606 21810
rect 30658 21758 30772 21810
rect 30604 21756 30772 21758
rect 30940 22148 30996 22158
rect 31388 22148 31444 22206
rect 30940 22146 31444 22148
rect 30940 22094 30942 22146
rect 30994 22094 31444 22146
rect 30940 22092 31444 22094
rect 29708 21074 29764 21084
rect 29820 21586 29876 21598
rect 29820 21534 29822 21586
rect 29874 21534 29876 21586
rect 29820 21028 29876 21534
rect 30268 21588 30324 21598
rect 29372 20972 29652 21028
rect 29260 20860 29540 20916
rect 29484 20802 29540 20860
rect 29484 20750 29486 20802
rect 29538 20750 29540 20802
rect 29484 20738 29540 20750
rect 29596 20804 29652 20972
rect 29820 20962 29876 20972
rect 29932 21476 29988 21486
rect 29596 20748 29876 20804
rect 29596 20578 29652 20590
rect 29596 20526 29598 20578
rect 29650 20526 29652 20578
rect 29596 19460 29652 20526
rect 29708 20580 29764 20590
rect 29708 20486 29764 20524
rect 29596 19394 29652 19404
rect 29708 19348 29764 19358
rect 29708 19254 29764 19292
rect 29148 19236 29204 19246
rect 29596 19236 29652 19246
rect 29148 19142 29204 19180
rect 29484 19234 29652 19236
rect 29484 19182 29598 19234
rect 29650 19182 29652 19234
rect 29484 19180 29652 19182
rect 29484 19124 29540 19180
rect 29596 19170 29652 19180
rect 29484 19058 29540 19068
rect 29372 19010 29428 19022
rect 29372 18958 29374 19010
rect 29426 18958 29428 19010
rect 29372 18564 29428 18958
rect 29372 18498 29428 18508
rect 29708 19012 29764 19022
rect 29036 18274 29092 18284
rect 29260 18452 29316 18462
rect 28364 17780 28420 17790
rect 28364 17686 28420 17724
rect 28588 17780 28644 17790
rect 28252 17602 28308 17612
rect 28476 17556 28532 17566
rect 28588 17556 28644 17724
rect 29260 17778 29316 18396
rect 29708 18228 29764 18956
rect 29820 18676 29876 20748
rect 29932 19572 29988 21420
rect 30156 21028 30212 21038
rect 30044 20802 30100 20814
rect 30044 20750 30046 20802
rect 30098 20750 30100 20802
rect 30044 20580 30100 20750
rect 30044 20514 30100 20524
rect 30156 19908 30212 20972
rect 30268 20916 30324 21532
rect 30268 20850 30324 20860
rect 30156 19852 30324 19908
rect 29932 19506 29988 19516
rect 30156 19236 30212 19246
rect 30044 19234 30212 19236
rect 30044 19182 30158 19234
rect 30210 19182 30212 19234
rect 30044 19180 30212 19182
rect 30044 19012 30100 19180
rect 30156 19170 30212 19180
rect 30044 18946 30100 18956
rect 30268 19124 30324 19852
rect 30604 19684 30660 21756
rect 30940 21588 30996 22092
rect 31500 22036 31556 23100
rect 30940 21522 30996 21532
rect 31052 21980 31556 22036
rect 31612 22258 31668 22270
rect 31612 22206 31614 22258
rect 31666 22206 31668 22258
rect 30716 20916 30772 20926
rect 30716 20822 30772 20860
rect 31052 20020 31108 21980
rect 31612 21924 31668 22206
rect 31276 21868 31668 21924
rect 31276 21586 31332 21868
rect 31276 21534 31278 21586
rect 31330 21534 31332 21586
rect 31276 20916 31332 21534
rect 31388 21586 31444 21598
rect 31388 21534 31390 21586
rect 31442 21534 31444 21586
rect 31388 21476 31444 21534
rect 31500 21588 31556 21598
rect 31500 21494 31556 21532
rect 31388 21410 31444 21420
rect 31612 21476 31668 21486
rect 31724 21476 31780 24332
rect 31948 23548 32004 31052
rect 32060 30996 32116 32510
rect 32060 30930 32116 30940
rect 32060 30324 32116 30334
rect 32172 30324 32228 32732
rect 32284 32722 32340 32732
rect 32396 31778 32452 33292
rect 32844 33124 32900 33134
rect 32844 33122 33012 33124
rect 32844 33070 32846 33122
rect 32898 33070 33012 33122
rect 32844 33068 33012 33070
rect 32844 33058 32900 33068
rect 32396 31726 32398 31778
rect 32450 31726 32452 31778
rect 32396 31714 32452 31726
rect 32620 32450 32676 32462
rect 32620 32398 32622 32450
rect 32674 32398 32676 32450
rect 32620 31668 32676 32398
rect 32620 31602 32676 31612
rect 32060 30322 32228 30324
rect 32060 30270 32062 30322
rect 32114 30270 32228 30322
rect 32060 30268 32228 30270
rect 32620 30882 32676 30894
rect 32620 30830 32622 30882
rect 32674 30830 32676 30882
rect 32060 30258 32116 30268
rect 32508 29988 32564 29998
rect 32620 29988 32676 30830
rect 32508 29986 32676 29988
rect 32508 29934 32510 29986
rect 32562 29934 32676 29986
rect 32508 29932 32676 29934
rect 32508 29922 32564 29932
rect 32172 29428 32228 29438
rect 32172 29334 32228 29372
rect 32060 28644 32116 28654
rect 32396 28644 32452 28654
rect 32060 28642 32452 28644
rect 32060 28590 32062 28642
rect 32114 28590 32398 28642
rect 32450 28590 32452 28642
rect 32060 28588 32452 28590
rect 32060 28578 32116 28588
rect 32284 28084 32340 28094
rect 32172 28028 32284 28084
rect 32060 27970 32116 27982
rect 32060 27918 32062 27970
rect 32114 27918 32116 27970
rect 32060 27748 32116 27918
rect 32060 27682 32116 27692
rect 32172 27746 32228 28028
rect 32284 28018 32340 28028
rect 32172 27694 32174 27746
rect 32226 27694 32228 27746
rect 32172 27682 32228 27694
rect 32284 27858 32340 27870
rect 32284 27806 32286 27858
rect 32338 27806 32340 27858
rect 32284 27748 32340 27806
rect 32284 27682 32340 27692
rect 32396 26962 32452 28588
rect 32508 27860 32564 27870
rect 32508 27766 32564 27804
rect 32396 26910 32398 26962
rect 32450 26910 32452 26962
rect 32060 26852 32116 26862
rect 32060 26514 32116 26796
rect 32060 26462 32062 26514
rect 32114 26462 32116 26514
rect 32060 26450 32116 26462
rect 32060 25732 32116 25742
rect 32060 25618 32116 25676
rect 32060 25566 32062 25618
rect 32114 25566 32116 25618
rect 32060 25554 32116 25566
rect 32396 25172 32452 26910
rect 32508 26852 32564 26862
rect 32508 26514 32564 26796
rect 32508 26462 32510 26514
rect 32562 26462 32564 26514
rect 32508 26450 32564 26462
rect 32620 25508 32676 29932
rect 32956 29204 33012 33068
rect 33180 32788 33236 33404
rect 33516 33348 33572 35756
rect 33628 35746 33684 35756
rect 33740 35476 33796 38670
rect 34076 38668 34132 40236
rect 34188 40226 34244 40236
rect 34636 39844 34692 40350
rect 34636 39778 34692 39788
rect 34972 40404 35028 40414
rect 34412 39620 34468 39630
rect 34860 39620 34916 39630
rect 33852 38612 33908 38622
rect 33852 37378 33908 38556
rect 33964 38612 34132 38668
rect 34188 39618 34916 39620
rect 34188 39566 34414 39618
rect 34466 39566 34862 39618
rect 34914 39566 34916 39618
rect 34188 39564 34916 39566
rect 33964 38162 34020 38612
rect 33964 38110 33966 38162
rect 34018 38110 34020 38162
rect 33964 38052 34020 38110
rect 33964 37986 34020 37996
rect 33852 37326 33854 37378
rect 33906 37326 33908 37378
rect 33852 37314 33908 37326
rect 34076 37268 34132 37278
rect 34076 36596 34132 37212
rect 33740 35410 33796 35420
rect 33852 35812 33908 35822
rect 33628 33348 33684 33358
rect 33572 33346 33684 33348
rect 33572 33294 33630 33346
rect 33682 33294 33684 33346
rect 33572 33292 33684 33294
rect 33516 33254 33572 33292
rect 33628 33282 33684 33292
rect 33180 32722 33236 32732
rect 33292 33236 33348 33246
rect 33292 32786 33348 33180
rect 33292 32734 33294 32786
rect 33346 32734 33348 32786
rect 33292 32722 33348 32734
rect 33180 32452 33236 32462
rect 33180 32358 33236 32396
rect 33740 32450 33796 32462
rect 33740 32398 33742 32450
rect 33794 32398 33796 32450
rect 33628 32340 33684 32350
rect 33404 32338 33684 32340
rect 33404 32286 33630 32338
rect 33682 32286 33684 32338
rect 33404 32284 33684 32286
rect 33404 32116 33460 32284
rect 33628 32274 33684 32284
rect 33068 32060 33460 32116
rect 33628 32116 33684 32126
rect 33068 31890 33124 32060
rect 33068 31838 33070 31890
rect 33122 31838 33124 31890
rect 33068 31826 33124 31838
rect 33180 30996 33236 31006
rect 33068 30322 33124 30334
rect 33068 30270 33070 30322
rect 33122 30270 33124 30322
rect 33068 29652 33124 30270
rect 33068 29586 33124 29596
rect 33180 29540 33236 30940
rect 33292 30882 33348 30894
rect 33292 30830 33294 30882
rect 33346 30830 33348 30882
rect 33292 29764 33348 30830
rect 33404 30770 33460 30782
rect 33404 30718 33406 30770
rect 33458 30718 33460 30770
rect 33404 30212 33460 30718
rect 33404 30146 33460 30156
rect 33292 29698 33348 29708
rect 33516 29652 33572 29662
rect 33404 29540 33460 29550
rect 33180 29538 33460 29540
rect 33180 29486 33406 29538
rect 33458 29486 33460 29538
rect 33180 29484 33460 29486
rect 33068 29428 33124 29438
rect 33068 29334 33124 29372
rect 32956 29148 33348 29204
rect 33180 28530 33236 28542
rect 33180 28478 33182 28530
rect 33234 28478 33236 28530
rect 33180 28084 33236 28478
rect 33180 28018 33236 28028
rect 33068 27746 33124 27758
rect 33068 27694 33070 27746
rect 33122 27694 33124 27746
rect 32732 26292 32788 26302
rect 32732 25730 32788 26236
rect 33068 26180 33124 27694
rect 33180 27636 33236 27646
rect 33180 27542 33236 27580
rect 33292 26852 33348 29148
rect 33292 26786 33348 26796
rect 33404 26292 33460 29484
rect 33516 29428 33572 29596
rect 33516 27970 33572 29372
rect 33628 29204 33684 32060
rect 33740 31892 33796 32398
rect 33740 31826 33796 31836
rect 33852 31332 33908 35756
rect 33852 31266 33908 31276
rect 33964 34020 34020 34030
rect 33852 30994 33908 31006
rect 33852 30942 33854 30994
rect 33906 30942 33908 30994
rect 33852 30436 33908 30942
rect 33852 30370 33908 30380
rect 33964 29988 34020 33964
rect 34076 32116 34132 36540
rect 34188 35700 34244 39564
rect 34412 39554 34468 39564
rect 34860 39554 34916 39564
rect 34860 38836 34916 38846
rect 34972 38836 35028 40348
rect 35196 40290 35252 40572
rect 35196 40238 35198 40290
rect 35250 40238 35252 40290
rect 35196 40180 35252 40238
rect 35308 40180 35364 40910
rect 35420 40964 35476 40974
rect 35420 40870 35476 40908
rect 35644 40962 35700 40974
rect 35644 40910 35646 40962
rect 35698 40910 35700 40962
rect 35308 40124 35588 40180
rect 35196 40114 35252 40124
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35308 39844 35364 39854
rect 35308 39618 35364 39788
rect 35308 39566 35310 39618
rect 35362 39566 35364 39618
rect 35308 38948 35364 39566
rect 35420 39620 35476 39630
rect 35532 39620 35588 40124
rect 35644 39732 35700 40910
rect 36204 40962 36260 40974
rect 36204 40910 36206 40962
rect 36258 40910 36260 40962
rect 36092 40516 36148 40526
rect 35644 39676 35812 39732
rect 35420 39618 35532 39620
rect 35420 39566 35422 39618
rect 35474 39566 35532 39618
rect 35420 39564 35532 39566
rect 35420 39554 35476 39564
rect 35532 39526 35588 39564
rect 35532 39394 35588 39406
rect 35532 39342 35534 39394
rect 35586 39342 35588 39394
rect 35420 38948 35476 38958
rect 35308 38892 35420 38948
rect 35420 38854 35476 38892
rect 34860 38834 35028 38836
rect 34860 38782 34862 38834
rect 34914 38782 35028 38834
rect 34860 38780 35028 38782
rect 34300 38724 34356 38762
rect 34300 38658 34356 38668
rect 34860 38164 34916 38780
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34860 38098 34916 38108
rect 35196 38220 35476 38276
rect 35196 38164 35252 38220
rect 35196 38098 35252 38108
rect 34860 37940 34916 37950
rect 34860 37846 34916 37884
rect 34972 37938 35028 37950
rect 34972 37886 34974 37938
rect 35026 37886 35028 37938
rect 34412 37826 34468 37838
rect 34412 37774 34414 37826
rect 34466 37774 34468 37826
rect 34412 37156 34468 37774
rect 34412 37090 34468 37100
rect 34972 37604 35028 37886
rect 34972 36708 35028 37548
rect 34972 36642 35028 36652
rect 35084 37938 35140 37950
rect 35084 37886 35086 37938
rect 35138 37886 35140 37938
rect 34300 36372 34356 36382
rect 34300 36278 34356 36316
rect 34188 35634 34244 35644
rect 35084 35140 35140 37886
rect 35420 37044 35476 38220
rect 35532 38164 35588 39342
rect 35644 39396 35700 39406
rect 35644 39302 35700 39340
rect 35756 39394 35812 39676
rect 35756 39342 35758 39394
rect 35810 39342 35812 39394
rect 35756 39172 35812 39342
rect 35980 39620 36036 39630
rect 35868 39172 35924 39182
rect 35532 38098 35588 38108
rect 35644 39116 35868 39172
rect 35644 38050 35700 39116
rect 35868 39106 35924 39116
rect 35644 37998 35646 38050
rect 35698 37998 35700 38050
rect 35644 37986 35700 37998
rect 35756 38500 35812 38510
rect 35756 37940 35812 38444
rect 35756 37846 35812 37884
rect 35868 37828 35924 37838
rect 35868 37734 35924 37772
rect 35980 37826 36036 39564
rect 36092 38836 36148 40460
rect 36204 40292 36260 40910
rect 36204 40226 36260 40236
rect 36316 39732 36372 41022
rect 36876 41076 36932 41086
rect 36988 41076 37044 41086
rect 36932 41074 37044 41076
rect 36932 41022 36990 41074
rect 37042 41022 37044 41074
rect 36932 41020 37044 41022
rect 36428 40404 36484 40414
rect 36428 39842 36484 40348
rect 36540 40292 36596 40302
rect 36596 40236 36708 40292
rect 36540 40226 36596 40236
rect 36428 39790 36430 39842
rect 36482 39790 36484 39842
rect 36428 39778 36484 39790
rect 36204 39676 36372 39732
rect 36204 38948 36260 39676
rect 36316 39508 36372 39518
rect 36316 39414 36372 39452
rect 36316 38948 36372 38958
rect 36204 38946 36372 38948
rect 36204 38894 36318 38946
rect 36370 38894 36372 38946
rect 36204 38892 36372 38894
rect 36092 38780 36260 38836
rect 36204 38722 36260 38780
rect 36204 38670 36206 38722
rect 36258 38670 36260 38722
rect 36204 38658 36260 38670
rect 35980 37774 35982 37826
rect 36034 37774 36036 37826
rect 35980 37716 36036 37774
rect 35980 37650 36036 37660
rect 36092 38500 36148 38510
rect 35980 37156 36036 37166
rect 36092 37156 36148 38444
rect 36204 38052 36260 38062
rect 36316 38052 36372 38892
rect 36652 38834 36708 40236
rect 36652 38782 36654 38834
rect 36706 38782 36708 38834
rect 36260 37996 36372 38052
rect 36428 38500 36484 38510
rect 36204 37958 36260 37996
rect 36428 37266 36484 38444
rect 36428 37214 36430 37266
rect 36482 37214 36484 37266
rect 36428 37202 36484 37214
rect 35980 37154 36148 37156
rect 35980 37102 35982 37154
rect 36034 37102 36148 37154
rect 35980 37100 36148 37102
rect 35980 37090 36036 37100
rect 35420 36988 35588 37044
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35532 35140 35588 36988
rect 35084 35084 35252 35140
rect 34748 35026 34804 35038
rect 34748 34974 34750 35026
rect 34802 34974 34804 35026
rect 34748 34916 34804 34974
rect 35084 34916 35140 34926
rect 34748 34914 35140 34916
rect 34748 34862 35086 34914
rect 35138 34862 35140 34914
rect 34748 34860 35140 34862
rect 34748 34130 34804 34860
rect 35084 34850 35140 34860
rect 34748 34078 34750 34130
rect 34802 34078 34804 34130
rect 34748 34066 34804 34078
rect 34524 34020 34580 34030
rect 34524 34018 34692 34020
rect 34524 33966 34526 34018
rect 34578 33966 34692 34018
rect 34524 33964 34692 33966
rect 34524 33954 34580 33964
rect 34300 33236 34356 33246
rect 34300 33142 34356 33180
rect 34300 32788 34356 32798
rect 34300 32694 34356 32732
rect 34076 32050 34132 32060
rect 34188 32562 34244 32574
rect 34188 32510 34190 32562
rect 34242 32510 34244 32562
rect 34188 31444 34244 32510
rect 34524 32562 34580 32574
rect 34524 32510 34526 32562
rect 34578 32510 34580 32562
rect 34412 32452 34468 32462
rect 34412 32358 34468 32396
rect 34188 31378 34244 31388
rect 34076 31332 34132 31342
rect 34076 31218 34132 31276
rect 34524 31332 34580 32510
rect 34524 31266 34580 31276
rect 34076 31166 34078 31218
rect 34130 31166 34132 31218
rect 34076 31154 34132 31166
rect 34412 31108 34468 31118
rect 34412 31014 34468 31052
rect 33964 29922 34020 29932
rect 34188 30996 34244 31006
rect 33740 29428 33796 29438
rect 33740 29334 33796 29372
rect 33964 29426 34020 29438
rect 33964 29374 33966 29426
rect 34018 29374 34020 29426
rect 33852 29316 33908 29326
rect 33852 29222 33908 29260
rect 33628 29148 33796 29204
rect 33516 27918 33518 27970
rect 33570 27918 33572 27970
rect 33516 27906 33572 27918
rect 33628 27972 33684 27982
rect 33628 27878 33684 27916
rect 33740 26908 33796 29148
rect 33852 27972 33908 27982
rect 33964 27972 34020 29374
rect 33852 27970 34020 27972
rect 33852 27918 33854 27970
rect 33906 27918 34020 27970
rect 33852 27916 34020 27918
rect 34076 28644 34132 28654
rect 34076 27970 34132 28588
rect 34076 27918 34078 27970
rect 34130 27918 34132 27970
rect 33852 27636 33908 27916
rect 34076 27906 34132 27918
rect 33852 27570 33908 27580
rect 33404 26226 33460 26236
rect 33628 26852 33796 26908
rect 34076 27524 34132 27534
rect 33068 26086 33124 26124
rect 33068 25844 33124 25854
rect 32732 25678 32734 25730
rect 32786 25678 32788 25730
rect 32732 25666 32788 25678
rect 32844 25732 32900 25742
rect 32396 25106 32452 25116
rect 32508 25452 32676 25508
rect 32060 24724 32116 24734
rect 32060 24630 32116 24668
rect 31948 23492 32116 23548
rect 31948 23268 32004 23278
rect 31948 23174 32004 23212
rect 31948 22930 32004 22942
rect 31948 22878 31950 22930
rect 32002 22878 32004 22930
rect 31948 22820 32004 22878
rect 31836 22764 32004 22820
rect 31836 22370 31892 22764
rect 32060 22708 32116 23492
rect 31836 22318 31838 22370
rect 31890 22318 31892 22370
rect 31836 22148 31892 22318
rect 31836 22082 31892 22092
rect 31948 22652 32116 22708
rect 31948 22260 32004 22652
rect 32060 22484 32116 22494
rect 32396 22484 32452 22494
rect 32060 22482 32452 22484
rect 32060 22430 32062 22482
rect 32114 22430 32398 22482
rect 32450 22430 32452 22482
rect 32060 22428 32452 22430
rect 32060 22418 32116 22428
rect 32396 22418 32452 22428
rect 32172 22260 32228 22270
rect 31948 22204 32172 22260
rect 31948 21924 32004 22204
rect 32172 22166 32228 22204
rect 31836 21868 32004 21924
rect 31836 21588 31892 21868
rect 32172 21812 32228 21822
rect 31948 21756 32172 21812
rect 31948 21698 32004 21756
rect 32172 21746 32228 21756
rect 31948 21646 31950 21698
rect 32002 21646 32004 21698
rect 31948 21634 32004 21646
rect 31836 21522 31892 21532
rect 32508 21588 32564 25452
rect 32844 25396 32900 25676
rect 33068 25732 33124 25788
rect 33068 25730 33348 25732
rect 33068 25678 33070 25730
rect 33122 25678 33348 25730
rect 33068 25676 33348 25678
rect 33068 25666 33124 25676
rect 32620 25394 32900 25396
rect 32620 25342 32846 25394
rect 32898 25342 32900 25394
rect 32620 25340 32900 25342
rect 32620 24946 32676 25340
rect 32844 25330 32900 25340
rect 33180 25172 33236 25182
rect 32620 24894 32622 24946
rect 32674 24894 32676 24946
rect 32620 23378 32676 24894
rect 32956 24948 33012 24958
rect 32956 24050 33012 24892
rect 33180 24722 33236 25116
rect 33180 24670 33182 24722
rect 33234 24670 33236 24722
rect 33180 24658 33236 24670
rect 32956 23998 32958 24050
rect 33010 23998 33012 24050
rect 32956 23986 33012 23998
rect 32620 23326 32622 23378
rect 32674 23326 32676 23378
rect 32620 23314 32676 23326
rect 33292 23378 33348 25676
rect 33516 25620 33572 25630
rect 33516 25526 33572 25564
rect 33292 23326 33294 23378
rect 33346 23326 33348 23378
rect 33292 23314 33348 23326
rect 33404 25394 33460 25406
rect 33404 25342 33406 25394
rect 33458 25342 33460 25394
rect 32620 22932 32676 22942
rect 33404 22932 33460 25342
rect 33516 23714 33572 23726
rect 33516 23662 33518 23714
rect 33570 23662 33572 23714
rect 33516 23492 33572 23662
rect 33516 23426 33572 23436
rect 33628 23380 33684 26852
rect 33852 26180 33908 26190
rect 33908 26124 34020 26180
rect 33852 26114 33908 26124
rect 33740 25508 33796 25518
rect 33740 25414 33796 25452
rect 33964 25506 34020 26124
rect 33964 25454 33966 25506
rect 34018 25454 34020 25506
rect 33964 25396 34020 25454
rect 33964 25330 34020 25340
rect 33852 24610 33908 24622
rect 33852 24558 33854 24610
rect 33906 24558 33908 24610
rect 33852 24164 33908 24558
rect 33964 24164 34020 24174
rect 33852 24108 33964 24164
rect 33964 24098 34020 24108
rect 33852 23828 33908 23838
rect 33852 23826 34020 23828
rect 33852 23774 33854 23826
rect 33906 23774 34020 23826
rect 33852 23772 34020 23774
rect 33852 23762 33908 23772
rect 33628 23314 33684 23324
rect 33740 23714 33796 23726
rect 33740 23662 33742 23714
rect 33794 23662 33796 23714
rect 33740 23268 33796 23662
rect 33964 23492 34020 23772
rect 33964 23426 34020 23436
rect 33740 23212 34020 23268
rect 33628 23044 33684 23054
rect 33740 23044 33796 23212
rect 33628 23042 33796 23044
rect 33628 22990 33630 23042
rect 33682 22990 33796 23042
rect 33628 22988 33796 22990
rect 33852 23044 33908 23054
rect 33628 22978 33684 22988
rect 33852 22950 33908 22988
rect 32620 22930 33460 22932
rect 32620 22878 32622 22930
rect 32674 22878 33460 22930
rect 32620 22876 33460 22878
rect 33516 22932 33572 22942
rect 32620 22866 32676 22876
rect 33292 22594 33348 22606
rect 33292 22542 33294 22594
rect 33346 22542 33348 22594
rect 32620 22260 32676 22270
rect 32620 22166 32676 22204
rect 33068 22260 33124 22270
rect 33068 22166 33124 22204
rect 33068 21812 33124 21822
rect 33068 21718 33124 21756
rect 33292 21810 33348 22542
rect 33292 21758 33294 21810
rect 33346 21758 33348 21810
rect 33292 21746 33348 21758
rect 31668 21420 31780 21476
rect 32396 21476 32452 21486
rect 31612 21410 31668 21420
rect 32396 21382 32452 21420
rect 31276 20850 31332 20860
rect 31052 19954 31108 19964
rect 31612 20580 31668 20590
rect 31164 19908 31220 19918
rect 31164 19906 31556 19908
rect 31164 19854 31166 19906
rect 31218 19854 31556 19906
rect 31164 19852 31556 19854
rect 31164 19842 31220 19852
rect 31052 19796 31108 19806
rect 30604 19618 30660 19628
rect 30940 19794 31108 19796
rect 30940 19742 31054 19794
rect 31106 19742 31108 19794
rect 30940 19740 31108 19742
rect 30604 19460 30660 19470
rect 30492 19348 30548 19358
rect 30492 19254 30548 19292
rect 30604 19234 30660 19404
rect 30604 19182 30606 19234
rect 30658 19182 30660 19234
rect 30604 19170 30660 19182
rect 29820 18620 30100 18676
rect 29708 18162 29764 18172
rect 29820 18452 29876 18462
rect 29260 17726 29262 17778
rect 29314 17726 29316 17778
rect 28476 17554 28644 17556
rect 28476 17502 28478 17554
rect 28530 17502 28644 17554
rect 28476 17500 28644 17502
rect 29036 17668 29092 17678
rect 28476 17490 28532 17500
rect 28140 17378 28196 17388
rect 28140 16772 28196 16782
rect 27468 16380 27972 16436
rect 28028 16660 28084 16670
rect 27356 16212 27412 16222
rect 27132 16210 27412 16212
rect 27132 16158 27358 16210
rect 27410 16158 27412 16210
rect 27132 16156 27412 16158
rect 27132 15314 27188 16156
rect 27356 16146 27412 16156
rect 27468 16098 27524 16380
rect 27692 16212 27748 16222
rect 27468 16046 27470 16098
rect 27522 16046 27524 16098
rect 27244 15988 27300 15998
rect 27244 15894 27300 15932
rect 27132 15262 27134 15314
rect 27186 15262 27188 15314
rect 27132 15250 27188 15262
rect 27468 14532 27524 16046
rect 27580 16100 27636 16110
rect 27580 15314 27636 16044
rect 27692 15986 27748 16156
rect 28028 16098 28084 16604
rect 28028 16046 28030 16098
rect 28082 16046 28084 16098
rect 28028 15988 28084 16046
rect 27692 15934 27694 15986
rect 27746 15934 27748 15986
rect 27692 15922 27748 15934
rect 27804 15932 28028 15988
rect 27804 15540 27860 15932
rect 28028 15922 28084 15932
rect 27580 15262 27582 15314
rect 27634 15262 27636 15314
rect 27580 15250 27636 15262
rect 27692 15484 27860 15540
rect 27692 15148 27748 15484
rect 27356 14476 27524 14532
rect 27580 15092 27748 15148
rect 27804 15316 27860 15326
rect 26572 13906 26628 13916
rect 26684 14028 27300 14084
rect 26684 13970 26740 14028
rect 26684 13918 26686 13970
rect 26738 13918 26740 13970
rect 26684 13906 26740 13918
rect 26012 13636 26068 13646
rect 25900 13634 26068 13636
rect 25900 13582 26014 13634
rect 26066 13582 26068 13634
rect 25900 13580 26068 13582
rect 25452 13522 25508 13534
rect 25788 13524 25844 13534
rect 25452 13470 25454 13522
rect 25506 13470 25508 13522
rect 25452 12628 25508 13470
rect 25452 12562 25508 12572
rect 25564 13522 25844 13524
rect 25564 13470 25790 13522
rect 25842 13470 25844 13522
rect 25564 13468 25844 13470
rect 25340 11554 25396 11564
rect 25452 12404 25508 12414
rect 25564 12404 25620 13468
rect 25788 13458 25844 13468
rect 25452 12402 25620 12404
rect 25452 12350 25454 12402
rect 25506 12350 25620 12402
rect 25452 12348 25620 12350
rect 25676 12404 25732 12414
rect 25900 12404 25956 13580
rect 26012 13570 26068 13580
rect 26572 13636 26628 13646
rect 26460 13188 26516 13198
rect 25676 12402 26404 12404
rect 25676 12350 25678 12402
rect 25730 12350 26404 12402
rect 25676 12348 26404 12350
rect 25452 11172 25508 12348
rect 25676 12338 25732 12348
rect 26124 12180 26180 12190
rect 26124 12086 26180 12124
rect 25564 12068 25620 12078
rect 25564 11974 25620 12012
rect 26348 11956 26404 12348
rect 26460 12178 26516 13132
rect 26572 13074 26628 13580
rect 26572 13022 26574 13074
rect 26626 13022 26628 13074
rect 26572 13010 26628 13022
rect 26908 12404 26964 14028
rect 27244 13970 27300 14028
rect 27244 13918 27246 13970
rect 27298 13918 27300 13970
rect 27244 13906 27300 13918
rect 27020 13748 27076 13758
rect 27076 13692 27188 13748
rect 27020 13654 27076 13692
rect 26908 12348 27076 12404
rect 26460 12126 26462 12178
rect 26514 12126 26516 12178
rect 26460 12114 26516 12126
rect 26796 12292 26852 12302
rect 26796 12066 26852 12236
rect 26796 12014 26798 12066
rect 26850 12014 26852 12066
rect 26796 12002 26852 12014
rect 26908 12180 26964 12190
rect 26348 11900 26628 11956
rect 25788 11620 25844 11630
rect 25452 11116 25620 11172
rect 25340 10612 25396 10622
rect 25340 10610 25508 10612
rect 25340 10558 25342 10610
rect 25394 10558 25508 10610
rect 25340 10556 25508 10558
rect 25340 10546 25396 10556
rect 25340 9268 25396 9278
rect 25228 9266 25396 9268
rect 25228 9214 25342 9266
rect 25394 9214 25396 9266
rect 25228 9212 25396 9214
rect 25340 9156 25396 9212
rect 25340 9090 25396 9100
rect 24780 8978 24836 8988
rect 25228 9042 25284 9054
rect 25228 8990 25230 9042
rect 25282 8990 25284 9042
rect 24668 8530 24724 8540
rect 25228 8260 25284 8990
rect 25228 8194 25284 8204
rect 24892 8148 24948 8158
rect 24556 7410 24612 7420
rect 24780 7924 24836 7934
rect 24780 7364 24836 7868
rect 23996 7252 24052 7262
rect 24556 7252 24612 7262
rect 24780 7252 24836 7308
rect 23996 7250 24500 7252
rect 23996 7198 23998 7250
rect 24050 7198 24500 7250
rect 23996 7196 24500 7198
rect 23996 7186 24052 7196
rect 24220 6692 24276 6702
rect 24276 6636 24388 6692
rect 24220 6626 24276 6636
rect 24220 6020 24276 6030
rect 24220 5926 24276 5964
rect 23772 5170 23828 5180
rect 24332 5124 24388 6636
rect 24444 5906 24500 7196
rect 24556 7250 24836 7252
rect 24556 7198 24558 7250
rect 24610 7198 24836 7250
rect 24556 7196 24836 7198
rect 24556 7186 24612 7196
rect 24892 7028 24948 8092
rect 25228 8036 25284 8046
rect 25228 7586 25284 7980
rect 25228 7534 25230 7586
rect 25282 7534 25284 7586
rect 25228 7522 25284 7534
rect 25340 7812 25396 7822
rect 25340 7474 25396 7756
rect 25340 7422 25342 7474
rect 25394 7422 25396 7474
rect 25340 7410 25396 7422
rect 24444 5854 24446 5906
rect 24498 5854 24500 5906
rect 24444 5842 24500 5854
rect 24556 6972 24948 7028
rect 24108 5122 24388 5124
rect 24108 5070 24334 5122
rect 24386 5070 24388 5122
rect 24108 5068 24388 5070
rect 24108 4340 24164 5068
rect 24332 5058 24388 5068
rect 24556 4562 24612 6972
rect 25452 6802 25508 10556
rect 25564 9716 25620 11116
rect 25788 10948 25844 11564
rect 26572 11506 26628 11900
rect 26572 11454 26574 11506
rect 26626 11454 26628 11506
rect 26572 11442 26628 11454
rect 26908 11394 26964 12124
rect 26908 11342 26910 11394
rect 26962 11342 26964 11394
rect 26908 11330 26964 11342
rect 25788 10882 25844 10892
rect 26460 11172 26516 11182
rect 26012 10500 26068 10510
rect 25676 10498 26068 10500
rect 25676 10446 26014 10498
rect 26066 10446 26068 10498
rect 25676 10444 26068 10446
rect 25676 9938 25732 10444
rect 26012 10434 26068 10444
rect 25788 10276 25844 10286
rect 25788 10050 25844 10220
rect 25788 9998 25790 10050
rect 25842 9998 25844 10050
rect 25788 9986 25844 9998
rect 26460 10050 26516 11116
rect 26460 9998 26462 10050
rect 26514 9998 26516 10050
rect 26460 9986 26516 9998
rect 26684 10500 26740 10510
rect 25676 9886 25678 9938
rect 25730 9886 25732 9938
rect 25676 9874 25732 9886
rect 26684 9938 26740 10444
rect 26684 9886 26686 9938
rect 26738 9886 26740 9938
rect 26684 9874 26740 9886
rect 26124 9716 26180 9726
rect 25564 9714 26180 9716
rect 25564 9662 25566 9714
rect 25618 9662 26126 9714
rect 26178 9662 26180 9714
rect 25564 9660 26180 9662
rect 25564 9650 25620 9660
rect 26124 9650 26180 9660
rect 25564 9268 25620 9278
rect 25564 9174 25620 9212
rect 27020 9268 27076 12348
rect 27132 9826 27188 13692
rect 27356 13636 27412 14476
rect 27580 14420 27636 15092
rect 27804 14644 27860 15260
rect 27916 14644 27972 14654
rect 27804 14642 27972 14644
rect 27804 14590 27918 14642
rect 27970 14590 27972 14642
rect 27804 14588 27972 14590
rect 27916 14578 27972 14588
rect 28028 14532 28084 14542
rect 28140 14532 28196 16716
rect 28364 16210 28420 16222
rect 28364 16158 28366 16210
rect 28418 16158 28420 16210
rect 28252 16100 28308 16110
rect 28252 16006 28308 16044
rect 28028 14530 28196 14532
rect 28028 14478 28030 14530
rect 28082 14478 28196 14530
rect 28028 14476 28196 14478
rect 28252 15426 28308 15438
rect 28252 15374 28254 15426
rect 28306 15374 28308 15426
rect 28028 14466 28084 14476
rect 27804 14420 27860 14430
rect 27580 14418 27860 14420
rect 27580 14366 27806 14418
rect 27858 14366 27860 14418
rect 27580 14364 27860 14366
rect 27804 14354 27860 14364
rect 27356 13570 27412 13580
rect 27468 14306 27524 14318
rect 27468 14254 27470 14306
rect 27522 14254 27524 14306
rect 27468 13412 27524 14254
rect 27468 13346 27524 13356
rect 27692 13748 27748 13758
rect 27244 13076 27300 13086
rect 27692 13076 27748 13692
rect 28252 13748 28308 15374
rect 28364 14530 28420 16158
rect 28476 16212 28532 16222
rect 28476 15986 28532 16156
rect 28476 15934 28478 15986
rect 28530 15934 28532 15986
rect 28476 15922 28532 15934
rect 28588 16100 28644 16110
rect 28364 14478 28366 14530
rect 28418 14478 28420 14530
rect 28364 14466 28420 14478
rect 28252 13682 28308 13692
rect 28028 13634 28084 13646
rect 28028 13582 28030 13634
rect 28082 13582 28084 13634
rect 27916 13522 27972 13534
rect 27916 13470 27918 13522
rect 27970 13470 27972 13522
rect 27804 13188 27860 13198
rect 27916 13188 27972 13470
rect 27860 13132 27972 13188
rect 28028 13300 28084 13582
rect 27804 13122 27860 13132
rect 27244 13074 27748 13076
rect 27244 13022 27246 13074
rect 27298 13022 27748 13074
rect 27244 13020 27748 13022
rect 27244 13010 27300 13020
rect 27692 12962 27748 13020
rect 27692 12910 27694 12962
rect 27746 12910 27748 12962
rect 27692 12898 27748 12910
rect 27916 12850 27972 12862
rect 27916 12798 27918 12850
rect 27970 12798 27972 12850
rect 27916 12292 27972 12798
rect 28028 12852 28084 13244
rect 28364 13634 28420 13646
rect 28364 13582 28366 13634
rect 28418 13582 28420 13634
rect 28364 13522 28420 13582
rect 28364 13470 28366 13522
rect 28418 13470 28420 13522
rect 28364 13076 28420 13470
rect 28364 13010 28420 13020
rect 28588 12962 28644 16044
rect 29036 15314 29092 17612
rect 29148 17556 29204 17566
rect 29148 16210 29204 17500
rect 29260 17444 29316 17726
rect 29260 17378 29316 17388
rect 29596 17892 29652 17902
rect 29596 16548 29652 17836
rect 29820 16770 29876 18396
rect 30044 18116 30100 18620
rect 30156 18340 30212 18350
rect 30268 18340 30324 19068
rect 30828 19122 30884 19134
rect 30828 19070 30830 19122
rect 30882 19070 30884 19122
rect 30380 19012 30436 19050
rect 30380 18946 30436 18956
rect 30828 19012 30884 19070
rect 30828 18946 30884 18956
rect 30828 18564 30884 18574
rect 30716 18452 30772 18462
rect 30828 18452 30884 18508
rect 30716 18450 30884 18452
rect 30716 18398 30718 18450
rect 30770 18398 30884 18450
rect 30716 18396 30884 18398
rect 30716 18386 30772 18396
rect 30156 18338 30324 18340
rect 30156 18286 30158 18338
rect 30210 18286 30324 18338
rect 30156 18284 30324 18286
rect 30604 18340 30660 18350
rect 30156 18274 30212 18284
rect 30604 18246 30660 18284
rect 30940 18228 30996 19740
rect 31052 19730 31108 19740
rect 31276 19348 31332 19358
rect 31276 19254 31332 19292
rect 31164 19122 31220 19134
rect 31164 19070 31166 19122
rect 31218 19070 31220 19122
rect 31164 19012 31220 19070
rect 31388 19124 31444 19134
rect 31388 19030 31444 19068
rect 31164 18676 31220 18956
rect 31052 18620 31220 18676
rect 31276 18900 31332 18910
rect 31052 18452 31108 18620
rect 31276 18562 31332 18844
rect 31388 18676 31444 18686
rect 31500 18676 31556 19852
rect 31612 19906 31668 20524
rect 31612 19854 31614 19906
rect 31666 19854 31668 19906
rect 31612 19796 31668 19854
rect 31612 19730 31668 19740
rect 32060 19906 32116 19918
rect 32060 19854 32062 19906
rect 32114 19854 32116 19906
rect 32060 19348 32116 19854
rect 31836 19010 31892 19022
rect 31836 18958 31838 19010
rect 31890 18958 31892 19010
rect 31388 18674 31556 18676
rect 31388 18622 31390 18674
rect 31442 18622 31556 18674
rect 31388 18620 31556 18622
rect 31612 18676 31668 18686
rect 31388 18610 31444 18620
rect 31276 18510 31278 18562
rect 31330 18510 31332 18562
rect 31052 18386 31108 18396
rect 31164 18450 31220 18462
rect 31164 18398 31166 18450
rect 31218 18398 31220 18450
rect 30716 18172 30996 18228
rect 31052 18228 31108 18238
rect 31164 18228 31220 18398
rect 31108 18172 31220 18228
rect 30044 18060 30324 18116
rect 29820 16718 29822 16770
rect 29874 16718 29876 16770
rect 29820 16706 29876 16718
rect 30044 17666 30100 17678
rect 30044 17614 30046 17666
rect 30098 17614 30100 17666
rect 29596 16482 29652 16492
rect 29148 16158 29150 16210
rect 29202 16158 29204 16210
rect 29148 16146 29204 16158
rect 29036 15262 29038 15314
rect 29090 15262 29092 15314
rect 29036 15250 29092 15262
rect 29260 15874 29316 15886
rect 29260 15822 29262 15874
rect 29314 15822 29316 15874
rect 29260 15316 29316 15822
rect 29932 15540 29988 15550
rect 29260 15250 29316 15260
rect 29596 15426 29652 15438
rect 29596 15374 29598 15426
rect 29650 15374 29652 15426
rect 29372 14532 29428 14542
rect 29260 14476 29372 14532
rect 28812 13748 28868 13758
rect 28812 13654 28868 13692
rect 29260 13746 29316 14476
rect 29372 14438 29428 14476
rect 29260 13694 29262 13746
rect 29314 13694 29316 13746
rect 29260 13682 29316 13694
rect 28588 12910 28590 12962
rect 28642 12910 28644 12962
rect 28588 12898 28644 12910
rect 29484 13412 29540 13422
rect 29484 12962 29540 13356
rect 29484 12910 29486 12962
rect 29538 12910 29540 12962
rect 29484 12898 29540 12910
rect 28028 12786 28084 12796
rect 27916 12226 27972 12236
rect 28476 12738 28532 12750
rect 28476 12686 28478 12738
rect 28530 12686 28532 12738
rect 28364 11396 28420 11406
rect 28476 11396 28532 12686
rect 29260 12738 29316 12750
rect 29260 12686 29262 12738
rect 29314 12686 29316 12738
rect 28924 12066 28980 12078
rect 28924 12014 28926 12066
rect 28978 12014 28980 12066
rect 28364 11394 28532 11396
rect 28364 11342 28366 11394
rect 28418 11342 28532 11394
rect 28364 11340 28532 11342
rect 28364 11330 28420 11340
rect 27244 11170 27300 11182
rect 27244 11118 27246 11170
rect 27298 11118 27300 11170
rect 27244 10500 27300 11118
rect 27244 10434 27300 10444
rect 27356 11170 27412 11182
rect 27356 11118 27358 11170
rect 27410 11118 27412 11170
rect 27356 10276 27412 11118
rect 27468 11172 27524 11182
rect 27468 11078 27524 11116
rect 28028 11172 28084 11182
rect 28028 11078 28084 11116
rect 28364 10612 28420 10622
rect 28140 10500 28196 10510
rect 28140 10406 28196 10444
rect 27356 10210 27412 10220
rect 27804 10164 27860 10174
rect 27132 9774 27134 9826
rect 27186 9774 27188 9826
rect 27132 9762 27188 9774
rect 27468 9940 27524 9950
rect 27468 9714 27524 9884
rect 27804 9826 27860 10108
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27804 9762 27860 9774
rect 28140 9826 28196 9838
rect 28140 9774 28142 9826
rect 28194 9774 28196 9826
rect 28140 9716 28196 9774
rect 27468 9662 27470 9714
rect 27522 9662 27524 9714
rect 27468 9650 27524 9662
rect 27916 9660 28140 9716
rect 27132 9268 27188 9278
rect 27020 9212 27132 9268
rect 25900 9156 25956 9166
rect 25900 9062 25956 9100
rect 25788 9042 25844 9054
rect 25788 8990 25790 9042
rect 25842 8990 25844 9042
rect 25788 8428 25844 8990
rect 26460 8930 26516 8942
rect 26460 8878 26462 8930
rect 26514 8878 26516 8930
rect 25564 8372 25620 8382
rect 25564 7474 25620 8316
rect 25564 7422 25566 7474
rect 25618 7422 25620 7474
rect 25564 7410 25620 7422
rect 25676 8372 25844 8428
rect 25900 8818 25956 8830
rect 26348 8820 26404 8830
rect 25900 8766 25902 8818
rect 25954 8766 25956 8818
rect 25676 7364 25732 8372
rect 25676 7270 25732 7308
rect 25788 8036 25844 8046
rect 25452 6750 25454 6802
rect 25506 6750 25508 6802
rect 25452 6692 25508 6750
rect 25452 6626 25508 6636
rect 25452 6020 25508 6030
rect 25452 6018 25732 6020
rect 25452 5966 25454 6018
rect 25506 5966 25732 6018
rect 25452 5964 25732 5966
rect 25452 5954 25508 5964
rect 25564 5794 25620 5806
rect 25564 5742 25566 5794
rect 25618 5742 25620 5794
rect 25564 5460 25620 5742
rect 25004 5404 25620 5460
rect 25004 5234 25060 5404
rect 25004 5182 25006 5234
rect 25058 5182 25060 5234
rect 25004 5170 25060 5182
rect 25228 5236 25284 5246
rect 24556 4510 24558 4562
rect 24610 4510 24612 4562
rect 24556 4498 24612 4510
rect 24668 4452 24724 4462
rect 24668 4358 24724 4396
rect 25228 4450 25284 5180
rect 25228 4398 25230 4450
rect 25282 4398 25284 4450
rect 25228 4386 25284 4398
rect 25676 4452 25732 5964
rect 25788 6018 25844 7980
rect 25788 5966 25790 6018
rect 25842 5966 25844 6018
rect 25788 5954 25844 5966
rect 25900 5906 25956 8766
rect 26124 8818 26404 8820
rect 26124 8766 26350 8818
rect 26402 8766 26404 8818
rect 26124 8764 26404 8766
rect 26124 7812 26180 8764
rect 26348 8754 26404 8764
rect 26460 8428 26516 8878
rect 27020 8428 27076 9212
rect 27132 9174 27188 9212
rect 27916 8930 27972 9660
rect 28140 9650 28196 9660
rect 28364 9266 28420 10556
rect 28476 9828 28532 11340
rect 28588 11396 28644 11406
rect 28588 11302 28644 11340
rect 28812 11172 28868 11182
rect 28812 10722 28868 11116
rect 28924 10836 28980 12014
rect 29260 11732 29316 12686
rect 29260 11666 29316 11676
rect 29372 12738 29428 12750
rect 29372 12686 29374 12738
rect 29426 12686 29428 12738
rect 29372 11508 29428 12686
rect 29372 11442 29428 11452
rect 29484 11732 29540 11742
rect 28924 10770 28980 10780
rect 29148 11394 29204 11406
rect 29148 11342 29150 11394
rect 29202 11342 29204 11394
rect 28812 10670 28814 10722
rect 28866 10670 28868 10722
rect 28812 10658 28868 10670
rect 29148 10724 29204 11342
rect 29148 10164 29204 10668
rect 29372 10612 29428 10622
rect 29484 10612 29540 11676
rect 29428 10556 29540 10612
rect 29596 11394 29652 15374
rect 29932 14644 29988 15484
rect 30044 15148 30100 17614
rect 30268 17332 30324 18060
rect 30716 17778 30772 18172
rect 31052 18162 31108 18172
rect 31276 17892 31332 18510
rect 31500 18452 31556 18462
rect 31612 18452 31668 18620
rect 31500 18450 31668 18452
rect 31500 18398 31502 18450
rect 31554 18398 31668 18450
rect 31500 18396 31668 18398
rect 31724 18450 31780 18462
rect 31724 18398 31726 18450
rect 31778 18398 31780 18450
rect 31500 18386 31556 18396
rect 31276 17826 31332 17836
rect 30716 17726 30718 17778
rect 30770 17726 30772 17778
rect 30716 17714 30772 17726
rect 31724 17780 31780 18398
rect 31836 18228 31892 18958
rect 32060 18788 32116 19292
rect 32508 19906 32564 21532
rect 33180 21474 33236 21486
rect 33180 21422 33182 21474
rect 33234 21422 33236 21474
rect 33180 21028 33236 21422
rect 32844 20972 33236 21028
rect 32844 20914 32900 20972
rect 32844 20862 32846 20914
rect 32898 20862 32900 20914
rect 32844 20850 32900 20862
rect 32508 19854 32510 19906
rect 32562 19854 32564 19906
rect 32172 19012 32228 19022
rect 32172 18918 32228 18956
rect 32060 18722 32116 18732
rect 31948 18676 32004 18686
rect 31948 18564 32004 18620
rect 32060 18564 32116 18574
rect 31948 18562 32116 18564
rect 31948 18510 32062 18562
rect 32114 18510 32116 18562
rect 31948 18508 32116 18510
rect 32060 18498 32116 18508
rect 32508 18564 32564 19854
rect 32620 20356 32676 20366
rect 32620 19236 32676 20300
rect 33180 19908 33236 19918
rect 33180 19796 33236 19852
rect 32620 19142 32676 19180
rect 32956 19740 33236 19796
rect 32844 18900 32900 18910
rect 32956 18900 33012 19740
rect 33516 19460 33572 22876
rect 33628 22820 33684 22830
rect 33628 22594 33684 22764
rect 33628 22542 33630 22594
rect 33682 22542 33684 22594
rect 33628 22530 33684 22542
rect 33964 22370 34020 23212
rect 34076 23156 34132 27468
rect 34188 24612 34244 30940
rect 34524 30996 34580 31006
rect 34636 30996 34692 33964
rect 35196 33908 35252 35084
rect 35420 35028 35476 35038
rect 35532 35028 35588 35084
rect 35420 35026 35588 35028
rect 35420 34974 35422 35026
rect 35474 34974 35588 35026
rect 35420 34972 35588 34974
rect 35644 36708 35700 36718
rect 35420 34962 35476 34972
rect 35644 34018 35700 36652
rect 36428 36596 36484 36606
rect 36092 36594 36484 36596
rect 36092 36542 36430 36594
rect 36482 36542 36484 36594
rect 36092 36540 36484 36542
rect 35980 36484 36036 36494
rect 35980 34690 36036 36428
rect 36092 35028 36148 36540
rect 36428 36530 36484 36540
rect 36652 36484 36708 38782
rect 36764 38724 36820 38734
rect 36876 38724 36932 41020
rect 36988 41010 37044 41020
rect 37100 40964 37156 41358
rect 37100 40898 37156 40908
rect 37212 40740 37268 41916
rect 37436 41970 37492 42028
rect 37436 41918 37438 41970
rect 37490 41918 37492 41970
rect 37436 41906 37492 41918
rect 37100 40684 37268 40740
rect 37548 40740 37604 42252
rect 37660 42196 37716 42206
rect 37660 41074 37716 42140
rect 37884 41748 37940 46510
rect 38332 46562 38388 46574
rect 38332 46510 38334 46562
rect 38386 46510 38388 46562
rect 37996 46450 38052 46462
rect 37996 46398 37998 46450
rect 38050 46398 38052 46450
rect 37996 45220 38052 46398
rect 38108 45220 38164 45230
rect 37996 45218 38164 45220
rect 37996 45166 38110 45218
rect 38162 45166 38164 45218
rect 37996 45164 38164 45166
rect 38108 45154 38164 45164
rect 38332 44660 38388 46510
rect 38444 46450 38500 46462
rect 38444 46398 38446 46450
rect 38498 46398 38500 46450
rect 38444 46002 38500 46398
rect 38668 46450 38724 47068
rect 38892 46788 38948 47180
rect 39228 47170 39284 47180
rect 40348 47236 40404 47246
rect 38668 46398 38670 46450
rect 38722 46398 38724 46450
rect 38668 46386 38724 46398
rect 38780 46732 38948 46788
rect 38444 45950 38446 46002
rect 38498 45950 38500 46002
rect 38444 45938 38500 45950
rect 38332 44594 38388 44604
rect 38332 44436 38388 44446
rect 38332 44342 38388 44380
rect 38332 43540 38388 43550
rect 38220 43426 38276 43438
rect 38220 43374 38222 43426
rect 38274 43374 38276 43426
rect 37884 41682 37940 41692
rect 38108 43204 38164 43214
rect 38108 41972 38164 43148
rect 37660 41022 37662 41074
rect 37714 41022 37716 41074
rect 37660 41010 37716 41022
rect 36988 40180 37044 40190
rect 36988 39618 37044 40124
rect 36988 39566 36990 39618
rect 37042 39566 37044 39618
rect 36988 39554 37044 39566
rect 36820 38668 36932 38724
rect 37100 38668 37156 40684
rect 37324 40404 37380 40414
rect 37324 40310 37380 40348
rect 37212 39620 37268 39630
rect 37212 39526 37268 39564
rect 37436 39620 37492 39630
rect 37548 39620 37604 40684
rect 37996 40962 38052 40974
rect 37996 40910 37998 40962
rect 38050 40910 38052 40962
rect 37884 40404 37940 40414
rect 37436 39618 37548 39620
rect 37436 39566 37438 39618
rect 37490 39566 37548 39618
rect 37436 39564 37548 39566
rect 37436 39554 37492 39564
rect 37548 39526 37604 39564
rect 37660 39618 37716 39630
rect 37660 39566 37662 39618
rect 37714 39566 37716 39618
rect 37324 39508 37380 39518
rect 37324 39414 37380 39452
rect 37660 39172 37716 39566
rect 37660 39106 37716 39116
rect 37548 39060 37604 39070
rect 36764 38658 36820 38668
rect 37100 38612 37268 38668
rect 36652 36418 36708 36428
rect 36876 38276 36932 38286
rect 36876 37380 36932 38220
rect 36988 38164 37044 38174
rect 36988 38070 37044 38108
rect 36092 35026 36260 35028
rect 36092 34974 36094 35026
rect 36146 34974 36260 35026
rect 36092 34972 36260 34974
rect 36092 34962 36148 34972
rect 35980 34638 35982 34690
rect 36034 34638 36036 34690
rect 35980 34626 36036 34638
rect 36204 34242 36260 34972
rect 36204 34190 36206 34242
rect 36258 34190 36260 34242
rect 36204 34178 36260 34190
rect 35644 33966 35646 34018
rect 35698 33966 35700 34018
rect 35644 33954 35700 33966
rect 35084 33852 35252 33908
rect 35084 33572 35140 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35084 33506 35140 33516
rect 34748 33460 34804 33470
rect 34748 32674 34804 33404
rect 34748 32622 34750 32674
rect 34802 32622 34804 32674
rect 34748 32610 34804 32622
rect 36428 33460 36484 33470
rect 36204 32452 36260 32462
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 31890 35252 31902
rect 35196 31838 35198 31890
rect 35250 31838 35252 31890
rect 35196 31668 35252 31838
rect 35868 31892 35924 31902
rect 35868 31798 35924 31836
rect 35980 31780 36036 31790
rect 35980 31686 36036 31724
rect 35532 31668 35588 31678
rect 35196 31666 35588 31668
rect 35196 31614 35534 31666
rect 35586 31614 35588 31666
rect 35196 31612 35588 31614
rect 34580 30940 34692 30996
rect 34748 31444 34804 31454
rect 34748 31218 34804 31388
rect 34748 31166 34750 31218
rect 34802 31166 34804 31218
rect 34524 30930 34580 30940
rect 34412 30772 34468 30782
rect 34412 29426 34468 30716
rect 34748 29650 34804 31166
rect 35084 31332 35140 31342
rect 34860 29764 34916 29774
rect 34916 29708 35028 29764
rect 34860 29698 34916 29708
rect 34748 29598 34750 29650
rect 34802 29598 34804 29650
rect 34748 29586 34804 29598
rect 34972 29650 35028 29708
rect 34972 29598 34974 29650
rect 35026 29598 35028 29650
rect 34972 29586 35028 29598
rect 35084 29650 35140 31276
rect 35196 30772 35252 31612
rect 35532 31602 35588 31612
rect 35756 31554 35812 31566
rect 35756 31502 35758 31554
rect 35810 31502 35812 31554
rect 35756 31332 35812 31502
rect 36092 31554 36148 31566
rect 36092 31502 36094 31554
rect 36146 31502 36148 31554
rect 36092 31444 36148 31502
rect 36092 31378 36148 31388
rect 35756 31266 35812 31276
rect 35308 30996 35364 31006
rect 35308 30902 35364 30940
rect 35196 30706 35252 30716
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 30212 35252 30222
rect 35196 30118 35252 30156
rect 35980 30212 36036 30222
rect 36204 30212 36260 32396
rect 36428 31780 36484 33404
rect 36428 31724 36820 31780
rect 35980 30210 36260 30212
rect 35980 30158 35982 30210
rect 36034 30158 36260 30210
rect 35980 30156 36260 30158
rect 36316 31556 36372 31566
rect 36316 30210 36372 31500
rect 36652 31108 36708 31118
rect 36316 30158 36318 30210
rect 36370 30158 36372 30210
rect 35980 30146 36036 30156
rect 36316 30146 36372 30158
rect 36540 30548 36596 30558
rect 36428 30100 36484 30110
rect 36428 30006 36484 30044
rect 35084 29598 35086 29650
rect 35138 29598 35140 29650
rect 35084 29586 35140 29598
rect 36428 29652 36484 29662
rect 36428 29558 36484 29596
rect 36540 29650 36596 30492
rect 36540 29598 36542 29650
rect 36594 29598 36596 29650
rect 36540 29586 36596 29598
rect 34860 29540 34916 29550
rect 34860 29446 34916 29484
rect 36652 29538 36708 31052
rect 36652 29486 36654 29538
rect 36706 29486 36708 29538
rect 34412 29374 34414 29426
rect 34466 29374 34468 29426
rect 34412 29362 34468 29374
rect 35196 29428 35252 29438
rect 35196 29334 35252 29372
rect 35980 29428 36036 29438
rect 35980 29426 36260 29428
rect 35980 29374 35982 29426
rect 36034 29374 36260 29426
rect 35980 29372 36260 29374
rect 35980 29362 36036 29372
rect 35756 29316 35812 29326
rect 35644 29202 35700 29214
rect 35644 29150 35646 29202
rect 35698 29150 35700 29202
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34636 28868 34692 28878
rect 34412 27860 34468 27870
rect 34412 27766 34468 27804
rect 34636 27858 34692 28812
rect 35308 28756 35364 28766
rect 35084 28700 35308 28756
rect 35084 27860 35140 28700
rect 35308 28662 35364 28700
rect 34636 27806 34638 27858
rect 34690 27806 34692 27858
rect 34636 27794 34692 27806
rect 34748 27858 35140 27860
rect 34748 27806 35086 27858
rect 35138 27806 35140 27858
rect 34748 27804 35140 27806
rect 34748 26908 34804 27804
rect 35084 27794 35140 27804
rect 35644 27972 35700 29150
rect 35756 28866 35812 29260
rect 35980 29204 36036 29214
rect 35980 29110 36036 29148
rect 35756 28814 35758 28866
rect 35810 28814 35812 28866
rect 35756 28802 35812 28814
rect 35980 28756 36036 28766
rect 36036 28700 36148 28756
rect 35980 28690 36036 28700
rect 35868 28644 35924 28654
rect 35868 28550 35924 28588
rect 36092 28642 36148 28700
rect 36092 28590 36094 28642
rect 36146 28590 36148 28642
rect 36092 28578 36148 28590
rect 35196 27468 35460 27478
rect 34524 26852 34804 26908
rect 34860 27412 34916 27422
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34300 25506 34356 25518
rect 34300 25454 34302 25506
rect 34354 25454 34356 25506
rect 34300 25396 34356 25454
rect 34524 25508 34580 26852
rect 34524 25414 34580 25452
rect 34636 26292 34692 26302
rect 34636 25506 34692 26236
rect 34636 25454 34638 25506
rect 34690 25454 34692 25506
rect 34636 25442 34692 25454
rect 34300 25330 34356 25340
rect 34860 25172 34916 27356
rect 35644 27076 35700 27916
rect 35756 28532 35812 28542
rect 35756 28082 35812 28476
rect 35756 28030 35758 28082
rect 35810 28030 35812 28082
rect 35756 27188 35812 28030
rect 36204 27972 36260 29372
rect 36204 27906 36260 27916
rect 36540 27858 36596 27870
rect 36540 27806 36542 27858
rect 36594 27806 36596 27858
rect 35756 27122 35812 27132
rect 36204 27748 36260 27758
rect 35644 27010 35700 27020
rect 36204 27074 36260 27692
rect 36204 27022 36206 27074
rect 36258 27022 36260 27074
rect 36204 27010 36260 27022
rect 36316 27748 36372 27758
rect 36540 27748 36596 27806
rect 36316 27746 36596 27748
rect 36316 27694 36318 27746
rect 36370 27694 36596 27746
rect 36316 27692 36596 27694
rect 36316 26404 36372 27692
rect 36652 26908 36708 29486
rect 36764 29426 36820 31724
rect 36764 29374 36766 29426
rect 36818 29374 36820 29426
rect 36764 29362 36820 29374
rect 36876 27858 36932 37324
rect 37100 37826 37156 37838
rect 37100 37774 37102 37826
rect 37154 37774 37156 37826
rect 37100 37378 37156 37774
rect 37100 37326 37102 37378
rect 37154 37326 37156 37378
rect 37100 37314 37156 37326
rect 36988 35700 37044 35710
rect 36988 35606 37044 35644
rect 37212 35140 37268 38612
rect 37548 38162 37604 39004
rect 37884 38500 37940 40348
rect 37884 38434 37940 38444
rect 37996 39618 38052 40910
rect 38108 40404 38164 41916
rect 38220 41860 38276 43374
rect 38332 42754 38388 43484
rect 38332 42702 38334 42754
rect 38386 42702 38388 42754
rect 38332 42196 38388 42702
rect 38668 43204 38724 43214
rect 38668 42756 38724 43148
rect 38780 42980 38836 46732
rect 38780 42914 38836 42924
rect 38892 46562 38948 46574
rect 39340 46564 39396 46574
rect 39788 46564 39844 46574
rect 38892 46510 38894 46562
rect 38946 46510 38948 46562
rect 38892 46450 38948 46510
rect 38892 46398 38894 46450
rect 38946 46398 38948 46450
rect 38780 42756 38836 42766
rect 38668 42754 38836 42756
rect 38668 42702 38782 42754
rect 38834 42702 38836 42754
rect 38668 42700 38836 42702
rect 38780 42690 38836 42700
rect 38444 42530 38500 42542
rect 38444 42478 38446 42530
rect 38498 42478 38500 42530
rect 38444 42420 38500 42478
rect 38556 42532 38612 42542
rect 38556 42438 38612 42476
rect 38668 42530 38724 42542
rect 38668 42478 38670 42530
rect 38722 42478 38724 42530
rect 38444 42354 38500 42364
rect 38556 42196 38612 42206
rect 38332 42194 38612 42196
rect 38332 42142 38558 42194
rect 38610 42142 38612 42194
rect 38332 42140 38612 42142
rect 38220 41794 38276 41804
rect 38444 41972 38500 41982
rect 38444 41300 38500 41916
rect 38556 41636 38612 42140
rect 38668 42196 38724 42478
rect 38668 42130 38724 42140
rect 38892 41972 38948 46398
rect 38556 41570 38612 41580
rect 38668 41970 38948 41972
rect 38668 41918 38894 41970
rect 38946 41918 38948 41970
rect 38668 41916 38948 41918
rect 38556 41300 38612 41310
rect 38444 41298 38612 41300
rect 38444 41246 38558 41298
rect 38610 41246 38612 41298
rect 38444 41244 38612 41246
rect 38556 41234 38612 41244
rect 38108 40310 38164 40348
rect 38220 40852 38276 40862
rect 37996 39566 37998 39618
rect 38050 39566 38052 39618
rect 37548 38110 37550 38162
rect 37602 38110 37604 38162
rect 37548 38098 37604 38110
rect 37660 38388 37716 38398
rect 37548 36482 37604 36494
rect 37548 36430 37550 36482
rect 37602 36430 37604 36482
rect 37324 36372 37380 36382
rect 37324 36278 37380 36316
rect 37548 35812 37604 36430
rect 37548 35746 37604 35756
rect 37212 35074 37268 35084
rect 37548 35588 37604 35598
rect 37324 35028 37380 35038
rect 37324 34934 37380 34972
rect 37436 34244 37492 34254
rect 37436 34150 37492 34188
rect 36988 34130 37044 34142
rect 36988 34078 36990 34130
rect 37042 34078 37044 34130
rect 36988 34020 37044 34078
rect 36988 33954 37044 33964
rect 36988 33346 37044 33358
rect 36988 33294 36990 33346
rect 37042 33294 37044 33346
rect 36988 32452 37044 33294
rect 37548 32564 37604 35532
rect 37548 32498 37604 32508
rect 36988 32386 37044 32396
rect 37324 31668 37380 31678
rect 37324 31574 37380 31612
rect 37212 31554 37268 31566
rect 37212 31502 37214 31554
rect 37266 31502 37268 31554
rect 37212 31108 37268 31502
rect 37436 31556 37492 31566
rect 37436 31462 37492 31500
rect 37548 31554 37604 31566
rect 37548 31502 37550 31554
rect 37602 31502 37604 31554
rect 37212 31042 37268 31052
rect 37548 30548 37604 31502
rect 37548 30482 37604 30492
rect 36988 30322 37044 30334
rect 36988 30270 36990 30322
rect 37042 30270 37044 30322
rect 36988 29764 37044 30270
rect 37660 29988 37716 38332
rect 37884 36260 37940 36270
rect 37884 36166 37940 36204
rect 37996 35924 38052 39566
rect 38108 38836 38164 38846
rect 38220 38836 38276 40796
rect 38668 40628 38724 41916
rect 38892 41906 38948 41916
rect 39004 46562 39396 46564
rect 39004 46510 39342 46562
rect 39394 46510 39396 46562
rect 39004 46508 39396 46510
rect 39004 41188 39060 46508
rect 39340 46498 39396 46508
rect 39452 46562 39844 46564
rect 39452 46510 39790 46562
rect 39842 46510 39844 46562
rect 39452 46508 39844 46510
rect 39228 42754 39284 42766
rect 39228 42702 39230 42754
rect 39282 42702 39284 42754
rect 39116 42644 39172 42654
rect 39116 41412 39172 42588
rect 39228 41972 39284 42702
rect 39452 42194 39508 46508
rect 39788 46498 39844 46508
rect 40236 44996 40292 45006
rect 39900 44994 40292 44996
rect 39900 44942 40238 44994
rect 40290 44942 40292 44994
rect 39900 44940 40292 44942
rect 39900 44212 39956 44940
rect 40236 44930 40292 44940
rect 39452 42142 39454 42194
rect 39506 42142 39508 42194
rect 39228 41906 39284 41916
rect 39340 41970 39396 41982
rect 39340 41918 39342 41970
rect 39394 41918 39396 41970
rect 39340 41636 39396 41918
rect 39452 41636 39508 42142
rect 39676 42196 39732 42206
rect 39676 42102 39732 42140
rect 39900 42082 39956 44156
rect 40348 43652 40404 47180
rect 41020 47236 41076 47246
rect 41020 47142 41076 47180
rect 41020 46676 41076 46686
rect 41020 46582 41076 46620
rect 40460 46562 40516 46574
rect 40460 46510 40462 46562
rect 40514 46510 40516 46562
rect 40460 44660 40516 46510
rect 41244 46114 41300 47404
rect 41916 47460 41972 47470
rect 41916 47366 41972 47404
rect 42140 47460 42196 47470
rect 42140 47366 42196 47404
rect 41580 47346 41636 47358
rect 41580 47294 41582 47346
rect 41634 47294 41636 47346
rect 41356 47236 41412 47246
rect 41356 47142 41412 47180
rect 41468 47234 41524 47246
rect 41468 47182 41470 47234
rect 41522 47182 41524 47234
rect 41244 46062 41246 46114
rect 41298 46062 41300 46114
rect 41244 46050 41300 46062
rect 41356 46676 41412 46686
rect 40572 46004 40628 46014
rect 40572 46002 41188 46004
rect 40572 45950 40574 46002
rect 40626 45950 41188 46002
rect 40572 45948 41188 45950
rect 40572 45938 40628 45948
rect 41132 45220 41188 45948
rect 41244 45220 41300 45230
rect 41132 45218 41300 45220
rect 41132 45166 41246 45218
rect 41298 45166 41300 45218
rect 41132 45164 41300 45166
rect 41356 45220 41412 46620
rect 41468 45444 41524 47182
rect 41580 46116 41636 47294
rect 42028 47236 42084 47246
rect 41692 47234 42084 47236
rect 41692 47182 42030 47234
rect 42082 47182 42084 47234
rect 41692 47180 42084 47182
rect 41692 46786 41748 47180
rect 42028 47170 42084 47180
rect 41692 46734 41694 46786
rect 41746 46734 41748 46786
rect 41692 46722 41748 46734
rect 41580 46050 41636 46060
rect 41692 46228 41748 46238
rect 41580 45892 41636 45902
rect 41692 45892 41748 46172
rect 41580 45890 41748 45892
rect 41580 45838 41582 45890
rect 41634 45838 41748 45890
rect 41580 45836 41748 45838
rect 41580 45826 41636 45836
rect 41468 45378 41524 45388
rect 41356 45164 41524 45220
rect 40460 44604 40628 44660
rect 40460 44434 40516 44446
rect 40460 44382 40462 44434
rect 40514 44382 40516 44434
rect 40460 44100 40516 44382
rect 40572 44324 40628 44604
rect 41132 44436 41188 44474
rect 41132 44370 41188 44380
rect 41020 44324 41076 44334
rect 40572 44322 41076 44324
rect 40572 44270 41022 44322
rect 41074 44270 41076 44322
rect 40572 44268 41076 44270
rect 41244 44324 41300 45164
rect 41356 44996 41412 45006
rect 41356 44902 41412 44940
rect 41356 44324 41412 44334
rect 41244 44322 41412 44324
rect 41244 44270 41358 44322
rect 41410 44270 41412 44322
rect 41244 44268 41412 44270
rect 40460 44034 40516 44044
rect 40348 43596 40516 43652
rect 40348 43426 40404 43438
rect 40348 43374 40350 43426
rect 40402 43374 40404 43426
rect 40348 43204 40404 43374
rect 40348 43138 40404 43148
rect 39900 42030 39902 42082
rect 39954 42030 39956 42082
rect 39900 42018 39956 42030
rect 40012 42642 40068 42654
rect 40012 42590 40014 42642
rect 40066 42590 40068 42642
rect 39564 41860 39620 41870
rect 39564 41858 39732 41860
rect 39564 41806 39566 41858
rect 39618 41806 39732 41858
rect 39564 41804 39732 41806
rect 39564 41794 39620 41804
rect 39676 41748 39732 41804
rect 39676 41682 39732 41692
rect 39452 41580 39620 41636
rect 39340 41570 39396 41580
rect 39116 41356 39396 41412
rect 38668 39618 38724 40572
rect 38668 39566 38670 39618
rect 38722 39566 38724 39618
rect 38332 39396 38388 39406
rect 38388 39340 38500 39396
rect 38332 39302 38388 39340
rect 38108 38834 38276 38836
rect 38108 38782 38110 38834
rect 38162 38782 38276 38834
rect 38108 38780 38276 38782
rect 38332 39060 38388 39070
rect 38108 38770 38164 38780
rect 38332 36482 38388 39004
rect 38332 36430 38334 36482
rect 38386 36430 38388 36482
rect 38332 36418 38388 36430
rect 38444 37268 38500 39340
rect 38668 38836 38724 39566
rect 38444 36482 38500 37212
rect 38444 36430 38446 36482
rect 38498 36430 38500 36482
rect 38444 36418 38500 36430
rect 38556 38780 38724 38836
rect 38780 40964 38836 40974
rect 38780 38834 38836 40908
rect 39004 40626 39060 41132
rect 39004 40574 39006 40626
rect 39058 40574 39060 40626
rect 39004 40562 39060 40574
rect 38892 40404 38948 40414
rect 38892 40402 39060 40404
rect 38892 40350 38894 40402
rect 38946 40350 39060 40402
rect 38892 40348 39060 40350
rect 38892 40338 38948 40348
rect 38780 38782 38782 38834
rect 38834 38782 38836 38834
rect 38556 36260 38612 38780
rect 38780 38770 38836 38782
rect 38892 39508 38948 39518
rect 38892 38836 38948 39452
rect 38892 38770 38948 38780
rect 39004 39394 39060 40348
rect 39228 40402 39284 40414
rect 39228 40350 39230 40402
rect 39282 40350 39284 40402
rect 39004 39342 39006 39394
rect 39058 39342 39060 39394
rect 39004 39284 39060 39342
rect 38892 38612 38948 38622
rect 38892 37940 38948 38556
rect 38668 37884 38892 37940
rect 38668 36482 38724 37884
rect 38892 37874 38948 37884
rect 38892 37716 38948 37726
rect 38780 37660 38892 37716
rect 38780 36594 38836 37660
rect 38892 37650 38948 37660
rect 39004 37492 39060 39228
rect 39116 40290 39172 40302
rect 39116 40238 39118 40290
rect 39170 40238 39172 40290
rect 39116 38724 39172 40238
rect 39228 39732 39284 40350
rect 39228 39396 39284 39676
rect 39228 39330 39284 39340
rect 39116 38658 39172 38668
rect 39228 38948 39284 38958
rect 38780 36542 38782 36594
rect 38834 36542 38836 36594
rect 38780 36530 38836 36542
rect 38892 37436 39004 37492
rect 38668 36430 38670 36482
rect 38722 36430 38724 36482
rect 38668 36418 38724 36430
rect 38892 36482 38948 37436
rect 39004 37426 39060 37436
rect 39228 37154 39284 38892
rect 39228 37102 39230 37154
rect 39282 37102 39284 37154
rect 39228 37090 39284 37102
rect 38892 36430 38894 36482
rect 38946 36430 38948 36482
rect 38892 36418 38948 36430
rect 38556 36204 38836 36260
rect 37996 35858 38052 35868
rect 38668 35812 38724 35822
rect 38668 35718 38724 35756
rect 38556 35700 38612 35710
rect 38108 34804 38164 34814
rect 38108 34020 38164 34748
rect 38444 34020 38500 34030
rect 38108 34018 38500 34020
rect 38108 33966 38446 34018
rect 38498 33966 38500 34018
rect 38108 33964 38500 33966
rect 37772 33236 37828 33246
rect 37772 33142 37828 33180
rect 37996 33012 38052 33022
rect 37884 32956 37996 33012
rect 37660 29922 37716 29932
rect 37772 31666 37828 31678
rect 37772 31614 37774 31666
rect 37826 31614 37828 31666
rect 36988 29698 37044 29708
rect 37660 29764 37716 29774
rect 37660 29428 37716 29708
rect 37772 29428 37828 31614
rect 37884 30212 37940 32956
rect 37996 32946 38052 32956
rect 37884 30146 37940 30156
rect 37996 32564 38052 32574
rect 37996 31106 38052 32508
rect 37996 31054 37998 31106
rect 38050 31054 38052 31106
rect 37660 29426 37828 29428
rect 37660 29374 37662 29426
rect 37714 29374 37828 29426
rect 37660 29372 37828 29374
rect 37660 29362 37716 29372
rect 36988 29314 37044 29326
rect 36988 29262 36990 29314
rect 37042 29262 37044 29314
rect 36988 28530 37044 29262
rect 36988 28478 36990 28530
rect 37042 28478 37044 28530
rect 36988 28466 37044 28478
rect 37324 28642 37380 28654
rect 37324 28590 37326 28642
rect 37378 28590 37380 28642
rect 36876 27806 36878 27858
rect 36930 27806 36932 27858
rect 36876 27794 36932 27806
rect 36988 27972 37044 27982
rect 36988 27412 37044 27916
rect 36988 27356 37156 27412
rect 36988 27076 37044 27114
rect 36988 27010 37044 27020
rect 37100 26962 37156 27356
rect 37324 27074 37380 28590
rect 37324 27022 37326 27074
rect 37378 27022 37380 27074
rect 37324 27010 37380 27022
rect 37436 28532 37492 28542
rect 37100 26910 37102 26962
rect 37154 26910 37156 26962
rect 37100 26908 37156 26910
rect 37436 26908 37492 28476
rect 36204 26348 36372 26404
rect 36540 26852 36708 26908
rect 36988 26852 37156 26908
rect 37324 26852 37492 26908
rect 37548 27636 37604 27646
rect 35980 26290 36036 26302
rect 35980 26238 35982 26290
rect 36034 26238 36036 26290
rect 35196 26180 35252 26190
rect 35084 26178 35252 26180
rect 35084 26126 35198 26178
rect 35250 26126 35252 26178
rect 35084 26124 35252 26126
rect 35084 25620 35140 26124
rect 35196 26114 35252 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35532 25620 35588 25630
rect 35084 25564 35252 25620
rect 34972 25508 35028 25518
rect 35028 25452 35140 25508
rect 34972 25442 35028 25452
rect 35084 25394 35140 25452
rect 35084 25342 35086 25394
rect 35138 25342 35140 25394
rect 35084 25330 35140 25342
rect 35196 25284 35252 25564
rect 35532 25526 35588 25564
rect 35644 25508 35700 25518
rect 35644 25414 35700 25452
rect 35868 25506 35924 25518
rect 35868 25454 35870 25506
rect 35922 25454 35924 25506
rect 35532 25284 35588 25294
rect 35196 25282 35588 25284
rect 35196 25230 35534 25282
rect 35586 25230 35588 25282
rect 35196 25228 35588 25230
rect 35532 25218 35588 25228
rect 34860 25116 35140 25172
rect 34188 23380 34244 24556
rect 34860 24164 34916 24174
rect 34860 24070 34916 24108
rect 34412 23940 34468 23950
rect 34972 23940 35028 23950
rect 34412 23938 34692 23940
rect 34412 23886 34414 23938
rect 34466 23886 34692 23938
rect 34412 23884 34692 23886
rect 34412 23874 34468 23884
rect 34524 23714 34580 23726
rect 34524 23662 34526 23714
rect 34578 23662 34580 23714
rect 34412 23492 34468 23502
rect 34188 23324 34356 23380
rect 34188 23156 34244 23166
rect 34076 23154 34244 23156
rect 34076 23102 34190 23154
rect 34242 23102 34244 23154
rect 34076 23100 34244 23102
rect 34188 23090 34244 23100
rect 34188 22932 34244 22942
rect 33964 22318 33966 22370
rect 34018 22318 34020 22370
rect 33964 21924 34020 22318
rect 33964 21858 34020 21868
rect 34076 22876 34188 22932
rect 34076 21810 34132 22876
rect 34188 22866 34244 22876
rect 34188 22372 34244 22382
rect 34188 21924 34244 22316
rect 34188 21858 34244 21868
rect 34076 21758 34078 21810
rect 34130 21758 34132 21810
rect 34076 21746 34132 21758
rect 33740 21586 33796 21598
rect 34188 21588 34244 21598
rect 33740 21534 33742 21586
rect 33794 21534 33796 21586
rect 33740 21476 33796 21534
rect 33964 21586 34244 21588
rect 33964 21534 34190 21586
rect 34242 21534 34244 21586
rect 33964 21532 34244 21534
rect 33852 21476 33908 21486
rect 33740 21420 33852 21476
rect 33852 21410 33908 21420
rect 33516 19394 33572 19404
rect 33628 20802 33684 20814
rect 33628 20750 33630 20802
rect 33682 20750 33684 20802
rect 33628 20692 33684 20750
rect 33628 19236 33684 20636
rect 33852 20578 33908 20590
rect 33852 20526 33854 20578
rect 33906 20526 33908 20578
rect 33852 20244 33908 20526
rect 33964 20580 34020 21532
rect 34188 21522 34244 21532
rect 34076 21364 34132 21374
rect 34076 21270 34132 21308
rect 34188 21140 34244 21150
rect 34188 20802 34244 21084
rect 34188 20750 34190 20802
rect 34242 20750 34244 20802
rect 34188 20738 34244 20750
rect 34076 20580 34132 20590
rect 33964 20578 34132 20580
rect 33964 20526 34078 20578
rect 34130 20526 34132 20578
rect 33964 20524 34132 20526
rect 33852 20178 33908 20188
rect 33292 19234 33684 19236
rect 33292 19182 33630 19234
rect 33682 19182 33684 19234
rect 33292 19180 33684 19182
rect 32900 18844 33012 18900
rect 33068 19122 33124 19134
rect 33068 19070 33070 19122
rect 33122 19070 33124 19122
rect 32844 18834 32900 18844
rect 32508 18498 32564 18508
rect 31836 18162 31892 18172
rect 32284 18450 32340 18462
rect 32284 18398 32286 18450
rect 32338 18398 32340 18450
rect 31724 17714 31780 17724
rect 30268 16996 30324 17276
rect 32284 17556 32340 18398
rect 32844 17780 32900 17790
rect 33068 17780 33124 19070
rect 33180 19010 33236 19022
rect 33180 18958 33182 19010
rect 33234 18958 33236 19010
rect 33180 18452 33236 18958
rect 33180 18386 33236 18396
rect 33292 18450 33348 19180
rect 33628 19170 33684 19180
rect 33852 19794 33908 19806
rect 33852 19742 33854 19794
rect 33906 19742 33908 19794
rect 33292 18398 33294 18450
rect 33346 18398 33348 18450
rect 33292 18386 33348 18398
rect 33852 19012 33908 19742
rect 34076 19012 34132 20524
rect 34300 20580 34356 23324
rect 34412 22708 34468 23436
rect 34524 23380 34580 23662
rect 34524 23314 34580 23324
rect 34524 22932 34580 22942
rect 34524 22838 34580 22876
rect 34412 22652 34580 22708
rect 34300 20514 34356 20524
rect 34412 21026 34468 21038
rect 34412 20974 34414 21026
rect 34466 20974 34468 21026
rect 34300 20244 34356 20254
rect 34188 20020 34244 20030
rect 34188 19926 34244 19964
rect 34300 19346 34356 20188
rect 34412 20018 34468 20974
rect 34412 19966 34414 20018
rect 34466 19966 34468 20018
rect 34412 19954 34468 19966
rect 34524 20020 34580 22652
rect 34636 22484 34692 23884
rect 34972 23846 35028 23884
rect 35084 23548 35140 25116
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 23940 35252 23950
rect 35196 23846 35252 23884
rect 35420 23938 35476 23950
rect 35420 23886 35422 23938
rect 35474 23886 35476 23938
rect 35420 23604 35476 23886
rect 35868 23828 35924 25454
rect 35980 25172 36036 26238
rect 36204 26068 36260 26348
rect 36204 26002 36260 26012
rect 36316 26178 36372 26190
rect 36316 26126 36318 26178
rect 36370 26126 36372 26178
rect 36316 25506 36372 26126
rect 36316 25454 36318 25506
rect 36370 25454 36372 25506
rect 36316 25442 36372 25454
rect 36428 25396 36484 25406
rect 36428 25302 36484 25340
rect 35980 25106 36036 25116
rect 36316 25284 36372 25294
rect 36316 24724 36372 25228
rect 35980 24722 36372 24724
rect 35980 24670 36318 24722
rect 36370 24670 36372 24722
rect 35980 24668 36372 24670
rect 35980 24610 36036 24668
rect 36316 24658 36372 24668
rect 35980 24558 35982 24610
rect 36034 24558 36036 24610
rect 35980 24546 36036 24558
rect 36428 24612 36484 24622
rect 36316 24500 36372 24510
rect 36204 24498 36372 24500
rect 36204 24446 36318 24498
rect 36370 24446 36372 24498
rect 36204 24444 36372 24446
rect 36092 24052 36148 24062
rect 36092 23958 36148 23996
rect 35868 23762 35924 23772
rect 36204 23604 36260 24444
rect 36316 24434 36372 24444
rect 36428 24050 36484 24556
rect 36428 23998 36430 24050
rect 36482 23998 36484 24050
rect 36428 23986 36484 23998
rect 35420 23548 36260 23604
rect 35084 23492 35364 23548
rect 35084 23380 35140 23390
rect 34748 23044 34804 23054
rect 34804 22988 35028 23044
rect 34748 22950 34804 22988
rect 34636 22390 34692 22428
rect 34524 19954 34580 19964
rect 34636 21476 34692 21486
rect 34300 19294 34302 19346
rect 34354 19294 34356 19346
rect 34300 19282 34356 19294
rect 34636 19796 34692 21420
rect 34860 21028 34916 21038
rect 34972 21028 35028 22988
rect 35084 22372 35140 23324
rect 35308 23268 35364 23492
rect 36540 23378 36596 26852
rect 36764 25844 36820 25854
rect 36652 25508 36708 25518
rect 36652 24834 36708 25452
rect 36652 24782 36654 24834
rect 36706 24782 36708 24834
rect 36652 24770 36708 24782
rect 36540 23326 36542 23378
rect 36594 23326 36596 23378
rect 36540 23314 36596 23326
rect 35420 23268 35476 23278
rect 35308 23266 35476 23268
rect 35308 23214 35422 23266
rect 35474 23214 35476 23266
rect 35308 23212 35476 23214
rect 35420 23156 35476 23212
rect 35420 23090 35476 23100
rect 35980 23044 36036 23054
rect 35980 22950 36036 22988
rect 36204 22930 36260 22942
rect 36204 22878 36206 22930
rect 36258 22878 36260 22930
rect 35644 22820 35700 22830
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35532 22764 35644 22820
rect 35196 22372 35252 22382
rect 35084 22370 35252 22372
rect 35084 22318 35198 22370
rect 35250 22318 35252 22370
rect 35084 22316 35252 22318
rect 35196 22306 35252 22316
rect 35532 22258 35588 22764
rect 35644 22754 35700 22764
rect 36204 22372 36260 22878
rect 36764 22820 36820 25788
rect 36988 25618 37044 26852
rect 36988 25566 36990 25618
rect 37042 25566 37044 25618
rect 36988 25284 37044 25566
rect 37212 25508 37268 25518
rect 37212 25414 37268 25452
rect 36988 25218 37044 25228
rect 37100 24612 37156 24622
rect 36988 24556 37100 24612
rect 36876 23940 36932 23950
rect 36876 23266 36932 23884
rect 36988 23378 37044 24556
rect 37100 24518 37156 24556
rect 37324 24052 37380 26852
rect 37548 25620 37604 27580
rect 37660 26962 37716 26974
rect 37660 26910 37662 26962
rect 37714 26910 37716 26962
rect 37660 26852 37716 26910
rect 37660 25844 37716 26796
rect 37660 25778 37716 25788
rect 37772 25732 37828 29372
rect 37884 29426 37940 29438
rect 37884 29374 37886 29426
rect 37938 29374 37940 29426
rect 37884 25956 37940 29374
rect 37996 29428 38052 31054
rect 38108 31780 38164 33964
rect 38444 33954 38500 33964
rect 38556 32564 38612 35644
rect 38780 35588 38836 36204
rect 39340 35924 39396 41356
rect 39452 40516 39508 40526
rect 39452 40422 39508 40460
rect 38556 32498 38612 32508
rect 38668 35532 38836 35588
rect 39116 35868 39396 35924
rect 39452 39394 39508 39406
rect 39452 39342 39454 39394
rect 39506 39342 39508 39394
rect 38668 35476 38724 35532
rect 38444 32452 38500 32462
rect 38444 31890 38500 32396
rect 38444 31838 38446 31890
rect 38498 31838 38500 31890
rect 38444 31826 38500 31838
rect 38108 30324 38164 31724
rect 38220 31554 38276 31566
rect 38220 31502 38222 31554
rect 38274 31502 38276 31554
rect 38220 31444 38276 31502
rect 38332 31556 38388 31566
rect 38556 31556 38612 31566
rect 38332 31462 38388 31500
rect 38444 31554 38612 31556
rect 38444 31502 38558 31554
rect 38610 31502 38612 31554
rect 38444 31500 38612 31502
rect 38220 31378 38276 31388
rect 38444 31332 38500 31500
rect 38556 31490 38612 31500
rect 38444 31266 38500 31276
rect 38668 31108 38724 35420
rect 38892 35140 38948 35150
rect 38892 34020 38948 35084
rect 38892 34018 39060 34020
rect 38892 33966 38894 34018
rect 38946 33966 39060 34018
rect 38892 33964 39060 33966
rect 38892 33954 38948 33964
rect 38892 32564 38948 32574
rect 38892 32470 38948 32508
rect 38668 31042 38724 31052
rect 38780 31666 38836 31678
rect 38780 31614 38782 31666
rect 38834 31614 38836 31666
rect 38108 30258 38164 30268
rect 38220 30212 38276 30222
rect 38780 30212 38836 31614
rect 38892 31668 38948 31678
rect 39004 31668 39060 33964
rect 38948 31612 39060 31668
rect 39116 31890 39172 35868
rect 39340 35698 39396 35710
rect 39340 35646 39342 35698
rect 39394 35646 39396 35698
rect 39340 35028 39396 35646
rect 39452 35588 39508 39342
rect 39564 37380 39620 41580
rect 39900 40628 39956 40638
rect 40012 40628 40068 42590
rect 40348 42532 40404 42542
rect 40348 41970 40404 42476
rect 40348 41918 40350 41970
rect 40402 41918 40404 41970
rect 40348 41906 40404 41918
rect 40236 41860 40292 41870
rect 40236 41766 40292 41804
rect 40460 41188 40516 43596
rect 40796 42308 40852 44268
rect 41020 44258 41076 44268
rect 41356 44258 41412 44268
rect 40908 44100 40964 44110
rect 40908 44098 41188 44100
rect 40908 44046 40910 44098
rect 40962 44046 41188 44098
rect 40908 44044 41188 44046
rect 40908 44034 40964 44044
rect 41020 43876 41076 43886
rect 41020 43538 41076 43820
rect 41020 43486 41022 43538
rect 41074 43486 41076 43538
rect 41020 43474 41076 43486
rect 40796 42242 40852 42252
rect 41132 41636 41188 44044
rect 41244 44098 41300 44110
rect 41244 44046 41246 44098
rect 41298 44046 41300 44098
rect 41244 42196 41300 44046
rect 41468 43876 41524 45164
rect 41692 45218 41748 45836
rect 41804 45892 41860 45902
rect 41804 45330 41860 45836
rect 41804 45278 41806 45330
rect 41858 45278 41860 45330
rect 41804 45266 41860 45278
rect 41692 45166 41694 45218
rect 41746 45166 41748 45218
rect 41692 45154 41748 45166
rect 41468 43810 41524 43820
rect 41804 44882 41860 44894
rect 41804 44830 41806 44882
rect 41858 44830 41860 44882
rect 41692 43428 41748 43438
rect 41692 43334 41748 43372
rect 41804 42756 41860 44830
rect 42252 44436 42308 47628
rect 42364 47590 42420 47628
rect 44492 47572 44548 47582
rect 44828 47572 44884 48188
rect 48188 48020 48244 48860
rect 45388 47684 45444 47694
rect 45388 47590 45444 47628
rect 47516 47684 47572 47694
rect 47572 47628 47684 47684
rect 47516 47618 47572 47628
rect 44492 47570 44660 47572
rect 44492 47518 44494 47570
rect 44546 47518 44660 47570
rect 44492 47516 44660 47518
rect 44492 47506 44548 47516
rect 42812 47460 42868 47470
rect 43708 47460 43764 47470
rect 44156 47460 44212 47470
rect 42812 47458 43092 47460
rect 42812 47406 42814 47458
rect 42866 47406 43092 47458
rect 42812 47404 43092 47406
rect 42812 47394 42868 47404
rect 42924 47234 42980 47246
rect 42924 47182 42926 47234
rect 42978 47182 42980 47234
rect 42588 45892 42644 45902
rect 42588 45778 42644 45836
rect 42588 45726 42590 45778
rect 42642 45726 42644 45778
rect 42588 45714 42644 45726
rect 42700 45890 42756 45902
rect 42700 45838 42702 45890
rect 42754 45838 42756 45890
rect 42028 44380 42308 44436
rect 42364 45218 42420 45230
rect 42364 45166 42366 45218
rect 42418 45166 42420 45218
rect 42364 44436 42420 45166
rect 42476 44994 42532 45006
rect 42476 44942 42478 44994
rect 42530 44942 42532 44994
rect 42476 44548 42532 44942
rect 42700 44996 42756 45838
rect 42700 44930 42756 44940
rect 42588 44884 42644 44894
rect 42588 44790 42644 44828
rect 42476 44482 42532 44492
rect 42028 43092 42084 44380
rect 42364 44370 42420 44380
rect 42476 44324 42532 44334
rect 42700 44324 42756 44334
rect 42476 44322 42756 44324
rect 42476 44270 42478 44322
rect 42530 44270 42702 44322
rect 42754 44270 42756 44322
rect 42476 44268 42756 44270
rect 42476 44258 42532 44268
rect 42700 44258 42756 44268
rect 42924 44324 42980 47182
rect 43036 46004 43092 47404
rect 43708 47458 43876 47460
rect 43708 47406 43710 47458
rect 43762 47406 43876 47458
rect 43708 47404 43876 47406
rect 43708 47394 43764 47404
rect 43036 45890 43092 45948
rect 43036 45838 43038 45890
rect 43090 45838 43092 45890
rect 43036 45826 43092 45838
rect 43820 46562 43876 47404
rect 43820 46510 43822 46562
rect 43874 46510 43876 46562
rect 43260 45668 43316 45678
rect 43484 45668 43540 45678
rect 43260 45666 43428 45668
rect 43260 45614 43262 45666
rect 43314 45614 43428 45666
rect 43260 45612 43428 45614
rect 43260 45602 43316 45612
rect 42924 44258 42980 44268
rect 43036 45556 43092 45566
rect 43036 44322 43092 45500
rect 43036 44270 43038 44322
rect 43090 44270 43092 44322
rect 43036 44258 43092 44270
rect 43260 44996 43316 45006
rect 43260 44322 43316 44940
rect 43260 44270 43262 44322
rect 43314 44270 43316 44322
rect 43260 44258 43316 44270
rect 42140 44210 42196 44222
rect 42140 44158 42142 44210
rect 42194 44158 42196 44210
rect 42140 43316 42196 44158
rect 42252 44100 42308 44110
rect 42252 44098 42868 44100
rect 42252 44046 42254 44098
rect 42306 44046 42868 44098
rect 42252 44044 42868 44046
rect 42252 44034 42308 44044
rect 42140 43250 42196 43260
rect 42588 43428 42644 43438
rect 42028 43036 42308 43092
rect 41804 42690 41860 42700
rect 42140 42866 42196 42878
rect 42140 42814 42142 42866
rect 42194 42814 42196 42866
rect 41244 42130 41300 42140
rect 42140 42084 42196 42814
rect 41132 41570 41188 41580
rect 41356 42028 42196 42084
rect 39900 40626 40068 40628
rect 39900 40574 39902 40626
rect 39954 40574 40068 40626
rect 39900 40572 40068 40574
rect 40348 40628 40404 40638
rect 40460 40628 40516 41132
rect 41244 41188 41300 41198
rect 41244 40852 41300 41132
rect 41356 40964 41412 42028
rect 41692 41970 41748 42028
rect 42252 41972 42308 43036
rect 42588 42866 42644 43372
rect 42588 42814 42590 42866
rect 42642 42814 42644 42866
rect 42588 42802 42644 42814
rect 42476 42756 42532 42766
rect 42476 42662 42532 42700
rect 42812 42756 42868 44044
rect 43148 44098 43204 44110
rect 43148 44046 43150 44098
rect 43202 44046 43204 44098
rect 42812 42662 42868 42700
rect 42924 42754 42980 42766
rect 42924 42702 42926 42754
rect 42978 42702 42980 42754
rect 42700 42644 42756 42654
rect 42700 42082 42756 42588
rect 42700 42030 42702 42082
rect 42754 42030 42756 42082
rect 42700 42018 42756 42030
rect 41692 41918 41694 41970
rect 41746 41918 41748 41970
rect 41692 41906 41748 41918
rect 42140 41916 42308 41972
rect 41468 41860 41524 41870
rect 41804 41860 41860 41870
rect 41468 41858 41636 41860
rect 41468 41806 41470 41858
rect 41522 41806 41636 41858
rect 41468 41804 41636 41806
rect 41468 41794 41524 41804
rect 41580 41524 41636 41804
rect 41804 41766 41860 41804
rect 41580 41468 41972 41524
rect 41356 40908 41748 40964
rect 41244 40796 41636 40852
rect 40348 40626 40516 40628
rect 40348 40574 40350 40626
rect 40402 40574 40516 40626
rect 40348 40572 40516 40574
rect 41020 40628 41076 40638
rect 39900 40562 39956 40572
rect 40348 40562 40404 40572
rect 41020 40534 41076 40572
rect 39676 40404 39732 40414
rect 39676 39620 39732 40348
rect 39788 40290 39844 40302
rect 39788 40238 39790 40290
rect 39842 40238 39844 40290
rect 39788 39844 39844 40238
rect 41468 40292 41524 40302
rect 41468 40198 41524 40236
rect 41580 40068 41636 40796
rect 41468 40012 41636 40068
rect 39788 39778 39844 39788
rect 41244 39844 41300 39854
rect 39788 39620 39844 39630
rect 39676 39618 39844 39620
rect 39676 39566 39790 39618
rect 39842 39566 39844 39618
rect 39676 39564 39844 39566
rect 39788 39554 39844 39564
rect 40572 39508 40628 39518
rect 40348 39506 40628 39508
rect 40348 39454 40574 39506
rect 40626 39454 40628 39506
rect 40348 39452 40628 39454
rect 40348 39058 40404 39452
rect 40572 39442 40628 39452
rect 41020 39284 41076 39294
rect 40348 39006 40350 39058
rect 40402 39006 40404 39058
rect 40348 38994 40404 39006
rect 40684 39172 40740 39182
rect 40012 38948 40068 38958
rect 39900 38722 39956 38734
rect 39900 38670 39902 38722
rect 39954 38670 39956 38722
rect 39788 38610 39844 38622
rect 39788 38558 39790 38610
rect 39842 38558 39844 38610
rect 39676 38164 39732 38174
rect 39788 38164 39844 38558
rect 39676 38162 39844 38164
rect 39676 38110 39678 38162
rect 39730 38110 39844 38162
rect 39676 38108 39844 38110
rect 39676 38098 39732 38108
rect 39900 37716 39956 38670
rect 39900 37650 39956 37660
rect 39676 37492 39732 37502
rect 40012 37492 40068 38892
rect 40236 38724 40292 38762
rect 40236 38658 40292 38668
rect 40348 38500 40404 38510
rect 39676 37398 39732 37436
rect 39788 37436 40068 37492
rect 40236 38052 40292 38062
rect 39564 37314 39620 37324
rect 39788 37266 39844 37436
rect 40236 37378 40292 37996
rect 40348 38050 40404 38444
rect 40348 37998 40350 38050
rect 40402 37998 40404 38050
rect 40348 37986 40404 37998
rect 40236 37326 40238 37378
rect 40290 37326 40292 37378
rect 40236 37314 40292 37326
rect 39788 37214 39790 37266
rect 39842 37214 39844 37266
rect 39676 35812 39732 35822
rect 39452 35494 39508 35532
rect 39564 35756 39676 35812
rect 39340 34244 39396 34972
rect 39452 35028 39508 35038
rect 39564 35028 39620 35756
rect 39676 35746 39732 35756
rect 39452 35026 39620 35028
rect 39452 34974 39454 35026
rect 39506 34974 39620 35026
rect 39452 34972 39620 34974
rect 39676 35252 39732 35262
rect 39452 34962 39508 34972
rect 39564 34244 39620 34254
rect 39340 34242 39620 34244
rect 39340 34190 39566 34242
rect 39618 34190 39620 34242
rect 39340 34188 39620 34190
rect 39228 34130 39284 34142
rect 39228 34078 39230 34130
rect 39282 34078 39284 34130
rect 39228 33012 39284 34078
rect 39564 33908 39620 34188
rect 39564 33842 39620 33852
rect 39228 32946 39284 32956
rect 39116 31838 39118 31890
rect 39170 31838 39172 31890
rect 38892 31602 38948 31612
rect 39116 31444 39172 31838
rect 39676 31780 39732 35196
rect 39788 34804 39844 37214
rect 40012 37268 40068 37278
rect 40012 37174 40068 37212
rect 39900 37156 39956 37166
rect 39900 37062 39956 37100
rect 40012 36594 40068 36606
rect 40012 36542 40014 36594
rect 40066 36542 40068 36594
rect 39900 36482 39956 36494
rect 39900 36430 39902 36482
rect 39954 36430 39956 36482
rect 39900 35140 39956 36430
rect 39900 35074 39956 35084
rect 39788 34738 39844 34748
rect 40012 34356 40068 36542
rect 40348 36372 40404 36382
rect 40348 36370 40628 36372
rect 40348 36318 40350 36370
rect 40402 36318 40628 36370
rect 40348 36316 40628 36318
rect 40348 36306 40404 36316
rect 40124 36036 40180 36046
rect 40124 35922 40180 35980
rect 40124 35870 40126 35922
rect 40178 35870 40180 35922
rect 40124 35476 40180 35870
rect 40236 35924 40292 35934
rect 40572 35924 40628 36316
rect 40684 36370 40740 39116
rect 41020 39058 41076 39228
rect 41020 39006 41022 39058
rect 41074 39006 41076 39058
rect 41020 38994 41076 39006
rect 41132 39172 41188 39182
rect 41132 39058 41188 39116
rect 41132 39006 41134 39058
rect 41186 39006 41188 39058
rect 41132 38994 41188 39006
rect 41244 39058 41300 39788
rect 41244 39006 41246 39058
rect 41298 39006 41300 39058
rect 41244 38994 41300 39006
rect 41356 39732 41412 39742
rect 41356 39058 41412 39676
rect 41356 39006 41358 39058
rect 41410 39006 41412 39058
rect 41356 38994 41412 39006
rect 40908 38050 40964 38062
rect 40908 37998 40910 38050
rect 40962 37998 40964 38050
rect 40908 37380 40964 37998
rect 41020 37940 41076 37950
rect 41020 37490 41076 37884
rect 41020 37438 41022 37490
rect 41074 37438 41076 37490
rect 41020 37426 41076 37438
rect 41244 37828 41300 37838
rect 40908 37314 40964 37324
rect 40908 37156 40964 37166
rect 40908 37062 40964 37100
rect 40908 36596 40964 36606
rect 40908 36482 40964 36540
rect 40908 36430 40910 36482
rect 40962 36430 40964 36482
rect 40908 36418 40964 36430
rect 40684 36318 40686 36370
rect 40738 36318 40740 36370
rect 40684 36306 40740 36318
rect 40572 35868 40964 35924
rect 40236 35830 40292 35868
rect 40908 35810 40964 35868
rect 40908 35758 40910 35810
rect 40962 35758 40964 35810
rect 40908 35746 40964 35758
rect 41244 35700 41300 37772
rect 41468 37154 41524 40012
rect 41580 38948 41636 38958
rect 41692 38948 41748 40908
rect 41804 40516 41860 40526
rect 41804 40422 41860 40460
rect 41916 40404 41972 41468
rect 42140 41412 42196 41916
rect 42252 41746 42308 41758
rect 42252 41694 42254 41746
rect 42306 41694 42308 41746
rect 42252 41636 42308 41694
rect 42364 41748 42420 41758
rect 42588 41748 42644 41758
rect 42364 41654 42420 41692
rect 42476 41746 42644 41748
rect 42476 41694 42590 41746
rect 42642 41694 42644 41746
rect 42476 41692 42644 41694
rect 42252 41570 42308 41580
rect 42140 41356 42308 41412
rect 42140 41188 42196 41198
rect 42140 41094 42196 41132
rect 42252 40404 42308 41356
rect 42364 40964 42420 40974
rect 42364 40626 42420 40908
rect 42364 40574 42366 40626
rect 42418 40574 42420 40626
rect 42364 40562 42420 40574
rect 41916 40348 42084 40404
rect 42252 40348 42420 40404
rect 41916 40180 41972 40190
rect 41916 40086 41972 40124
rect 42028 39956 42084 40348
rect 41916 39900 42084 39956
rect 42252 40178 42308 40190
rect 42252 40126 42254 40178
rect 42306 40126 42308 40178
rect 41580 38946 41748 38948
rect 41580 38894 41582 38946
rect 41634 38894 41748 38946
rect 41580 38892 41748 38894
rect 41804 39172 41860 39182
rect 41580 38882 41636 38892
rect 41580 37940 41636 37950
rect 41580 37846 41636 37884
rect 41468 37102 41470 37154
rect 41522 37102 41524 37154
rect 41356 36258 41412 36270
rect 41356 36206 41358 36258
rect 41410 36206 41412 36258
rect 41356 35812 41412 36206
rect 41356 35746 41412 35756
rect 41132 35698 41300 35700
rect 41132 35646 41246 35698
rect 41298 35646 41300 35698
rect 41132 35644 41300 35646
rect 40348 35476 40404 35486
rect 40124 35420 40292 35476
rect 40236 35252 40292 35420
rect 40348 35382 40404 35420
rect 40236 35186 40292 35196
rect 40236 34916 40292 34926
rect 40236 34822 40292 34860
rect 41020 34916 41076 34926
rect 40684 34412 40964 34468
rect 40236 34356 40292 34366
rect 40012 34354 40292 34356
rect 40012 34302 40238 34354
rect 40290 34302 40292 34354
rect 40012 34300 40292 34302
rect 39900 34242 39956 34254
rect 39900 34190 39902 34242
rect 39954 34190 39956 34242
rect 39900 33460 39956 34190
rect 39900 33394 39956 33404
rect 40012 33124 40068 33134
rect 40012 33122 40180 33124
rect 40012 33070 40014 33122
rect 40066 33070 40180 33122
rect 40012 33068 40180 33070
rect 40012 33058 40068 33068
rect 40012 31780 40068 31790
rect 39676 31778 40068 31780
rect 39676 31726 40014 31778
rect 40066 31726 40068 31778
rect 39676 31724 40068 31726
rect 39116 31378 39172 31388
rect 39340 31668 39396 31678
rect 37996 27748 38052 29372
rect 37996 27682 38052 27692
rect 38108 29988 38164 29998
rect 38108 28196 38164 29932
rect 38108 27188 38164 28140
rect 38220 27858 38276 30156
rect 38444 30156 38836 30212
rect 38892 31332 38948 31342
rect 38332 29426 38388 29438
rect 38332 29374 38334 29426
rect 38386 29374 38388 29426
rect 38332 28532 38388 29374
rect 38444 29314 38500 30156
rect 38444 29262 38446 29314
rect 38498 29262 38500 29314
rect 38444 28756 38500 29262
rect 38444 28690 38500 28700
rect 38556 29202 38612 29214
rect 38556 29150 38558 29202
rect 38610 29150 38612 29202
rect 38332 28466 38388 28476
rect 38556 28420 38612 29150
rect 38668 29204 38724 29214
rect 38668 28642 38724 29148
rect 38668 28590 38670 28642
rect 38722 28590 38724 28642
rect 38668 28578 38724 28590
rect 38556 28364 38836 28420
rect 38220 27806 38222 27858
rect 38274 27806 38276 27858
rect 38220 27794 38276 27806
rect 38444 27858 38500 27870
rect 38444 27806 38446 27858
rect 38498 27806 38500 27858
rect 38332 27188 38388 27198
rect 38108 27186 38388 27188
rect 38108 27134 38334 27186
rect 38386 27134 38388 27186
rect 38108 27132 38388 27134
rect 38332 27122 38388 27132
rect 37996 26964 38052 26974
rect 37996 26870 38052 26908
rect 38444 26908 38500 27806
rect 38780 27858 38836 28364
rect 38780 27806 38782 27858
rect 38834 27806 38836 27858
rect 38780 27794 38836 27806
rect 38668 27748 38724 27758
rect 38444 26852 38612 26908
rect 38444 26180 38500 26190
rect 37884 25890 37940 25900
rect 37996 26178 38500 26180
rect 37996 26126 38446 26178
rect 38498 26126 38500 26178
rect 37996 26124 38500 26126
rect 37772 25676 37940 25732
rect 37548 25564 37716 25620
rect 37324 23938 37380 23996
rect 37324 23886 37326 23938
rect 37378 23886 37380 23938
rect 37324 23874 37380 23886
rect 37436 25508 37492 25518
rect 36988 23326 36990 23378
rect 37042 23326 37044 23378
rect 36988 23314 37044 23326
rect 37212 23380 37268 23390
rect 37436 23380 37492 25452
rect 37548 25282 37604 25294
rect 37548 25230 37550 25282
rect 37602 25230 37604 25282
rect 37548 24050 37604 25230
rect 37548 23998 37550 24050
rect 37602 23998 37604 24050
rect 37548 23940 37604 23998
rect 37548 23874 37604 23884
rect 37212 23378 37492 23380
rect 37212 23326 37214 23378
rect 37266 23326 37492 23378
rect 37212 23324 37492 23326
rect 37212 23314 37268 23324
rect 36876 23214 36878 23266
rect 36930 23214 36932 23266
rect 36876 23202 36932 23214
rect 37548 23266 37604 23278
rect 37548 23214 37550 23266
rect 37602 23214 37604 23266
rect 37324 22932 37380 22942
rect 36876 22820 36932 22830
rect 36764 22764 36876 22820
rect 36876 22754 36932 22764
rect 36764 22484 36820 22494
rect 36820 22428 36932 22484
rect 36764 22418 36820 22428
rect 36204 22306 36260 22316
rect 35532 22206 35534 22258
rect 35586 22206 35588 22258
rect 35532 22194 35588 22206
rect 36092 22146 36148 22158
rect 36428 22148 36484 22158
rect 36092 22094 36094 22146
rect 36146 22094 36148 22146
rect 35980 21812 36036 21822
rect 35980 21718 36036 21756
rect 35084 21588 35140 21598
rect 35084 21494 35140 21532
rect 35532 21586 35588 21598
rect 35532 21534 35534 21586
rect 35586 21534 35588 21586
rect 35532 21476 35588 21534
rect 35756 21476 35812 21486
rect 35532 21420 35756 21476
rect 35756 21410 35812 21420
rect 36092 21476 36148 22094
rect 36204 22092 36428 22148
rect 36204 21698 36260 22092
rect 36428 22054 36484 22092
rect 36652 21812 36708 21822
rect 36204 21646 36206 21698
rect 36258 21646 36260 21698
rect 36204 21634 36260 21646
rect 36316 21810 36708 21812
rect 36316 21758 36654 21810
rect 36706 21758 36708 21810
rect 36316 21756 36708 21758
rect 36092 21410 36148 21420
rect 35420 21364 35476 21374
rect 35868 21364 35924 21374
rect 35420 21362 35588 21364
rect 35420 21310 35422 21362
rect 35474 21310 35588 21362
rect 35420 21308 35588 21310
rect 35420 21298 35476 21308
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 21028 35140 21038
rect 34860 21026 35140 21028
rect 34860 20974 34862 21026
rect 34914 20974 35086 21026
rect 35138 20974 35140 21026
rect 34860 20972 35140 20974
rect 34860 20962 34916 20972
rect 35084 20962 35140 20972
rect 35420 21028 35476 21038
rect 35532 21028 35588 21308
rect 35868 21270 35924 21308
rect 35420 21026 35532 21028
rect 35420 20974 35422 21026
rect 35474 20974 35532 21026
rect 35420 20972 35532 20974
rect 35420 20962 35476 20972
rect 35532 20934 35588 20972
rect 35980 21028 36036 21038
rect 35196 20804 35252 20814
rect 35196 20690 35252 20748
rect 35980 20802 36036 20972
rect 35980 20750 35982 20802
rect 36034 20750 36036 20802
rect 35980 20738 36036 20750
rect 36316 20802 36372 21756
rect 36652 21746 36708 21756
rect 36540 21586 36596 21598
rect 36540 21534 36542 21586
rect 36594 21534 36596 21586
rect 36316 20750 36318 20802
rect 36370 20750 36372 20802
rect 36316 20738 36372 20750
rect 36428 21476 36484 21486
rect 35196 20638 35198 20690
rect 35250 20638 35252 20690
rect 35196 20626 35252 20638
rect 35756 20690 35812 20702
rect 35756 20638 35758 20690
rect 35810 20638 35812 20690
rect 34748 20580 34804 20590
rect 34748 20468 34804 20524
rect 35756 20580 35812 20638
rect 35756 20514 35812 20524
rect 35868 20578 35924 20590
rect 35868 20526 35870 20578
rect 35922 20526 35924 20578
rect 34748 20412 35140 20468
rect 35084 20018 35140 20412
rect 35868 20244 35924 20526
rect 35868 20178 35924 20188
rect 35084 19966 35086 20018
rect 35138 19966 35140 20018
rect 35084 19954 35140 19966
rect 34636 19236 34692 19740
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 36428 19346 36484 21420
rect 36428 19294 36430 19346
rect 36482 19294 36484 19346
rect 36428 19282 36484 19294
rect 34636 19170 34692 19180
rect 35420 19236 35476 19246
rect 34412 19012 34468 19022
rect 34076 18956 34244 19012
rect 32900 17724 33012 17780
rect 32844 17686 32900 17724
rect 32508 17668 32564 17678
rect 31724 17108 31780 17118
rect 30940 17106 31780 17108
rect 30940 17054 31726 17106
rect 31778 17054 31780 17106
rect 30940 17052 31780 17054
rect 30268 16902 30324 16940
rect 30604 16996 30660 17006
rect 30156 16772 30212 16782
rect 30156 16678 30212 16716
rect 30156 16436 30212 16446
rect 30156 16210 30212 16380
rect 30156 16158 30158 16210
rect 30210 16158 30212 16210
rect 30156 16146 30212 16158
rect 30604 16210 30660 16940
rect 30940 16994 30996 17052
rect 31724 17042 31780 17052
rect 31836 17108 31892 17118
rect 32284 17108 32340 17500
rect 31836 17106 32340 17108
rect 31836 17054 31838 17106
rect 31890 17054 32340 17106
rect 31836 17052 32340 17054
rect 32396 17612 32508 17668
rect 31836 17042 31892 17052
rect 32396 16996 32452 17612
rect 32508 17602 32564 17612
rect 30940 16942 30942 16994
rect 30994 16942 30996 16994
rect 30940 16930 30996 16942
rect 32284 16940 32452 16996
rect 31276 16884 31332 16894
rect 30604 16158 30606 16210
rect 30658 16158 30660 16210
rect 30604 16146 30660 16158
rect 30828 16658 30884 16670
rect 30828 16606 30830 16658
rect 30882 16606 30884 16658
rect 30828 15540 30884 16606
rect 31276 16660 31332 16828
rect 31500 16884 31556 16894
rect 31500 16790 31556 16828
rect 31612 16882 31668 16894
rect 31612 16830 31614 16882
rect 31666 16830 31668 16882
rect 31612 16660 31668 16830
rect 32060 16882 32116 16894
rect 32060 16830 32062 16882
rect 32114 16830 32116 16882
rect 31276 16604 31668 16660
rect 31724 16772 31780 16782
rect 30828 15474 30884 15484
rect 30604 15428 30660 15438
rect 30604 15334 30660 15372
rect 30828 15316 30884 15326
rect 30828 15222 30884 15260
rect 30716 15204 30772 15214
rect 30044 15092 30212 15148
rect 30044 14644 30100 14654
rect 29932 14642 30100 14644
rect 29932 14590 30046 14642
rect 30098 14590 30100 14642
rect 29932 14588 30100 14590
rect 30044 14578 30100 14588
rect 30156 14532 30212 15092
rect 30156 14466 30212 14476
rect 29932 13636 29988 13646
rect 29932 13542 29988 13580
rect 30268 13074 30324 13086
rect 30268 13022 30270 13074
rect 30322 13022 30324 13074
rect 29708 12964 29764 12974
rect 29932 12964 29988 12974
rect 29708 12962 29876 12964
rect 29708 12910 29710 12962
rect 29762 12910 29876 12962
rect 29708 12908 29876 12910
rect 29708 12898 29764 12908
rect 29708 12180 29764 12190
rect 29708 12086 29764 12124
rect 29596 11342 29598 11394
rect 29650 11342 29652 11394
rect 29372 10518 29428 10556
rect 29148 10098 29204 10108
rect 28476 9762 28532 9772
rect 29372 9826 29428 9838
rect 29372 9774 29374 9826
rect 29426 9774 29428 9826
rect 28588 9716 28644 9726
rect 29372 9716 29428 9774
rect 28588 9714 28980 9716
rect 28588 9662 28590 9714
rect 28642 9662 28980 9714
rect 28588 9660 28980 9662
rect 28588 9650 28644 9660
rect 28364 9214 28366 9266
rect 28418 9214 28420 9266
rect 28364 9202 28420 9214
rect 28924 9044 28980 9660
rect 29372 9650 29428 9660
rect 29596 9714 29652 11342
rect 29820 11284 29876 12908
rect 29932 12870 29988 12908
rect 30268 12516 30324 13022
rect 30380 13076 30436 13086
rect 30380 12962 30436 13020
rect 30380 12910 30382 12962
rect 30434 12910 30436 12962
rect 30380 12898 30436 12910
rect 30716 12850 30772 15148
rect 31724 14084 31780 16716
rect 32060 15428 32116 16830
rect 32284 16436 32340 16940
rect 32284 16370 32340 16380
rect 32396 16770 32452 16782
rect 32396 16718 32398 16770
rect 32450 16718 32452 16770
rect 32396 15988 32452 16718
rect 32508 16660 32564 16670
rect 32956 16660 33012 17724
rect 33068 17714 33124 17724
rect 33180 17892 33236 17902
rect 33852 17892 33908 18956
rect 33964 18452 34020 18462
rect 33964 18358 34020 18396
rect 33180 17890 33908 17892
rect 33180 17838 33182 17890
rect 33234 17838 33908 17890
rect 33180 17836 33908 17838
rect 33180 16884 33236 17836
rect 33516 17668 33572 17678
rect 33516 17574 33572 17612
rect 33852 17666 33908 17836
rect 34076 17892 34132 17902
rect 33964 17780 34020 17790
rect 33964 17686 34020 17724
rect 33852 17614 33854 17666
rect 33906 17614 33908 17666
rect 33852 17602 33908 17614
rect 34076 17666 34132 17836
rect 34076 17614 34078 17666
rect 34130 17614 34132 17666
rect 34076 17602 34132 17614
rect 33292 17556 33348 17566
rect 33292 17462 33348 17500
rect 33516 17444 33572 17454
rect 33404 17220 33460 17230
rect 33404 17106 33460 17164
rect 33404 17054 33406 17106
rect 33458 17054 33460 17106
rect 33404 17042 33460 17054
rect 33516 16994 33572 17388
rect 34076 17444 34132 17454
rect 33516 16942 33518 16994
rect 33570 16942 33572 16994
rect 33516 16930 33572 16942
rect 33964 16996 34020 17006
rect 33964 16902 34020 16940
rect 34076 16994 34132 17388
rect 34076 16942 34078 16994
rect 34130 16942 34132 16994
rect 34076 16930 34132 16942
rect 34188 16996 34244 18956
rect 34300 17556 34356 17566
rect 34300 17462 34356 17500
rect 34412 17444 34468 18956
rect 35420 18452 35476 19180
rect 35868 18900 35924 18910
rect 35420 18396 35700 18452
rect 34524 18340 34580 18350
rect 34524 17668 34580 18284
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 34524 17666 35028 17668
rect 34524 17614 34526 17666
rect 34578 17614 35028 17666
rect 34524 17612 35028 17614
rect 34524 17602 34580 17612
rect 34468 17388 34692 17444
rect 34412 17350 34468 17388
rect 34524 16996 34580 17006
rect 34188 16994 34580 16996
rect 34188 16942 34526 16994
rect 34578 16942 34580 16994
rect 34188 16940 34580 16942
rect 33180 16818 33236 16828
rect 34524 16884 34580 16940
rect 34636 16994 34692 17388
rect 34636 16942 34638 16994
rect 34690 16942 34692 16994
rect 34636 16930 34692 16942
rect 34972 16996 35028 17612
rect 35420 17556 35476 17566
rect 35420 17462 35476 17500
rect 35084 17444 35140 17454
rect 35084 17442 35252 17444
rect 35084 17390 35086 17442
rect 35138 17390 35252 17442
rect 35084 17388 35252 17390
rect 35084 17378 35140 17388
rect 35084 16996 35140 17006
rect 34972 16994 35140 16996
rect 34972 16942 35086 16994
rect 35138 16942 35140 16994
rect 34972 16940 35140 16942
rect 35084 16930 35140 16940
rect 34524 16818 34580 16828
rect 35196 16772 35252 17388
rect 35532 17332 35588 17342
rect 35532 17106 35588 17276
rect 35532 17054 35534 17106
rect 35586 17054 35588 17106
rect 35532 17042 35588 17054
rect 35196 16706 35252 16716
rect 33404 16660 33460 16670
rect 32508 16658 32900 16660
rect 32508 16606 32510 16658
rect 32562 16606 32900 16658
rect 32508 16604 32900 16606
rect 32956 16604 33348 16660
rect 32508 16594 32564 16604
rect 32396 15932 32564 15988
rect 31500 13748 31556 13758
rect 31388 13524 31444 13534
rect 30716 12798 30718 12850
rect 30770 12798 30772 12850
rect 30716 12786 30772 12798
rect 31052 12964 31108 12974
rect 30044 12460 30324 12516
rect 30044 11732 30100 12460
rect 30156 12292 30212 12302
rect 30156 12198 30212 12236
rect 31052 12292 31108 12908
rect 31388 12850 31444 13468
rect 31500 12962 31556 13692
rect 31500 12910 31502 12962
rect 31554 12910 31556 12962
rect 31500 12898 31556 12910
rect 31612 13076 31668 13086
rect 31388 12798 31390 12850
rect 31442 12798 31444 12850
rect 31388 12786 31444 12798
rect 31052 12198 31108 12236
rect 31164 12178 31220 12190
rect 31164 12126 31166 12178
rect 31218 12126 31220 12178
rect 30268 11956 30324 11966
rect 31164 11956 31220 12126
rect 31612 12178 31668 13020
rect 31612 12126 31614 12178
rect 31666 12126 31668 12178
rect 31612 12114 31668 12126
rect 30268 11954 31220 11956
rect 30268 11902 30270 11954
rect 30322 11902 31220 11954
rect 30268 11900 31220 11902
rect 30268 11890 30324 11900
rect 30044 11666 30100 11676
rect 30268 11732 30324 11742
rect 30268 11394 30324 11676
rect 30940 11508 30996 11518
rect 30940 11414 30996 11452
rect 30268 11342 30270 11394
rect 30322 11342 30324 11394
rect 30268 11330 30324 11342
rect 29820 11218 29876 11228
rect 30044 11172 30100 11182
rect 30044 10724 30100 11116
rect 30044 10610 30100 10668
rect 30044 10558 30046 10610
rect 30098 10558 30100 10610
rect 30044 10546 30100 10558
rect 31164 10610 31220 11900
rect 31164 10558 31166 10610
rect 31218 10558 31220 10610
rect 31164 10546 31220 10558
rect 31276 12066 31332 12078
rect 31276 12014 31278 12066
rect 31330 12014 31332 12066
rect 31276 11396 31332 12014
rect 31724 11788 31780 14028
rect 31836 15202 31892 15214
rect 31836 15150 31838 15202
rect 31890 15150 31892 15202
rect 31836 13860 31892 15150
rect 32060 15148 32116 15372
rect 32284 15540 32340 15550
rect 32284 15426 32340 15484
rect 32284 15374 32286 15426
rect 32338 15374 32340 15426
rect 32284 15362 32340 15374
rect 32396 15426 32452 15438
rect 32396 15374 32398 15426
rect 32450 15374 32452 15426
rect 31948 15092 32004 15102
rect 32060 15092 32228 15148
rect 31948 14998 32004 15036
rect 32172 14642 32228 15092
rect 32172 14590 32174 14642
rect 32226 14590 32228 14642
rect 32172 14578 32228 14590
rect 31836 13636 31892 13804
rect 32060 13636 32116 13646
rect 31836 13634 32116 13636
rect 31836 13582 32062 13634
rect 32114 13582 32116 13634
rect 31836 13580 32116 13582
rect 31836 13412 31892 13422
rect 31836 12402 31892 13356
rect 32060 12962 32116 13580
rect 32060 12910 32062 12962
rect 32114 12910 32116 12962
rect 32060 12898 32116 12910
rect 32396 12516 32452 15374
rect 32508 14980 32564 15932
rect 32508 14914 32564 14924
rect 32620 15314 32676 15326
rect 32620 15262 32622 15314
rect 32674 15262 32676 15314
rect 32620 13972 32676 15262
rect 32732 15316 32788 15326
rect 32732 14532 32788 15260
rect 32732 14438 32788 14476
rect 32508 13748 32564 13758
rect 32508 13654 32564 13692
rect 32620 13076 32676 13916
rect 32732 14196 32788 14206
rect 32732 13748 32788 14140
rect 32732 13682 32788 13692
rect 32844 13186 32900 16604
rect 32956 15428 33012 15438
rect 33180 15428 33236 15438
rect 33012 15426 33236 15428
rect 33012 15374 33182 15426
rect 33234 15374 33236 15426
rect 33012 15372 33236 15374
rect 32956 15362 33012 15372
rect 33180 15362 33236 15372
rect 33068 15204 33124 15242
rect 33068 15138 33124 15148
rect 33068 13748 33124 13758
rect 33068 13654 33124 13692
rect 33292 13746 33348 16604
rect 33404 16566 33460 16604
rect 33964 16658 34020 16670
rect 33964 16606 33966 16658
rect 34018 16606 34020 16658
rect 33516 15986 33572 15998
rect 33516 15934 33518 15986
rect 33570 15934 33572 15986
rect 33516 15316 33572 15934
rect 33516 15222 33572 15260
rect 33852 15540 33908 15550
rect 33852 15204 33908 15484
rect 33516 14980 33572 14990
rect 33516 14756 33572 14924
rect 33292 13694 33294 13746
rect 33346 13694 33348 13746
rect 33292 13682 33348 13694
rect 33404 14418 33460 14430
rect 33404 14366 33406 14418
rect 33458 14366 33460 14418
rect 32844 13134 32846 13186
rect 32898 13134 32900 13186
rect 32844 13122 32900 13134
rect 33292 13300 33348 13310
rect 32620 13020 32788 13076
rect 32732 12964 32788 13020
rect 33068 12964 33124 12974
rect 32732 12962 33124 12964
rect 32732 12910 33070 12962
rect 33122 12910 33124 12962
rect 32732 12908 33124 12910
rect 33068 12898 33124 12908
rect 33292 12964 33348 13244
rect 33404 13074 33460 14366
rect 33516 13970 33572 14700
rect 33516 13918 33518 13970
rect 33570 13918 33572 13970
rect 33516 13906 33572 13918
rect 33740 13860 33796 13870
rect 33740 13766 33796 13804
rect 33628 13634 33684 13646
rect 33852 13636 33908 15148
rect 33628 13582 33630 13634
rect 33682 13582 33684 13634
rect 33516 13524 33572 13534
rect 33628 13524 33684 13582
rect 33572 13468 33684 13524
rect 33740 13580 33908 13636
rect 33516 13458 33572 13468
rect 33740 13300 33796 13580
rect 33404 13022 33406 13074
rect 33458 13022 33460 13074
rect 33404 13010 33460 13022
rect 33516 13244 33796 13300
rect 33292 12870 33348 12908
rect 33516 12962 33572 13244
rect 33516 12910 33518 12962
rect 33570 12910 33572 12962
rect 33516 12898 33572 12910
rect 31836 12350 31838 12402
rect 31890 12350 31892 12402
rect 31836 12338 31892 12350
rect 32284 12460 32452 12516
rect 33404 12852 33460 12862
rect 31948 12180 32004 12190
rect 30716 10500 30772 10510
rect 29596 9662 29598 9714
rect 29650 9662 29652 9714
rect 29596 9650 29652 9662
rect 30604 10498 30772 10500
rect 30604 10446 30718 10498
rect 30770 10446 30772 10498
rect 30604 10444 30772 10446
rect 30268 9602 30324 9614
rect 30268 9550 30270 9602
rect 30322 9550 30324 9602
rect 27916 8878 27918 8930
rect 27970 8878 27972 8930
rect 27916 8866 27972 8878
rect 28700 8930 28756 8942
rect 28700 8878 28702 8930
rect 28754 8878 28756 8930
rect 26236 8372 26516 8428
rect 26796 8372 27076 8428
rect 28588 8820 28644 8830
rect 28140 8372 28196 8382
rect 26236 8370 26292 8372
rect 26236 8318 26238 8370
rect 26290 8318 26292 8370
rect 26236 8306 26292 8318
rect 26796 8258 26852 8372
rect 26796 8206 26798 8258
rect 26850 8206 26852 8258
rect 26796 8194 26852 8206
rect 26572 8148 26628 8158
rect 26572 8054 26628 8092
rect 27692 8146 27748 8158
rect 27692 8094 27694 8146
rect 27746 8094 27748 8146
rect 27580 8036 27636 8046
rect 27580 7942 27636 7980
rect 26124 7746 26180 7756
rect 25900 5854 25902 5906
rect 25954 5854 25956 5906
rect 25900 5842 25956 5854
rect 26012 7476 26068 7486
rect 25676 4386 25732 4396
rect 25788 4452 25844 4462
rect 26012 4452 26068 7420
rect 27132 7476 27188 7486
rect 27580 7476 27636 7486
rect 27692 7476 27748 8094
rect 28140 8146 28196 8316
rect 28364 8260 28420 8270
rect 28364 8166 28420 8204
rect 28588 8258 28644 8764
rect 28700 8372 28756 8878
rect 28700 8306 28756 8316
rect 28924 8428 28980 8988
rect 29372 9380 29428 9390
rect 29148 8820 29204 8830
rect 29148 8726 29204 8764
rect 28924 8372 29204 8428
rect 28588 8206 28590 8258
rect 28642 8206 28644 8258
rect 28588 8194 28644 8206
rect 28924 8260 28980 8372
rect 28924 8194 28980 8204
rect 29148 8258 29204 8372
rect 29148 8206 29150 8258
rect 29202 8206 29204 8258
rect 29148 8194 29204 8206
rect 28140 8094 28142 8146
rect 28194 8094 28196 8146
rect 28140 8082 28196 8094
rect 28476 8036 28532 8046
rect 28476 7942 28532 7980
rect 29260 8034 29316 8046
rect 29260 7982 29262 8034
rect 29314 7982 29316 8034
rect 26460 7364 26516 7374
rect 26460 7250 26516 7308
rect 26460 7198 26462 7250
rect 26514 7198 26516 7250
rect 26460 7186 26516 7198
rect 26908 6580 26964 6590
rect 26908 5906 26964 6524
rect 27132 6018 27188 7420
rect 27132 5966 27134 6018
rect 27186 5966 27188 6018
rect 27132 5954 27188 5966
rect 27244 7474 27748 7476
rect 27244 7422 27582 7474
rect 27634 7422 27748 7474
rect 27244 7420 27748 7422
rect 27804 7474 27860 7486
rect 27804 7422 27806 7474
rect 27858 7422 27860 7474
rect 26908 5854 26910 5906
rect 26962 5854 26964 5906
rect 26908 5842 26964 5854
rect 26572 5684 26628 5694
rect 26572 5590 26628 5628
rect 27020 5684 27076 5694
rect 26460 5124 26516 5134
rect 25788 4450 26068 4452
rect 25788 4398 25790 4450
rect 25842 4398 26068 4450
rect 25788 4396 26068 4398
rect 26348 4900 26404 4910
rect 25788 4386 25844 4396
rect 25452 4340 25508 4350
rect 23100 4274 23156 4284
rect 23772 4338 24500 4340
rect 23772 4286 24110 4338
rect 24162 4286 24500 4338
rect 23772 4284 24500 4286
rect 23324 4228 23380 4238
rect 23324 4134 23380 4172
rect 22988 3614 22990 3666
rect 23042 3614 23044 3666
rect 22988 3602 23044 3614
rect 23772 3554 23828 4284
rect 24108 4274 24164 4284
rect 23772 3502 23774 3554
rect 23826 3502 23828 3554
rect 23772 3490 23828 3502
rect 24444 3556 24500 4284
rect 25452 4246 25508 4284
rect 25340 4228 25396 4238
rect 25340 4134 25396 4172
rect 26236 4226 26292 4238
rect 26236 4174 26238 4226
rect 26290 4174 26292 4226
rect 24556 4116 24612 4126
rect 24556 4022 24612 4060
rect 26124 4116 26180 4126
rect 26124 4022 26180 4060
rect 26236 3780 26292 4174
rect 25340 3724 26292 3780
rect 25340 3666 25396 3724
rect 25340 3614 25342 3666
rect 25394 3614 25396 3666
rect 25340 3602 25396 3614
rect 24556 3556 24612 3566
rect 24444 3554 24612 3556
rect 24444 3502 24558 3554
rect 24610 3502 24612 3554
rect 24444 3500 24612 3502
rect 24556 3490 24612 3500
rect 24444 3332 24500 3342
rect 22540 2156 22708 2212
rect 22652 800 22708 2156
rect 24444 800 24500 3276
rect 26348 2436 26404 4844
rect 26460 4338 26516 5068
rect 26684 4452 26740 4462
rect 26684 4358 26740 4396
rect 26908 4450 26964 4462
rect 26908 4398 26910 4450
rect 26962 4398 26964 4450
rect 26460 4286 26462 4338
rect 26514 4286 26516 4338
rect 26460 4274 26516 4286
rect 26908 4228 26964 4398
rect 27020 4450 27076 5628
rect 27132 5236 27188 5246
rect 27244 5236 27300 7420
rect 27580 7410 27636 7420
rect 27804 6132 27860 7422
rect 28028 7474 28084 7486
rect 28028 7422 28030 7474
rect 28082 7422 28084 7474
rect 28028 6580 28084 7422
rect 28476 7476 28532 7486
rect 28476 7382 28532 7420
rect 29260 7476 29316 7982
rect 29260 7410 29316 7420
rect 28028 6514 28084 6524
rect 29036 6580 29092 6590
rect 29036 6486 29092 6524
rect 27692 6076 27860 6132
rect 28588 6468 28644 6478
rect 27468 5684 27524 5694
rect 27468 5346 27524 5628
rect 27468 5294 27470 5346
rect 27522 5294 27524 5346
rect 27468 5282 27524 5294
rect 27132 5234 27300 5236
rect 27132 5182 27134 5234
rect 27186 5182 27300 5234
rect 27132 5180 27300 5182
rect 27132 5170 27188 5180
rect 27580 5124 27636 5134
rect 27580 5030 27636 5068
rect 27692 5010 27748 6076
rect 28588 6018 28644 6412
rect 28588 5966 28590 6018
rect 28642 5966 28644 6018
rect 28588 5954 28644 5966
rect 27692 4958 27694 5010
rect 27746 4958 27748 5010
rect 27692 4676 27748 4958
rect 27020 4398 27022 4450
rect 27074 4398 27076 4450
rect 27020 4386 27076 4398
rect 27468 4620 27748 4676
rect 27804 5908 27860 5918
rect 27468 4228 27524 4620
rect 27580 4340 27636 4350
rect 27804 4340 27860 5852
rect 29260 5124 29316 5134
rect 29372 5124 29428 9324
rect 30156 9156 30212 9166
rect 30268 9156 30324 9550
rect 30156 9154 30324 9156
rect 30156 9102 30158 9154
rect 30210 9102 30324 9154
rect 30156 9100 30324 9102
rect 29820 9044 29876 9054
rect 29820 8950 29876 8988
rect 30044 9044 30100 9054
rect 30044 8950 30100 8988
rect 29596 8818 29652 8830
rect 29596 8766 29598 8818
rect 29650 8766 29652 8818
rect 29596 8428 29652 8766
rect 30156 8820 30212 9100
rect 29596 8372 30100 8428
rect 29484 6692 29540 6702
rect 29596 6692 29652 8372
rect 29484 6690 29652 6692
rect 29484 6638 29486 6690
rect 29538 6638 29652 6690
rect 29484 6636 29652 6638
rect 29708 8036 29764 8046
rect 29708 6690 29764 7980
rect 30044 7586 30100 8372
rect 30156 8146 30212 8764
rect 30156 8094 30158 8146
rect 30210 8094 30212 8146
rect 30156 8082 30212 8094
rect 30268 8036 30324 8046
rect 30268 7698 30324 7980
rect 30268 7646 30270 7698
rect 30322 7646 30324 7698
rect 30268 7634 30324 7646
rect 30492 7588 30548 7598
rect 30044 7534 30046 7586
rect 30098 7534 30100 7586
rect 30044 7522 30100 7534
rect 30380 7586 30548 7588
rect 30380 7534 30494 7586
rect 30546 7534 30548 7586
rect 30380 7532 30548 7534
rect 29708 6638 29710 6690
rect 29762 6638 29764 6690
rect 29484 6626 29540 6636
rect 29708 6626 29764 6638
rect 29932 7476 29988 7486
rect 30380 7476 30436 7532
rect 30492 7522 30548 7532
rect 29932 6578 29988 7420
rect 30156 7420 30436 7476
rect 30604 7476 30660 10444
rect 30716 10434 30772 10444
rect 30940 9828 30996 9838
rect 30940 9734 30996 9772
rect 31276 9826 31332 11340
rect 31612 11732 31780 11788
rect 31836 11844 31892 11854
rect 31388 11284 31444 11294
rect 31388 10612 31444 11228
rect 31612 10834 31668 11732
rect 31724 11620 31780 11630
rect 31836 11620 31892 11788
rect 31948 11732 32004 12124
rect 31948 11666 32004 11676
rect 31780 11564 31892 11620
rect 32284 11620 32340 12460
rect 32508 12348 33124 12404
rect 32396 12292 32452 12302
rect 32396 12198 32452 12236
rect 32508 12290 32564 12348
rect 32508 12238 32510 12290
rect 32562 12238 32564 12290
rect 32508 12226 32564 12238
rect 32844 12180 32900 12190
rect 31724 11554 31780 11564
rect 31836 11172 31892 11182
rect 31612 10782 31614 10834
rect 31666 10782 31668 10834
rect 31612 10770 31668 10782
rect 31724 10836 31780 10846
rect 31724 10742 31780 10780
rect 31836 10834 31892 11116
rect 31836 10782 31838 10834
rect 31890 10782 31892 10834
rect 31836 10770 31892 10782
rect 32284 10836 32340 11564
rect 32508 11732 32564 11742
rect 32508 11172 32564 11676
rect 32396 10836 32452 10846
rect 32284 10834 32452 10836
rect 32284 10782 32398 10834
rect 32450 10782 32452 10834
rect 32284 10780 32452 10782
rect 32396 10770 32452 10780
rect 32508 10722 32564 11116
rect 32508 10670 32510 10722
rect 32562 10670 32564 10722
rect 32508 10658 32564 10670
rect 31388 10518 31444 10556
rect 32172 10612 32228 10622
rect 32172 10518 32228 10556
rect 31276 9774 31278 9826
rect 31330 9774 31332 9826
rect 31276 9762 31332 9774
rect 32172 10164 32228 10174
rect 31500 9268 31556 9278
rect 31500 9174 31556 9212
rect 31052 9156 31108 9166
rect 31052 9062 31108 9100
rect 30716 9044 30772 9054
rect 30716 8950 30772 8988
rect 31612 9042 31668 9054
rect 31612 8990 31614 9042
rect 31666 8990 31668 9042
rect 31500 8820 31556 8830
rect 31500 8726 31556 8764
rect 31612 8484 31668 8990
rect 32172 9042 32228 10108
rect 32844 9826 32900 12124
rect 33068 11506 33124 12348
rect 33068 11454 33070 11506
rect 33122 11454 33124 11506
rect 33068 11442 33124 11454
rect 33404 11508 33460 12796
rect 33964 11732 34020 16606
rect 34524 16658 34580 16670
rect 34524 16606 34526 16658
rect 34578 16606 34580 16658
rect 34300 15202 34356 15214
rect 34300 15150 34302 15202
rect 34354 15150 34356 15202
rect 34188 15092 34244 15102
rect 34188 13746 34244 15036
rect 34300 14644 34356 15150
rect 34524 15204 34580 16606
rect 34972 16658 35028 16670
rect 34972 16606 34974 16658
rect 35026 16606 35028 16658
rect 34524 15092 34916 15148
rect 34300 14578 34356 14588
rect 34636 14084 34692 14094
rect 34188 13694 34190 13746
rect 34242 13694 34244 13746
rect 34188 13682 34244 13694
rect 34412 13972 34468 13982
rect 34412 13746 34468 13916
rect 34636 13970 34692 14028
rect 34636 13918 34638 13970
rect 34690 13918 34692 13970
rect 34636 13906 34692 13918
rect 34860 13970 34916 15092
rect 34860 13918 34862 13970
rect 34914 13918 34916 13970
rect 34860 13906 34916 13918
rect 34412 13694 34414 13746
rect 34466 13694 34468 13746
rect 34412 13682 34468 13694
rect 34748 13636 34804 13646
rect 34748 13542 34804 13580
rect 34972 13412 35028 16606
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35308 16098 35364 16110
rect 35308 16046 35310 16098
rect 35362 16046 35364 16098
rect 35308 15876 35364 16046
rect 35308 15810 35364 15820
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35532 14756 35588 14766
rect 35532 14642 35588 14700
rect 35532 14590 35534 14642
rect 35586 14590 35588 14642
rect 35532 14578 35588 14590
rect 35308 14532 35364 14542
rect 35364 14476 35476 14532
rect 35308 14466 35364 14476
rect 35420 13972 35476 14476
rect 35532 13972 35588 13982
rect 35420 13970 35588 13972
rect 35420 13918 35534 13970
rect 35586 13918 35588 13970
rect 35420 13916 35588 13918
rect 35532 13906 35588 13916
rect 34972 13346 35028 13356
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 34860 13188 34916 13198
rect 35644 13188 35700 18396
rect 35756 17444 35812 17454
rect 35756 17350 35812 17388
rect 35868 17332 35924 18844
rect 36540 18676 36596 21534
rect 36764 21586 36820 21598
rect 36764 21534 36766 21586
rect 36818 21534 36820 21586
rect 36764 21364 36820 21534
rect 36764 21298 36820 21308
rect 36316 18620 36596 18676
rect 35868 17266 35924 17276
rect 35980 18452 36036 18462
rect 35756 16996 35812 17006
rect 35756 16902 35812 16940
rect 35868 14532 35924 14542
rect 35980 14532 36036 18396
rect 36092 18340 36148 18350
rect 36092 18246 36148 18284
rect 36204 18004 36260 18014
rect 36092 17892 36148 17902
rect 36092 17554 36148 17836
rect 36092 17502 36094 17554
rect 36146 17502 36148 17554
rect 36092 17490 36148 17502
rect 36204 16884 36260 17948
rect 36316 17556 36372 18620
rect 36876 18564 36932 22428
rect 37100 22260 37156 22270
rect 36988 22204 37100 22260
rect 36988 21812 37044 22204
rect 37100 22166 37156 22204
rect 37212 22258 37268 22270
rect 37212 22206 37214 22258
rect 37266 22206 37268 22258
rect 36988 20804 37044 21756
rect 37212 22148 37268 22206
rect 37100 21586 37156 21598
rect 37100 21534 37102 21586
rect 37154 21534 37156 21586
rect 37100 21028 37156 21534
rect 37212 21476 37268 22092
rect 37324 22258 37380 22876
rect 37324 22206 37326 22258
rect 37378 22206 37380 22258
rect 37324 21924 37380 22206
rect 37324 21858 37380 21868
rect 37548 21812 37604 23214
rect 37548 21746 37604 21756
rect 37548 21586 37604 21598
rect 37548 21534 37550 21586
rect 37602 21534 37604 21586
rect 37212 21420 37380 21476
rect 37100 20972 37268 21028
rect 37100 20804 37156 20814
rect 37044 20802 37156 20804
rect 37044 20750 37102 20802
rect 37154 20750 37156 20802
rect 37044 20748 37156 20750
rect 36988 20710 37044 20748
rect 37100 20738 37156 20748
rect 36876 18498 36932 18508
rect 36988 20132 37044 20142
rect 36428 18452 36484 18462
rect 36428 18450 36708 18452
rect 36428 18398 36430 18450
rect 36482 18398 36708 18450
rect 36428 18396 36708 18398
rect 36428 18386 36484 18396
rect 36540 18228 36596 18238
rect 36540 18134 36596 18172
rect 36316 17490 36372 17500
rect 36092 16828 36260 16884
rect 36428 17444 36484 17454
rect 36092 14642 36148 16828
rect 36428 16660 36484 17388
rect 36540 16996 36596 17006
rect 36540 16882 36596 16940
rect 36540 16830 36542 16882
rect 36594 16830 36596 16882
rect 36540 16818 36596 16830
rect 36652 16882 36708 18396
rect 36988 18450 37044 20076
rect 36988 18398 36990 18450
rect 37042 18398 37044 18450
rect 36988 18340 37044 18398
rect 36988 18274 37044 18284
rect 37100 18226 37156 18238
rect 37100 18174 37102 18226
rect 37154 18174 37156 18226
rect 37100 17780 37156 18174
rect 36988 17778 37156 17780
rect 36988 17726 37102 17778
rect 37154 17726 37156 17778
rect 36988 17724 37156 17726
rect 36652 16830 36654 16882
rect 36706 16830 36708 16882
rect 36092 14590 36094 14642
rect 36146 14590 36148 14642
rect 36092 14578 36148 14590
rect 36316 16604 36484 16660
rect 36316 14644 36372 16604
rect 36652 16100 36708 16830
rect 36428 16044 36652 16100
rect 36876 17556 36932 17566
rect 36876 16100 36932 17500
rect 36988 16882 37044 17724
rect 37100 17714 37156 17724
rect 37212 17668 37268 20972
rect 37324 20804 37380 21420
rect 37324 20710 37380 20748
rect 37436 20690 37492 20702
rect 37436 20638 37438 20690
rect 37490 20638 37492 20690
rect 37436 19572 37492 20638
rect 37548 20692 37604 21534
rect 37548 20626 37604 20636
rect 37436 19506 37492 19516
rect 37548 18564 37604 18574
rect 37548 18470 37604 18508
rect 37212 17602 37268 17612
rect 37324 18228 37380 18238
rect 37324 17892 37380 18172
rect 37660 18116 37716 25564
rect 37772 25508 37828 25546
rect 37772 25442 37828 25452
rect 37772 25284 37828 25294
rect 37772 23828 37828 25228
rect 37884 23940 37940 25676
rect 37996 25618 38052 26124
rect 38444 26114 38500 26124
rect 37996 25566 37998 25618
rect 38050 25566 38052 25618
rect 37996 25554 38052 25566
rect 38220 25956 38276 25966
rect 38108 25508 38164 25518
rect 37996 24052 38052 24062
rect 38108 24052 38164 25452
rect 37996 24050 38164 24052
rect 37996 23998 37998 24050
rect 38050 23998 38164 24050
rect 37996 23996 38164 23998
rect 38220 25396 38276 25900
rect 37996 23986 38052 23996
rect 37884 23874 37940 23884
rect 37772 23716 37828 23772
rect 38220 23716 38276 25340
rect 38332 25506 38388 25518
rect 38332 25454 38334 25506
rect 38386 25454 38388 25506
rect 38332 25284 38388 25454
rect 38332 25218 38388 25228
rect 38444 24164 38500 24174
rect 38556 24164 38612 26852
rect 38444 24162 38612 24164
rect 38444 24110 38446 24162
rect 38498 24110 38612 24162
rect 38444 24108 38612 24110
rect 38444 24098 38500 24108
rect 38556 23940 38612 23950
rect 38556 23846 38612 23884
rect 38444 23716 38500 23726
rect 37772 23660 38052 23716
rect 38220 23714 38500 23716
rect 38220 23662 38446 23714
rect 38498 23662 38500 23714
rect 38220 23660 38500 23662
rect 37772 23492 37828 23502
rect 37772 22594 37828 23436
rect 37772 22542 37774 22594
rect 37826 22542 37828 22594
rect 37772 22530 37828 22542
rect 37884 23154 37940 23166
rect 37884 23102 37886 23154
rect 37938 23102 37940 23154
rect 37884 21252 37940 23102
rect 37884 21186 37940 21196
rect 37884 20578 37940 20590
rect 37884 20526 37886 20578
rect 37938 20526 37940 20578
rect 37884 20244 37940 20526
rect 37884 20178 37940 20188
rect 37660 18050 37716 18060
rect 37884 19572 37940 19582
rect 37324 17836 37828 17892
rect 37324 17666 37380 17836
rect 37324 17614 37326 17666
rect 37378 17614 37380 17666
rect 37324 17602 37380 17614
rect 37548 17666 37604 17678
rect 37548 17614 37550 17666
rect 37602 17614 37604 17666
rect 37548 16996 37604 17614
rect 37548 16930 37604 16940
rect 37660 17220 37716 17230
rect 36988 16830 36990 16882
rect 37042 16830 37044 16882
rect 36988 16212 37044 16830
rect 37436 16772 37492 16782
rect 37212 16212 37268 16222
rect 36988 16210 37268 16212
rect 36988 16158 37214 16210
rect 37266 16158 37268 16210
rect 36988 16156 37268 16158
rect 36876 16044 37156 16100
rect 36428 15202 36484 16044
rect 36652 16034 36708 16044
rect 36428 15150 36430 15202
rect 36482 15150 36484 15202
rect 36428 15138 36484 15150
rect 36988 15876 37044 15886
rect 36652 14868 36708 14878
rect 36540 14812 36652 14868
rect 36428 14644 36484 14654
rect 36316 14642 36484 14644
rect 36316 14590 36430 14642
rect 36482 14590 36484 14642
rect 36316 14588 36484 14590
rect 36428 14578 36484 14588
rect 35924 14476 36036 14532
rect 35868 14466 35924 14476
rect 36540 14420 36596 14812
rect 36652 14802 36708 14812
rect 36428 14364 36596 14420
rect 34300 12962 34356 12974
rect 34300 12910 34302 12962
rect 34354 12910 34356 12962
rect 34300 12852 34356 12910
rect 34860 12962 34916 13132
rect 34860 12910 34862 12962
rect 34914 12910 34916 12962
rect 34860 12898 34916 12910
rect 35420 13132 35700 13188
rect 35756 13746 35812 13758
rect 35756 13694 35758 13746
rect 35810 13694 35812 13746
rect 34300 12786 34356 12796
rect 34972 12852 35028 12862
rect 35308 12852 35364 12862
rect 34972 12850 35364 12852
rect 34972 12798 34974 12850
rect 35026 12798 35310 12850
rect 35362 12798 35364 12850
rect 34972 12796 35364 12798
rect 34972 12786 35028 12796
rect 35308 12786 35364 12796
rect 35420 12850 35476 13132
rect 35420 12798 35422 12850
rect 35474 12798 35476 12850
rect 35420 12786 35476 12798
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 33964 11666 34020 11676
rect 33516 11508 33572 11518
rect 33404 11506 33572 11508
rect 33404 11454 33518 11506
rect 33570 11454 33572 11506
rect 33404 11452 33572 11454
rect 33516 11442 33572 11452
rect 33068 11284 33124 11294
rect 33068 10610 33124 11228
rect 33068 10558 33070 10610
rect 33122 10558 33124 10610
rect 33068 10546 33124 10558
rect 33404 11060 33460 11070
rect 32844 9774 32846 9826
rect 32898 9774 32900 9826
rect 32844 9762 32900 9774
rect 32732 9716 32788 9726
rect 32508 9660 32732 9716
rect 32508 9154 32564 9660
rect 32732 9650 32788 9660
rect 32508 9102 32510 9154
rect 32562 9102 32564 9154
rect 32508 9090 32564 9102
rect 32172 8990 32174 9042
rect 32226 8990 32228 9042
rect 32172 8978 32228 8990
rect 33404 9044 33460 11004
rect 35532 11060 35588 13132
rect 35644 12738 35700 12750
rect 35644 12686 35646 12738
rect 35698 12686 35700 12738
rect 35644 11506 35700 12686
rect 35756 12290 35812 13694
rect 36092 13412 36148 13422
rect 36092 13074 36148 13356
rect 36092 13022 36094 13074
rect 36146 13022 36148 13074
rect 36092 13010 36148 13022
rect 36428 13074 36484 14364
rect 36428 13022 36430 13074
rect 36482 13022 36484 13074
rect 36316 12964 36372 12974
rect 36316 12870 36372 12908
rect 36428 12628 36484 13022
rect 36540 13634 36596 13646
rect 36540 13582 36542 13634
rect 36594 13582 36596 13634
rect 36540 13076 36596 13582
rect 36988 13076 37044 15820
rect 37100 14980 37156 16044
rect 37212 15202 37268 16156
rect 37324 16100 37380 16110
rect 37436 16100 37492 16716
rect 37548 16324 37604 16334
rect 37660 16324 37716 17164
rect 37548 16322 37716 16324
rect 37548 16270 37550 16322
rect 37602 16270 37716 16322
rect 37548 16268 37716 16270
rect 37548 16258 37604 16268
rect 37548 16100 37604 16110
rect 37436 16098 37604 16100
rect 37436 16046 37550 16098
rect 37602 16046 37604 16098
rect 37436 16044 37604 16046
rect 37324 16006 37380 16044
rect 37436 15876 37492 15886
rect 37212 15150 37214 15202
rect 37266 15150 37268 15202
rect 37212 15138 37268 15150
rect 37324 15652 37380 15662
rect 37100 14924 37268 14980
rect 37212 14420 37268 14924
rect 36988 13020 37156 13076
rect 36540 13010 36596 13020
rect 36428 12562 36484 12572
rect 36988 12850 37044 12862
rect 36988 12798 36990 12850
rect 37042 12798 37044 12850
rect 35756 12238 35758 12290
rect 35810 12238 35812 12290
rect 35756 12180 35812 12238
rect 35756 12114 35812 12124
rect 36988 11620 37044 12798
rect 37100 12180 37156 13020
rect 37212 12962 37268 14364
rect 37324 13412 37380 15596
rect 37436 14642 37492 15820
rect 37548 15314 37604 16044
rect 37548 15262 37550 15314
rect 37602 15262 37604 15314
rect 37548 15250 37604 15262
rect 37772 15316 37828 17836
rect 37884 16884 37940 19516
rect 37996 19124 38052 23660
rect 38444 23650 38500 23660
rect 38668 23380 38724 27692
rect 38892 27636 38948 31276
rect 38780 27580 38948 27636
rect 39004 31108 39060 31118
rect 38780 25732 38836 27580
rect 38892 26850 38948 26862
rect 38892 26798 38894 26850
rect 38946 26798 38948 26850
rect 38892 26628 38948 26798
rect 38892 26562 38948 26572
rect 39004 25844 39060 31052
rect 39116 30100 39172 30110
rect 39116 30006 39172 30044
rect 39340 29426 39396 31612
rect 39676 31556 39732 31566
rect 39676 31462 39732 31500
rect 39340 29374 39342 29426
rect 39394 29374 39396 29426
rect 39340 29362 39396 29374
rect 39676 30324 39732 30334
rect 39116 28530 39172 28542
rect 39116 28478 39118 28530
rect 39170 28478 39172 28530
rect 39116 27858 39172 28478
rect 39116 27806 39118 27858
rect 39170 27806 39172 27858
rect 39116 27794 39172 27806
rect 39340 27748 39396 27758
rect 39116 27188 39172 27198
rect 39116 25956 39172 27132
rect 39340 27074 39396 27692
rect 39340 27022 39342 27074
rect 39394 27022 39396 27074
rect 39340 26908 39396 27022
rect 39228 26852 39396 26908
rect 39676 26908 39732 30268
rect 39788 30210 39844 30222
rect 39788 30158 39790 30210
rect 39842 30158 39844 30210
rect 39788 27748 39844 30158
rect 40012 29540 40068 31724
rect 40124 29764 40180 33068
rect 40236 30100 40292 34300
rect 40460 33460 40516 33470
rect 40460 32228 40516 33404
rect 40460 32162 40516 32172
rect 40572 31554 40628 31566
rect 40572 31502 40574 31554
rect 40626 31502 40628 31554
rect 40572 30324 40628 31502
rect 40572 30258 40628 30268
rect 40684 30210 40740 34412
rect 40684 30158 40686 30210
rect 40738 30158 40740 30210
rect 40684 30146 40740 30158
rect 40796 34244 40852 34254
rect 40348 30100 40404 30110
rect 40236 30098 40404 30100
rect 40236 30046 40350 30098
rect 40402 30046 40404 30098
rect 40236 30044 40404 30046
rect 40348 30034 40404 30044
rect 40460 30100 40516 30110
rect 40796 30100 40852 34188
rect 40908 34242 40964 34412
rect 40908 34190 40910 34242
rect 40962 34190 40964 34242
rect 40908 34178 40964 34190
rect 41020 33572 41076 34860
rect 41132 34356 41188 35644
rect 41244 35634 41300 35644
rect 41468 35700 41524 37102
rect 41692 36372 41748 36382
rect 41692 36278 41748 36316
rect 41468 35634 41524 35644
rect 41692 35588 41748 35598
rect 41804 35588 41860 39116
rect 41916 37604 41972 39900
rect 42028 38724 42084 38762
rect 42028 38658 42084 38668
rect 42252 38164 42308 40126
rect 42364 39060 42420 40348
rect 42476 39396 42532 41692
rect 42588 41682 42644 41692
rect 42924 41412 42980 42702
rect 43036 41972 43092 41982
rect 43148 41972 43204 44046
rect 43372 43540 43428 45612
rect 43484 45574 43540 45612
rect 43820 45556 43876 46510
rect 43932 47234 43988 47246
rect 43932 47182 43934 47234
rect 43986 47182 43988 47234
rect 43932 45892 43988 47182
rect 44156 46002 44212 47404
rect 44380 46676 44436 46686
rect 44268 46228 44324 46238
rect 44268 46114 44324 46172
rect 44268 46062 44270 46114
rect 44322 46062 44324 46114
rect 44268 46050 44324 46062
rect 44156 45950 44158 46002
rect 44210 45950 44212 46002
rect 44156 45938 44212 45950
rect 43932 45798 43988 45836
rect 44380 45892 44436 46620
rect 44380 45826 44436 45836
rect 43820 45490 43876 45500
rect 43596 44322 43652 44334
rect 43596 44270 43598 44322
rect 43650 44270 43652 44322
rect 43596 44212 43652 44270
rect 43820 44324 43876 44334
rect 43820 44230 43876 44268
rect 43596 44146 43652 44156
rect 44268 44212 44324 44222
rect 44268 44118 44324 44156
rect 43932 44098 43988 44110
rect 43932 44046 43934 44098
rect 43986 44046 43988 44098
rect 43932 43764 43988 44046
rect 44044 44100 44100 44110
rect 44044 44006 44100 44044
rect 43932 43698 43988 43708
rect 43260 43484 43428 43540
rect 44492 43652 44548 43662
rect 44492 43538 44548 43596
rect 44492 43486 44494 43538
rect 44546 43486 44548 43538
rect 43260 42308 43316 43484
rect 44492 43474 44548 43486
rect 43820 43428 43876 43438
rect 43820 43426 44100 43428
rect 43820 43374 43822 43426
rect 43874 43374 44100 43426
rect 43820 43372 44100 43374
rect 43820 43362 43876 43372
rect 43372 43204 43428 43214
rect 43372 42978 43428 43148
rect 43372 42926 43374 42978
rect 43426 42926 43428 42978
rect 43372 42914 43428 42926
rect 44044 42868 44100 43372
rect 44380 43426 44436 43438
rect 44380 43374 44382 43426
rect 44434 43374 44436 43426
rect 44156 43316 44212 43326
rect 44268 43316 44324 43326
rect 44156 43314 44268 43316
rect 44156 43262 44158 43314
rect 44210 43262 44268 43314
rect 44156 43260 44268 43262
rect 44156 43250 44212 43260
rect 44156 42868 44212 42878
rect 44044 42866 44212 42868
rect 44044 42814 44158 42866
rect 44210 42814 44212 42866
rect 44044 42812 44212 42814
rect 44156 42802 44212 42812
rect 43596 42756 43652 42766
rect 43596 42644 43652 42700
rect 44044 42644 44100 42654
rect 43596 42642 44100 42644
rect 43596 42590 43598 42642
rect 43650 42590 44046 42642
rect 44098 42590 44100 42642
rect 43596 42588 44100 42590
rect 43596 42578 43652 42588
rect 44044 42578 44100 42588
rect 43484 42530 43540 42542
rect 43484 42478 43486 42530
rect 43538 42478 43540 42530
rect 43484 42420 43540 42478
rect 43596 42420 43652 42430
rect 43484 42364 43596 42420
rect 43596 42354 43652 42364
rect 43260 42252 43540 42308
rect 43260 42084 43316 42094
rect 43484 42084 43540 42252
rect 44156 42196 44212 42206
rect 44268 42196 44324 43260
rect 44212 42140 44324 42196
rect 44156 42130 44212 42140
rect 43484 42028 43652 42084
rect 43260 41990 43316 42028
rect 43092 41916 43204 41972
rect 43596 41970 43652 42028
rect 43596 41918 43598 41970
rect 43650 41918 43652 41970
rect 43036 41878 43092 41916
rect 43484 41860 43540 41870
rect 42812 41356 42980 41412
rect 43148 41858 43540 41860
rect 43148 41806 43486 41858
rect 43538 41806 43540 41858
rect 43148 41804 43540 41806
rect 42588 40516 42644 40526
rect 42588 40290 42644 40460
rect 42588 40238 42590 40290
rect 42642 40238 42644 40290
rect 42588 40226 42644 40238
rect 42700 40404 42756 40414
rect 42700 39730 42756 40348
rect 42700 39678 42702 39730
rect 42754 39678 42756 39730
rect 42700 39666 42756 39678
rect 42588 39396 42644 39406
rect 42476 39340 42588 39396
rect 42588 39330 42644 39340
rect 42476 39060 42532 39070
rect 42364 39058 42532 39060
rect 42364 39006 42478 39058
rect 42530 39006 42532 39058
rect 42364 39004 42532 39006
rect 42252 38098 42308 38108
rect 41916 37548 42084 37604
rect 41692 35586 41860 35588
rect 41692 35534 41694 35586
rect 41746 35534 41860 35586
rect 41692 35532 41860 35534
rect 41692 35522 41748 35532
rect 41244 35476 41300 35486
rect 41244 35474 41636 35476
rect 41244 35422 41246 35474
rect 41298 35422 41636 35474
rect 41244 35420 41636 35422
rect 41244 35410 41300 35420
rect 41580 35028 41636 35420
rect 41692 35028 41748 35038
rect 41580 35026 41748 35028
rect 41580 34974 41694 35026
rect 41746 34974 41748 35026
rect 41580 34972 41748 34974
rect 41692 34962 41748 34972
rect 41132 34262 41188 34300
rect 41020 33506 41076 33516
rect 41244 33906 41300 33918
rect 41244 33854 41246 33906
rect 41298 33854 41300 33906
rect 41244 33460 41300 33854
rect 41244 33394 41300 33404
rect 41468 33572 41524 33582
rect 40908 33236 40964 33246
rect 40908 32786 40964 33180
rect 40908 32734 40910 32786
rect 40962 32734 40964 32786
rect 40908 32722 40964 32734
rect 41468 32562 41524 33516
rect 41468 32510 41470 32562
rect 41522 32510 41524 32562
rect 41468 32498 41524 32510
rect 41020 32452 41076 32462
rect 41020 32358 41076 32396
rect 40908 32228 40964 32238
rect 40908 30994 40964 32172
rect 41132 31780 41188 31790
rect 41692 31780 41748 31790
rect 41132 31778 41636 31780
rect 41132 31726 41134 31778
rect 41186 31726 41636 31778
rect 41132 31724 41636 31726
rect 41132 31714 41188 31724
rect 41244 31554 41300 31566
rect 41244 31502 41246 31554
rect 41298 31502 41300 31554
rect 40908 30942 40910 30994
rect 40962 30942 40964 30994
rect 40908 30212 40964 30942
rect 41020 30996 41076 31006
rect 41244 30996 41300 31502
rect 41356 31556 41412 31566
rect 41356 31462 41412 31500
rect 41468 31554 41524 31566
rect 41468 31502 41470 31554
rect 41522 31502 41524 31554
rect 41468 31444 41524 31502
rect 41356 30996 41412 31006
rect 41020 30994 41412 30996
rect 41020 30942 41022 30994
rect 41074 30942 41358 30994
rect 41410 30942 41412 30994
rect 41020 30940 41412 30942
rect 41020 30930 41076 30940
rect 41132 30212 41188 30222
rect 40908 30210 41188 30212
rect 40908 30158 41134 30210
rect 41186 30158 41188 30210
rect 40908 30156 41188 30158
rect 41132 30146 41188 30156
rect 41244 30212 41300 30222
rect 40460 30098 40628 30100
rect 40460 30046 40462 30098
rect 40514 30046 40628 30098
rect 40460 30044 40628 30046
rect 40460 30034 40516 30044
rect 40124 29698 40180 29708
rect 40460 29764 40516 29774
rect 40572 29764 40628 30044
rect 40796 30034 40852 30044
rect 41132 29764 41188 29774
rect 40572 29708 41076 29764
rect 40348 29652 40404 29662
rect 40348 29558 40404 29596
rect 40012 29474 40068 29484
rect 39900 29426 39956 29438
rect 39900 29374 39902 29426
rect 39954 29374 39956 29426
rect 39900 28644 39956 29374
rect 39900 28578 39956 28588
rect 40012 29204 40068 29214
rect 39900 27748 39956 27758
rect 39788 27692 39900 27748
rect 39900 27682 39956 27692
rect 40012 27186 40068 29148
rect 40460 28756 40516 29708
rect 41020 29650 41076 29708
rect 41020 29598 41022 29650
rect 41074 29598 41076 29650
rect 41020 29586 41076 29598
rect 41132 29650 41188 29708
rect 41132 29598 41134 29650
rect 41186 29598 41188 29650
rect 41132 29586 41188 29598
rect 40460 28642 40516 28700
rect 40908 29540 40964 29550
rect 40908 29426 40964 29484
rect 40908 29374 40910 29426
rect 40962 29374 40964 29426
rect 40908 28756 40964 29374
rect 41244 28868 41300 30156
rect 41356 29650 41412 30940
rect 41468 30324 41524 31388
rect 41468 30258 41524 30268
rect 41580 30324 41636 31724
rect 41692 31686 41748 31724
rect 41692 31332 41748 31342
rect 41804 31332 41860 35532
rect 41916 37380 41972 37390
rect 41916 37266 41972 37324
rect 41916 37214 41918 37266
rect 41970 37214 41972 37266
rect 41916 34916 41972 37214
rect 41916 34850 41972 34860
rect 42028 34692 42084 37548
rect 42476 36484 42532 39004
rect 42700 38724 42756 38734
rect 42700 37378 42756 38668
rect 42812 37828 42868 41356
rect 42924 41188 42980 41198
rect 42924 40404 42980 41132
rect 42924 40310 42980 40348
rect 43148 40292 43204 41804
rect 43484 41794 43540 41804
rect 43596 41524 43652 41918
rect 43596 41458 43652 41468
rect 43820 41746 43876 41758
rect 43820 41694 43822 41746
rect 43874 41694 43876 41746
rect 43036 40236 43204 40292
rect 43372 40628 43428 40638
rect 42812 37762 42868 37772
rect 42924 38722 42980 38734
rect 42924 38670 42926 38722
rect 42978 38670 42980 38722
rect 42700 37326 42702 37378
rect 42754 37326 42756 37378
rect 42700 37314 42756 37326
rect 42476 36418 42532 36428
rect 42700 37044 42756 37054
rect 42028 34626 42084 34636
rect 42140 36258 42196 36270
rect 42140 36206 42142 36258
rect 42194 36206 42196 36258
rect 42140 34244 42196 36206
rect 42140 34178 42196 34188
rect 42476 34130 42532 34142
rect 42476 34078 42478 34130
rect 42530 34078 42532 34130
rect 42140 33796 42196 33806
rect 42140 32674 42196 33740
rect 42476 33236 42532 34078
rect 42588 33460 42644 33470
rect 42588 33366 42644 33404
rect 42476 33170 42532 33180
rect 42140 32622 42142 32674
rect 42194 32622 42196 32674
rect 42140 32610 42196 32622
rect 42252 31778 42308 31790
rect 42252 31726 42254 31778
rect 42306 31726 42308 31778
rect 42252 31668 42308 31726
rect 42588 31780 42644 31790
rect 42252 31602 42308 31612
rect 42476 31666 42532 31678
rect 42476 31614 42478 31666
rect 42530 31614 42532 31666
rect 41748 31276 41860 31332
rect 42364 31556 42420 31566
rect 41692 31266 41748 31276
rect 41916 30324 41972 30334
rect 41580 30322 41748 30324
rect 41580 30270 41582 30322
rect 41634 30270 41748 30322
rect 41580 30268 41748 30270
rect 41580 30258 41636 30268
rect 41356 29598 41358 29650
rect 41410 29598 41412 29650
rect 41356 29586 41412 29598
rect 41580 29876 41636 29886
rect 41244 28802 41300 28812
rect 41468 29316 41524 29326
rect 40908 28690 40964 28700
rect 40460 28590 40462 28642
rect 40514 28590 40516 28642
rect 40460 28578 40516 28590
rect 41356 28644 41412 28654
rect 40348 28532 40404 28542
rect 40348 28438 40404 28476
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 40012 27122 40068 27134
rect 39676 26852 39956 26908
rect 39228 26290 39284 26852
rect 39228 26238 39230 26290
rect 39282 26238 39284 26290
rect 39228 26226 39284 26238
rect 39788 26402 39844 26414
rect 39788 26350 39790 26402
rect 39842 26350 39844 26402
rect 39676 26178 39732 26190
rect 39676 26126 39678 26178
rect 39730 26126 39732 26178
rect 39564 26066 39620 26078
rect 39564 26014 39566 26066
rect 39618 26014 39620 26066
rect 39116 25900 39284 25956
rect 39004 25788 39172 25844
rect 38780 25676 39060 25732
rect 38892 25396 38948 25406
rect 38892 25302 38948 25340
rect 39004 24050 39060 25676
rect 39004 23998 39006 24050
rect 39058 23998 39060 24050
rect 39004 23986 39060 23998
rect 39004 23716 39060 23726
rect 38892 23380 38948 23390
rect 38668 23324 38892 23380
rect 38892 23286 38948 23324
rect 38220 23268 38276 23278
rect 38220 23174 38276 23212
rect 38332 23156 38388 23166
rect 38332 23062 38388 23100
rect 38892 22596 38948 22606
rect 38892 22502 38948 22540
rect 38332 22370 38388 22382
rect 38556 22372 38612 22382
rect 38332 22318 38334 22370
rect 38386 22318 38388 22370
rect 37996 19058 38052 19068
rect 38108 21924 38164 21934
rect 37996 17220 38052 17230
rect 38108 17220 38164 21868
rect 38220 21476 38276 21486
rect 38220 21382 38276 21420
rect 38332 21252 38388 22318
rect 38220 21196 38388 21252
rect 38444 22370 38612 22372
rect 38444 22318 38558 22370
rect 38610 22318 38612 22370
rect 38444 22316 38612 22318
rect 38220 20020 38276 21196
rect 38332 21028 38388 21038
rect 38444 21028 38500 22316
rect 38556 22306 38612 22316
rect 38332 21026 38500 21028
rect 38332 20974 38334 21026
rect 38386 20974 38500 21026
rect 38332 20972 38500 20974
rect 38332 20962 38388 20972
rect 38332 20804 38388 20814
rect 38332 20710 38388 20748
rect 38220 17668 38276 19964
rect 38444 19012 38500 20972
rect 38668 20804 38724 20814
rect 38668 20710 38724 20748
rect 38444 18946 38500 18956
rect 38556 19124 38612 19134
rect 38332 17668 38388 17678
rect 38220 17666 38388 17668
rect 38220 17614 38334 17666
rect 38386 17614 38388 17666
rect 38220 17612 38388 17614
rect 38332 17602 38388 17612
rect 38444 17668 38500 17678
rect 38052 17164 38164 17220
rect 37996 17154 38052 17164
rect 38444 16884 38500 17612
rect 37884 15538 37940 16828
rect 38220 16828 38500 16884
rect 37884 15486 37886 15538
rect 37938 15486 37940 15538
rect 37884 15474 37940 15486
rect 37996 15876 38052 15886
rect 38220 15876 38276 16828
rect 38556 15986 38612 19068
rect 38668 18562 38724 18574
rect 38668 18510 38670 18562
rect 38722 18510 38724 18562
rect 38668 16100 38724 18510
rect 39004 18116 39060 23660
rect 39116 23492 39172 25788
rect 39228 25732 39284 25900
rect 39228 25666 39284 25676
rect 39564 25508 39620 26014
rect 39564 25442 39620 25452
rect 39676 25284 39732 26126
rect 39788 25620 39844 26350
rect 39788 25554 39844 25564
rect 39228 25228 39732 25284
rect 39228 24834 39284 25228
rect 39228 24782 39230 24834
rect 39282 24782 39284 24834
rect 39228 24770 39284 24782
rect 39900 24050 39956 26852
rect 40236 26628 40292 26638
rect 40236 25508 40292 26572
rect 40348 26178 40404 26190
rect 40348 26126 40350 26178
rect 40402 26126 40404 26178
rect 40348 25732 40404 26126
rect 40348 25666 40404 25676
rect 41132 25844 41188 25854
rect 40908 25620 40964 25630
rect 40348 25508 40404 25518
rect 40236 25506 40404 25508
rect 40236 25454 40350 25506
rect 40402 25454 40404 25506
rect 40236 25452 40404 25454
rect 40348 25442 40404 25452
rect 40796 25508 40852 25518
rect 40796 25414 40852 25452
rect 40684 25396 40740 25406
rect 40460 25282 40516 25294
rect 40460 25230 40462 25282
rect 40514 25230 40516 25282
rect 40012 24724 40068 24734
rect 40012 24630 40068 24668
rect 39900 23998 39902 24050
rect 39954 23998 39956 24050
rect 39900 23986 39956 23998
rect 40236 23828 40292 23838
rect 39452 23714 39508 23726
rect 39452 23662 39454 23714
rect 39506 23662 39508 23714
rect 39452 23548 39508 23662
rect 39452 23492 39732 23548
rect 39116 23426 39172 23436
rect 39676 23156 39732 23492
rect 39228 23042 39284 23054
rect 39228 22990 39230 23042
rect 39282 22990 39284 23042
rect 39228 22820 39284 22990
rect 39676 23044 39732 23100
rect 40124 23044 40180 23054
rect 39676 23042 40180 23044
rect 39676 22990 39678 23042
rect 39730 22990 40126 23042
rect 40178 22990 40180 23042
rect 39676 22988 40180 22990
rect 39676 22978 39732 22988
rect 39228 22484 39284 22764
rect 39228 22418 39284 22428
rect 39564 22372 39620 22382
rect 39564 22370 40068 22372
rect 39564 22318 39566 22370
rect 39618 22318 40068 22370
rect 39564 22316 40068 22318
rect 39564 22306 39620 22316
rect 39228 22260 39284 22270
rect 39228 22166 39284 22204
rect 40012 22258 40068 22316
rect 40012 22206 40014 22258
rect 40066 22206 40068 22258
rect 39900 22148 39956 22158
rect 39676 22146 39956 22148
rect 39676 22094 39902 22146
rect 39954 22094 39956 22146
rect 39676 22092 39956 22094
rect 39452 21476 39508 21486
rect 39340 21252 39396 21262
rect 39228 20802 39284 20814
rect 39228 20750 39230 20802
rect 39282 20750 39284 20802
rect 39228 20580 39284 20750
rect 39228 19124 39284 20524
rect 39228 19058 39284 19068
rect 39004 18050 39060 18060
rect 38892 17666 38948 17678
rect 38892 17614 38894 17666
rect 38946 17614 38948 17666
rect 38892 17556 38948 17614
rect 39004 17668 39060 17706
rect 39004 17602 39060 17612
rect 39340 17556 39396 21196
rect 39452 20914 39508 21420
rect 39452 20862 39454 20914
rect 39506 20862 39508 20914
rect 39452 20850 39508 20862
rect 39676 20804 39732 22092
rect 39900 22082 39956 22092
rect 39900 21924 39956 21934
rect 39676 20710 39732 20748
rect 39788 20802 39844 20814
rect 39788 20750 39790 20802
rect 39842 20750 39844 20802
rect 39564 20692 39620 20702
rect 39564 19122 39620 20636
rect 39676 20356 39732 20366
rect 39676 20132 39732 20300
rect 39676 20066 39732 20076
rect 39564 19070 39566 19122
rect 39618 19070 39620 19122
rect 39564 17666 39620 19070
rect 39564 17614 39566 17666
rect 39618 17614 39620 17666
rect 39564 17602 39620 17614
rect 39788 17668 39844 20750
rect 39900 18116 39956 21868
rect 40012 21476 40068 22206
rect 40124 21812 40180 22988
rect 40236 22372 40292 23772
rect 40348 23716 40404 23726
rect 40348 23622 40404 23660
rect 40236 21924 40292 22316
rect 40236 21858 40292 21868
rect 40124 21746 40180 21756
rect 40348 21476 40404 21486
rect 40012 21474 40404 21476
rect 40012 21422 40350 21474
rect 40402 21422 40404 21474
rect 40012 21420 40404 21422
rect 40348 21410 40404 21420
rect 40124 21252 40180 21262
rect 40460 21252 40516 25230
rect 40684 24050 40740 25340
rect 40684 23998 40686 24050
rect 40738 23998 40740 24050
rect 40684 23986 40740 23998
rect 40908 23266 40964 25564
rect 41020 23716 41076 23726
rect 41020 23378 41076 23660
rect 41020 23326 41022 23378
rect 41074 23326 41076 23378
rect 41020 23314 41076 23326
rect 41132 23378 41188 25788
rect 41356 25508 41412 28588
rect 41468 26178 41524 29260
rect 41580 28754 41636 29820
rect 41692 28980 41748 30268
rect 41916 29988 41972 30268
rect 42028 30212 42084 30222
rect 42252 30212 42308 30222
rect 42028 30210 42308 30212
rect 42028 30158 42030 30210
rect 42082 30158 42254 30210
rect 42306 30158 42308 30210
rect 42028 30156 42308 30158
rect 42028 30146 42084 30156
rect 42252 30146 42308 30156
rect 41916 29932 42084 29988
rect 41916 29316 41972 29326
rect 41916 29222 41972 29260
rect 41804 29204 41860 29214
rect 41804 29110 41860 29148
rect 41692 28914 41748 28924
rect 41580 28702 41582 28754
rect 41634 28702 41636 28754
rect 41580 28690 41636 28702
rect 41468 26126 41470 26178
rect 41522 26126 41524 26178
rect 41468 26114 41524 26126
rect 41356 25442 41412 25452
rect 41916 25508 41972 25518
rect 41916 25394 41972 25452
rect 41916 25342 41918 25394
rect 41970 25342 41972 25394
rect 41916 25330 41972 25342
rect 42028 25396 42084 29932
rect 42364 29538 42420 31500
rect 42476 30436 42532 31614
rect 42588 31106 42644 31724
rect 42588 31054 42590 31106
rect 42642 31054 42644 31106
rect 42588 31042 42644 31054
rect 42700 30884 42756 36988
rect 42812 36484 42868 36494
rect 42812 36370 42868 36428
rect 42812 36318 42814 36370
rect 42866 36318 42868 36370
rect 42812 36306 42868 36318
rect 42924 36036 42980 38670
rect 42924 35970 42980 35980
rect 43036 34356 43092 40236
rect 43148 40068 43204 40078
rect 43148 39618 43204 40012
rect 43372 39730 43428 40572
rect 43820 40516 43876 41694
rect 44044 41748 44100 41758
rect 44044 41298 44100 41692
rect 44268 41748 44324 41758
rect 44268 41654 44324 41692
rect 44380 41636 44436 43374
rect 44492 42980 44548 42990
rect 44492 41970 44548 42924
rect 44492 41918 44494 41970
rect 44546 41918 44548 41970
rect 44492 41906 44548 41918
rect 44380 41570 44436 41580
rect 44044 41246 44046 41298
rect 44098 41246 44100 41298
rect 44044 41234 44100 41246
rect 44268 41300 44324 41310
rect 44268 41186 44324 41244
rect 44268 41134 44270 41186
rect 44322 41134 44324 41186
rect 44268 41122 44324 41134
rect 43820 40450 43876 40460
rect 43932 41074 43988 41086
rect 43932 41022 43934 41074
rect 43986 41022 43988 41074
rect 43932 40180 43988 41022
rect 44604 40964 44660 47516
rect 44828 47458 44884 47516
rect 44828 47406 44830 47458
rect 44882 47406 44884 47458
rect 44828 47394 44884 47406
rect 45612 47458 45668 47470
rect 45612 47406 45614 47458
rect 45666 47406 45668 47458
rect 45276 47348 45332 47358
rect 45052 47346 45332 47348
rect 45052 47294 45278 47346
rect 45330 47294 45332 47346
rect 45052 47292 45332 47294
rect 45052 46786 45108 47292
rect 45276 47282 45332 47292
rect 45052 46734 45054 46786
rect 45106 46734 45108 46786
rect 45052 46722 45108 46734
rect 45388 46116 45444 46126
rect 45276 45892 45332 45902
rect 44940 45778 44996 45790
rect 44940 45726 44942 45778
rect 44994 45726 44996 45778
rect 44828 45668 44884 45678
rect 44828 45574 44884 45612
rect 44940 44324 44996 45726
rect 45276 45218 45332 45836
rect 45276 45166 45278 45218
rect 45330 45166 45332 45218
rect 45276 45154 45332 45166
rect 45388 45890 45444 46060
rect 45388 45838 45390 45890
rect 45442 45838 45444 45890
rect 45388 44772 45444 45838
rect 45612 45666 45668 47406
rect 45836 47458 45892 47470
rect 46396 47460 46452 47470
rect 45836 47406 45838 47458
rect 45890 47406 45892 47458
rect 45612 45614 45614 45666
rect 45666 45614 45668 45666
rect 45612 45602 45668 45614
rect 45724 47236 45780 47246
rect 45724 45890 45780 47180
rect 45836 46228 45892 47406
rect 46284 47458 46452 47460
rect 46284 47406 46398 47458
rect 46450 47406 46452 47458
rect 46284 47404 46452 47406
rect 46172 47236 46228 47246
rect 46172 47142 46228 47180
rect 45836 46162 45892 46172
rect 45724 45838 45726 45890
rect 45778 45838 45780 45890
rect 45724 45220 45780 45838
rect 45836 46004 45892 46014
rect 45836 45890 45892 45948
rect 45836 45838 45838 45890
rect 45890 45838 45892 45890
rect 45836 45826 45892 45838
rect 46284 46002 46340 47404
rect 46396 47394 46452 47404
rect 46844 47348 46900 47358
rect 46284 45950 46286 46002
rect 46338 45950 46340 46002
rect 46284 45668 46340 45950
rect 45724 45154 45780 45164
rect 45836 45612 46340 45668
rect 46732 46004 46788 46014
rect 45836 44772 45892 45612
rect 46620 45220 46676 45230
rect 46060 44884 46116 44894
rect 45388 44706 45444 44716
rect 45612 44716 45892 44772
rect 45948 44772 46004 44782
rect 45612 44434 45668 44716
rect 45612 44382 45614 44434
rect 45666 44382 45668 44434
rect 45612 44370 45668 44382
rect 44940 44258 44996 44268
rect 45836 44324 45892 44334
rect 45836 44230 45892 44268
rect 44828 44210 44884 44222
rect 44828 44158 44830 44210
rect 44882 44158 44884 44210
rect 44828 44100 44884 44158
rect 45052 44212 45108 44222
rect 45108 44156 45556 44212
rect 45052 44118 45108 44156
rect 44828 44034 44884 44044
rect 44940 44098 44996 44110
rect 44940 44046 44942 44098
rect 44994 44046 44996 44098
rect 44716 43764 44772 43774
rect 44716 42980 44772 43708
rect 44828 43540 44884 43550
rect 44940 43540 44996 44046
rect 45500 44098 45556 44156
rect 45500 44046 45502 44098
rect 45554 44046 45556 44098
rect 45500 44034 45556 44046
rect 45948 43652 46004 44716
rect 46060 44324 46116 44828
rect 46620 44660 46676 45164
rect 46508 44324 46564 44334
rect 46060 44322 46452 44324
rect 46060 44270 46062 44322
rect 46114 44270 46452 44322
rect 46060 44268 46452 44270
rect 46060 44258 46116 44268
rect 46172 43652 46228 43662
rect 45948 43650 46228 43652
rect 45948 43598 46174 43650
rect 46226 43598 46228 43650
rect 45948 43596 46228 43598
rect 44940 43484 45668 43540
rect 44828 43446 44884 43484
rect 45052 43316 45108 43326
rect 45052 43222 45108 43260
rect 45388 43314 45444 43326
rect 45388 43262 45390 43314
rect 45442 43262 45444 43314
rect 44828 42980 44884 42990
rect 44716 42978 44884 42980
rect 44716 42926 44830 42978
rect 44882 42926 44884 42978
rect 44716 42924 44884 42926
rect 44716 41972 44772 41982
rect 44716 41878 44772 41916
rect 44828 41186 44884 42924
rect 44940 42978 44996 42990
rect 44940 42926 44942 42978
rect 44994 42926 44996 42978
rect 44940 42084 44996 42926
rect 45388 42980 45444 43262
rect 45388 42886 45444 42924
rect 45612 42980 45668 43484
rect 45836 43426 45892 43438
rect 45836 43374 45838 43426
rect 45890 43374 45892 43426
rect 45836 43316 45892 43374
rect 46172 43428 46228 43596
rect 46172 43362 46228 43372
rect 46396 43316 46452 44268
rect 46508 43540 46564 44268
rect 46620 44322 46676 44604
rect 46620 44270 46622 44322
rect 46674 44270 46676 44322
rect 46620 44258 46676 44270
rect 46732 44322 46788 45948
rect 46732 44270 46734 44322
rect 46786 44270 46788 44322
rect 46732 44258 46788 44270
rect 46732 43540 46788 43550
rect 46564 43538 46788 43540
rect 46564 43486 46734 43538
rect 46786 43486 46788 43538
rect 46564 43484 46788 43486
rect 46508 43474 46564 43484
rect 46732 43474 46788 43484
rect 46508 43316 46564 43326
rect 46396 43314 46564 43316
rect 46396 43262 46510 43314
rect 46562 43262 46564 43314
rect 46396 43260 46564 43262
rect 45612 42978 45780 42980
rect 45612 42926 45614 42978
rect 45666 42926 45780 42978
rect 45612 42924 45780 42926
rect 45612 42914 45668 42924
rect 45052 42644 45108 42654
rect 45052 42550 45108 42588
rect 44940 42018 44996 42028
rect 45052 42420 45108 42430
rect 44828 41134 44830 41186
rect 44882 41134 44884 41186
rect 44828 41122 44884 41134
rect 44940 41860 44996 41870
rect 45052 41860 45108 42364
rect 45724 41970 45780 42924
rect 45724 41918 45726 41970
rect 45778 41918 45780 41970
rect 45724 41906 45780 41918
rect 44940 41858 45108 41860
rect 44940 41806 44942 41858
rect 44994 41806 45108 41858
rect 44940 41804 45108 41806
rect 45276 41860 45332 41870
rect 43932 40114 43988 40124
rect 44044 40908 44660 40964
rect 44716 40964 44772 40974
rect 43372 39678 43374 39730
rect 43426 39678 43428 39730
rect 43372 39666 43428 39678
rect 43708 39732 43764 39742
rect 43148 39566 43150 39618
rect 43202 39566 43204 39618
rect 43148 39554 43204 39566
rect 43484 39620 43540 39630
rect 43260 39508 43316 39518
rect 43260 39414 43316 39452
rect 43372 39060 43428 39070
rect 43484 39060 43540 39564
rect 43708 39618 43764 39676
rect 43708 39566 43710 39618
rect 43762 39566 43764 39618
rect 43708 39554 43764 39566
rect 43596 39060 43652 39070
rect 43484 39058 43652 39060
rect 43484 39006 43598 39058
rect 43650 39006 43652 39058
rect 43484 39004 43652 39006
rect 43372 38836 43428 39004
rect 43596 38994 43652 39004
rect 43484 38836 43540 38846
rect 43932 38836 43988 38846
rect 43372 38834 43988 38836
rect 43372 38782 43486 38834
rect 43538 38782 43934 38834
rect 43986 38782 43988 38834
rect 43372 38780 43988 38782
rect 43484 38770 43540 38780
rect 43932 38770 43988 38780
rect 43708 38162 43764 38174
rect 43708 38110 43710 38162
rect 43762 38110 43764 38162
rect 43708 38052 43764 38110
rect 43708 37986 43764 37996
rect 43484 37380 43540 37390
rect 43484 36482 43540 37324
rect 44044 37044 44100 40908
rect 44716 40870 44772 40908
rect 44940 40628 44996 41804
rect 45276 41766 45332 41804
rect 45500 41746 45556 41758
rect 45500 41694 45502 41746
rect 45554 41694 45556 41746
rect 45500 41636 45556 41694
rect 45500 41570 45556 41580
rect 45388 41524 45444 41534
rect 45388 41186 45444 41468
rect 45388 41134 45390 41186
rect 45442 41134 45444 41186
rect 45388 41122 45444 41134
rect 45500 41188 45556 41198
rect 44604 40572 44996 40628
rect 45052 40962 45108 40974
rect 45052 40910 45054 40962
rect 45106 40910 45108 40962
rect 44156 40404 44212 40414
rect 44156 39730 44212 40348
rect 44156 39678 44158 39730
rect 44210 39678 44212 39730
rect 44156 39666 44212 39678
rect 44268 39284 44324 39294
rect 44268 39058 44324 39228
rect 44604 39172 44660 40572
rect 44940 40180 44996 40190
rect 44940 39620 44996 40124
rect 45052 40068 45108 40910
rect 45276 40962 45332 40974
rect 45276 40910 45278 40962
rect 45330 40910 45332 40962
rect 45276 40628 45332 40910
rect 45276 40562 45332 40572
rect 45052 40012 45332 40068
rect 45052 39620 45108 39630
rect 44940 39618 45108 39620
rect 44940 39566 45054 39618
rect 45106 39566 45108 39618
rect 44940 39564 45108 39566
rect 45052 39554 45108 39564
rect 45276 39618 45332 40012
rect 45276 39566 45278 39618
rect 45330 39566 45332 39618
rect 44828 39508 44884 39518
rect 44828 39414 44884 39452
rect 44716 39396 44772 39406
rect 44716 39302 44772 39340
rect 45164 39284 45220 39294
rect 45276 39284 45332 39566
rect 45388 39620 45444 39630
rect 45388 39526 45444 39564
rect 45220 39228 45332 39284
rect 45164 39218 45220 39228
rect 44604 39116 44772 39172
rect 44268 39006 44270 39058
rect 44322 39006 44324 39058
rect 44268 38994 44324 39006
rect 44156 38836 44212 38846
rect 44156 38742 44212 38780
rect 44380 38834 44436 38846
rect 44380 38782 44382 38834
rect 44434 38782 44436 38834
rect 44156 38164 44212 38174
rect 44156 38070 44212 38108
rect 44380 38052 44436 38782
rect 44604 38834 44660 38846
rect 44604 38782 44606 38834
rect 44658 38782 44660 38834
rect 44604 38612 44660 38782
rect 44604 38546 44660 38556
rect 44380 37986 44436 37996
rect 44268 37828 44324 37838
rect 44044 36978 44100 36988
rect 44156 37826 44324 37828
rect 44156 37774 44270 37826
rect 44322 37774 44324 37826
rect 44156 37772 44324 37774
rect 43484 36430 43486 36482
rect 43538 36430 43540 36482
rect 43484 36418 43540 36430
rect 43596 36932 43652 36942
rect 43596 36370 43652 36876
rect 44156 36596 44212 37772
rect 44268 37762 44324 37772
rect 43596 36318 43598 36370
rect 43650 36318 43652 36370
rect 43596 36306 43652 36318
rect 43708 36540 44212 36596
rect 43148 36260 43204 36270
rect 43148 36166 43204 36204
rect 43708 34356 43764 36540
rect 44044 36370 44100 36382
rect 44044 36318 44046 36370
rect 44098 36318 44100 36370
rect 43820 36260 43876 36270
rect 43820 36258 43988 36260
rect 43820 36206 43822 36258
rect 43874 36206 43988 36258
rect 43820 36204 43988 36206
rect 43820 36194 43876 36204
rect 43820 35140 43876 35150
rect 43820 35026 43876 35084
rect 43820 34974 43822 35026
rect 43874 34974 43876 35026
rect 43820 34962 43876 34974
rect 43932 35028 43988 36204
rect 43932 34962 43988 34972
rect 43932 34356 43988 34366
rect 43036 34300 43204 34356
rect 43708 34300 43876 34356
rect 43036 34132 43092 34142
rect 43036 34038 43092 34076
rect 42812 34018 42868 34030
rect 42812 33966 42814 34018
rect 42866 33966 42868 34018
rect 42812 32564 42868 33966
rect 42812 32498 42868 32508
rect 43148 31892 43204 34300
rect 43708 34132 43764 34142
rect 43820 34132 43876 34300
rect 43932 34262 43988 34300
rect 44044 34244 44100 36318
rect 44044 34178 44100 34188
rect 44156 36258 44212 36270
rect 44156 36206 44158 36258
rect 44210 36206 44212 36258
rect 44156 35138 44212 36206
rect 44380 36258 44436 36270
rect 44380 36206 44382 36258
rect 44434 36206 44436 36258
rect 44380 35252 44436 36206
rect 44380 35186 44436 35196
rect 44156 35086 44158 35138
rect 44210 35086 44212 35138
rect 43820 34076 43988 34132
rect 43708 34038 43764 34076
rect 43708 33908 43764 33918
rect 43372 33572 43428 33582
rect 43372 33346 43428 33516
rect 43708 33458 43764 33852
rect 43708 33406 43710 33458
rect 43762 33406 43764 33458
rect 43708 33394 43764 33406
rect 43372 33294 43374 33346
rect 43426 33294 43428 33346
rect 43372 33282 43428 33294
rect 43820 33122 43876 33134
rect 43820 33070 43822 33122
rect 43874 33070 43876 33122
rect 43148 31826 43204 31836
rect 43484 32564 43540 32574
rect 42924 31778 42980 31790
rect 42924 31726 42926 31778
rect 42978 31726 42980 31778
rect 42924 31444 42980 31726
rect 43036 31666 43092 31678
rect 43036 31614 43038 31666
rect 43090 31614 43092 31666
rect 43036 31556 43092 31614
rect 43036 31490 43092 31500
rect 43148 31556 43204 31566
rect 43148 31554 43428 31556
rect 43148 31502 43150 31554
rect 43202 31502 43428 31554
rect 43148 31500 43428 31502
rect 43148 31490 43204 31500
rect 42924 31378 42980 31388
rect 42700 30818 42756 30828
rect 43260 30436 43316 30446
rect 42476 30380 42980 30436
rect 42588 30212 42644 30222
rect 42812 30212 42868 30222
rect 42476 30156 42588 30212
rect 42644 30210 42868 30212
rect 42644 30158 42814 30210
rect 42866 30158 42868 30210
rect 42644 30156 42868 30158
rect 42476 29650 42532 30156
rect 42588 30146 42644 30156
rect 42812 30146 42868 30156
rect 42924 30212 42980 30380
rect 43260 30322 43316 30380
rect 43260 30270 43262 30322
rect 43314 30270 43316 30322
rect 43260 30258 43316 30270
rect 42924 30210 43092 30212
rect 42924 30158 42926 30210
rect 42978 30158 43092 30210
rect 42924 30156 43092 30158
rect 42924 30146 42980 30156
rect 42700 29986 42756 29998
rect 42700 29934 42702 29986
rect 42754 29934 42756 29986
rect 42700 29876 42756 29934
rect 42700 29810 42756 29820
rect 42812 29988 42868 29998
rect 42476 29598 42478 29650
rect 42530 29598 42532 29650
rect 42476 29586 42532 29598
rect 42700 29652 42756 29662
rect 42812 29652 42868 29932
rect 42700 29650 42868 29652
rect 42700 29598 42702 29650
rect 42754 29598 42868 29650
rect 42700 29596 42868 29598
rect 42700 29586 42756 29596
rect 42364 29486 42366 29538
rect 42418 29486 42420 29538
rect 42364 29474 42420 29486
rect 42924 29428 42980 29438
rect 42924 29334 42980 29372
rect 42812 29316 42868 29326
rect 42140 28980 42196 28990
rect 42140 27188 42196 28924
rect 42588 28642 42644 28654
rect 42588 28590 42590 28642
rect 42642 28590 42644 28642
rect 42588 28532 42644 28590
rect 42140 27186 42532 27188
rect 42140 27134 42142 27186
rect 42194 27134 42532 27186
rect 42140 27132 42532 27134
rect 42140 27122 42196 27132
rect 42476 27074 42532 27132
rect 42476 27022 42478 27074
rect 42530 27022 42532 27074
rect 42476 27010 42532 27022
rect 42588 26908 42644 28476
rect 42812 27186 42868 29260
rect 43036 29092 43092 30156
rect 43372 30100 43428 31500
rect 43484 31218 43540 32508
rect 43484 31166 43486 31218
rect 43538 31166 43540 31218
rect 43484 31154 43540 31166
rect 43820 31668 43876 33070
rect 43820 31108 43876 31612
rect 43596 31052 43876 31108
rect 43484 30996 43540 31006
rect 43484 30434 43540 30940
rect 43484 30382 43486 30434
rect 43538 30382 43540 30434
rect 43484 30370 43540 30382
rect 43596 30994 43652 31052
rect 43596 30942 43598 30994
rect 43650 30942 43652 30994
rect 43372 30034 43428 30044
rect 43596 29876 43652 30942
rect 43932 30996 43988 34076
rect 44044 33906 44100 33918
rect 44044 33854 44046 33906
rect 44098 33854 44100 33906
rect 44044 33796 44100 33854
rect 44044 33730 44100 33740
rect 43932 30930 43988 30940
rect 44044 31106 44100 31118
rect 44044 31054 44046 31106
rect 44098 31054 44100 31106
rect 43932 30322 43988 30334
rect 43932 30270 43934 30322
rect 43986 30270 43988 30322
rect 43596 29810 43652 29820
rect 43708 30210 43764 30222
rect 43708 30158 43710 30210
rect 43762 30158 43764 30210
rect 43036 29036 43540 29092
rect 43148 28868 43204 28878
rect 43148 28774 43204 28812
rect 43036 28642 43092 28654
rect 43036 28590 43038 28642
rect 43090 28590 43092 28642
rect 43036 27748 43092 28590
rect 43148 28532 43204 28542
rect 43148 28438 43204 28476
rect 43036 27692 43204 27748
rect 42812 27134 42814 27186
rect 42866 27134 42868 27186
rect 42812 27122 42868 27134
rect 42364 26852 42644 26908
rect 42028 25330 42084 25340
rect 42140 26516 42196 26526
rect 42140 26290 42196 26460
rect 42140 26238 42142 26290
rect 42194 26238 42196 26290
rect 41468 25284 41524 25294
rect 41356 24948 41412 24958
rect 41468 24948 41524 25228
rect 41356 24946 41524 24948
rect 41356 24894 41358 24946
rect 41410 24894 41524 24946
rect 41356 24892 41524 24894
rect 41916 25172 41972 25182
rect 41356 24882 41412 24892
rect 41580 24836 41636 24846
rect 41580 24742 41636 24780
rect 41692 24836 41748 24846
rect 41692 24834 41860 24836
rect 41692 24782 41694 24834
rect 41746 24782 41860 24834
rect 41692 24780 41860 24782
rect 41692 24770 41748 24780
rect 41468 24722 41524 24734
rect 41468 24670 41470 24722
rect 41522 24670 41524 24722
rect 41468 24612 41524 24670
rect 41468 23548 41524 24556
rect 41804 24612 41860 24780
rect 41916 24834 41972 25116
rect 41916 24782 41918 24834
rect 41970 24782 41972 24834
rect 41916 24770 41972 24782
rect 41804 24546 41860 24556
rect 42028 24052 42084 24062
rect 42028 23604 42084 23996
rect 41468 23492 41636 23548
rect 41132 23326 41134 23378
rect 41186 23326 41188 23378
rect 41132 23314 41188 23326
rect 40908 23214 40910 23266
rect 40962 23214 40964 23266
rect 40908 22596 40964 23214
rect 40908 22530 40964 22540
rect 40684 22370 40740 22382
rect 40684 22318 40686 22370
rect 40738 22318 40740 22370
rect 40684 22260 40740 22318
rect 41356 22372 41412 22382
rect 41356 22370 41524 22372
rect 41356 22318 41358 22370
rect 41410 22318 41524 22370
rect 41356 22316 41524 22318
rect 41356 22306 41412 22316
rect 40684 22194 40740 22204
rect 40908 22146 40964 22158
rect 40908 22094 40910 22146
rect 40962 22094 40964 22146
rect 40908 21588 40964 22094
rect 40908 21522 40964 21532
rect 41356 21812 41412 21822
rect 41356 21586 41412 21756
rect 41356 21534 41358 21586
rect 41410 21534 41412 21586
rect 41020 21476 41076 21486
rect 41020 21474 41300 21476
rect 41020 21422 41022 21474
rect 41074 21422 41300 21474
rect 41020 21420 41300 21422
rect 41020 21410 41076 21420
rect 40124 20914 40180 21196
rect 40124 20862 40126 20914
rect 40178 20862 40180 20914
rect 40124 20850 40180 20862
rect 40348 21196 40516 21252
rect 40908 21362 40964 21374
rect 40908 21310 40910 21362
rect 40962 21310 40964 21362
rect 40348 20802 40404 21196
rect 40908 20804 40964 21310
rect 40348 20750 40350 20802
rect 40402 20750 40404 20802
rect 40348 20738 40404 20750
rect 40572 20748 40964 20804
rect 40460 20692 40516 20702
rect 40124 19908 40180 19918
rect 40124 19906 40404 19908
rect 40124 19854 40126 19906
rect 40178 19854 40404 19906
rect 40124 19852 40404 19854
rect 40124 19842 40180 19852
rect 40348 19684 40404 19852
rect 40348 19618 40404 19628
rect 40236 18452 40292 18462
rect 40236 18358 40292 18396
rect 40460 18340 40516 20636
rect 40460 18274 40516 18284
rect 39900 18060 40292 18116
rect 39788 17602 39844 17612
rect 39900 17892 39956 17902
rect 38892 17490 38948 17500
rect 39116 17500 39396 17556
rect 39116 17442 39172 17500
rect 39116 17390 39118 17442
rect 39170 17390 39172 17442
rect 38892 16996 38948 17006
rect 38668 16034 38724 16044
rect 38780 16660 38836 16670
rect 38556 15934 38558 15986
rect 38610 15934 38612 15986
rect 38444 15876 38500 15886
rect 38556 15876 38612 15934
rect 38220 15820 38388 15876
rect 37772 15314 37940 15316
rect 37772 15262 37774 15314
rect 37826 15262 37940 15314
rect 37772 15260 37940 15262
rect 37772 15250 37828 15260
rect 37436 14590 37438 14642
rect 37490 14590 37492 14642
rect 37436 14578 37492 14590
rect 37660 15092 37716 15102
rect 37548 14532 37604 14542
rect 37324 13346 37380 13356
rect 37436 14418 37492 14430
rect 37436 14366 37438 14418
rect 37490 14366 37492 14418
rect 37212 12910 37214 12962
rect 37266 12910 37268 12962
rect 37212 12898 37268 12910
rect 37324 13076 37380 13086
rect 37324 12738 37380 13020
rect 37324 12686 37326 12738
rect 37378 12686 37380 12738
rect 37324 12674 37380 12686
rect 37100 12086 37156 12124
rect 37324 11844 37380 11854
rect 37436 11844 37492 14366
rect 37548 13188 37604 14476
rect 37548 13122 37604 13132
rect 37660 12962 37716 15036
rect 37884 14308 37940 15260
rect 37996 14530 38052 15820
rect 38108 14644 38164 14654
rect 38108 14550 38164 14588
rect 37996 14478 37998 14530
rect 38050 14478 38052 14530
rect 37996 14466 38052 14478
rect 38220 14530 38276 14542
rect 38220 14478 38222 14530
rect 38274 14478 38276 14530
rect 38220 14308 38276 14478
rect 37884 14252 38276 14308
rect 37660 12910 37662 12962
rect 37714 12910 37716 12962
rect 37660 12898 37716 12910
rect 37380 11788 37492 11844
rect 37884 12738 37940 12750
rect 37884 12686 37886 12738
rect 37938 12686 37940 12738
rect 37324 11778 37380 11788
rect 36988 11564 37716 11620
rect 35644 11454 35646 11506
rect 35698 11454 35700 11506
rect 35644 11442 35700 11454
rect 36428 11394 36484 11406
rect 36428 11342 36430 11394
rect 36482 11342 36484 11394
rect 35756 11284 35812 11294
rect 35532 10994 35588 11004
rect 35644 11228 35756 11284
rect 34076 10724 34132 10734
rect 33964 10668 34076 10724
rect 33516 10610 33572 10622
rect 33516 10558 33518 10610
rect 33570 10558 33572 10610
rect 33516 9940 33572 10558
rect 33516 9874 33572 9884
rect 33516 9716 33572 9726
rect 33516 9622 33572 9660
rect 33964 9268 34020 10668
rect 34076 10630 34132 10668
rect 34972 10724 35028 10734
rect 35196 10724 35252 10734
rect 34972 10630 35028 10668
rect 35084 10722 35252 10724
rect 35084 10670 35198 10722
rect 35250 10670 35252 10722
rect 35084 10668 35252 10670
rect 34412 10612 34468 10622
rect 34412 10518 34468 10556
rect 34524 10610 34580 10622
rect 34524 10558 34526 10610
rect 34578 10558 34580 10610
rect 34188 10498 34244 10510
rect 34188 10446 34190 10498
rect 34242 10446 34244 10498
rect 34188 10164 34244 10446
rect 34188 10098 34244 10108
rect 34524 9940 34580 10558
rect 33964 9212 34468 9268
rect 33852 9156 33908 9166
rect 33852 9062 33908 9100
rect 33964 9154 34020 9212
rect 33964 9102 33966 9154
rect 34018 9102 34020 9154
rect 33964 9090 34020 9102
rect 33404 8988 33572 9044
rect 32060 8818 32116 8830
rect 32060 8766 32062 8818
rect 32114 8766 32116 8818
rect 32060 8428 32116 8766
rect 31612 8418 31668 8428
rect 30044 6804 30100 6814
rect 30156 6804 30212 7420
rect 30604 7382 30660 7420
rect 30716 8372 30772 8382
rect 30716 8260 30772 8316
rect 31948 8372 32116 8428
rect 32396 8820 32452 8830
rect 33404 8820 33460 8830
rect 30940 8260 30996 8270
rect 30716 8258 30996 8260
rect 30716 8206 30942 8258
rect 30994 8206 30996 8258
rect 30716 8204 30996 8206
rect 30492 7362 30548 7374
rect 30492 7310 30494 7362
rect 30546 7310 30548 7362
rect 30492 6916 30548 7310
rect 30604 6916 30660 6926
rect 30492 6914 30660 6916
rect 30492 6862 30606 6914
rect 30658 6862 30660 6914
rect 30492 6860 30660 6862
rect 30604 6850 30660 6860
rect 30044 6802 30324 6804
rect 30044 6750 30046 6802
rect 30098 6750 30324 6802
rect 30044 6748 30324 6750
rect 30044 6738 30100 6748
rect 29932 6526 29934 6578
rect 29986 6526 29988 6578
rect 29932 6514 29988 6526
rect 29260 5122 29428 5124
rect 29260 5070 29262 5122
rect 29314 5070 29428 5122
rect 29260 5068 29428 5070
rect 29260 5058 29316 5068
rect 29596 5012 29652 5022
rect 29596 4918 29652 4956
rect 30268 5012 30324 6748
rect 30380 6690 30436 6702
rect 30380 6638 30382 6690
rect 30434 6638 30436 6690
rect 30380 6580 30436 6638
rect 30380 6514 30436 6524
rect 30492 6468 30548 6478
rect 30492 6374 30548 6412
rect 30716 6244 30772 8204
rect 30940 8194 30996 8204
rect 31612 7700 31668 7710
rect 31052 7476 31108 7486
rect 31052 7382 31108 7420
rect 31612 7474 31668 7644
rect 31612 7422 31614 7474
rect 31666 7422 31668 7474
rect 30828 7252 30884 7262
rect 30828 6916 30884 7196
rect 30828 6822 30884 6860
rect 30380 6188 30772 6244
rect 30940 6804 30996 6814
rect 30380 5346 30436 6188
rect 30716 5796 30772 5806
rect 30380 5294 30382 5346
rect 30434 5294 30436 5346
rect 30380 5282 30436 5294
rect 30492 5794 30772 5796
rect 30492 5742 30718 5794
rect 30770 5742 30772 5794
rect 30492 5740 30772 5742
rect 30492 5122 30548 5740
rect 30716 5730 30772 5740
rect 30828 5236 30884 5246
rect 30940 5236 30996 6748
rect 31276 6690 31332 6702
rect 31276 6638 31278 6690
rect 31330 6638 31332 6690
rect 31276 5908 31332 6638
rect 31276 5842 31332 5852
rect 31388 6244 31444 6254
rect 30828 5234 30996 5236
rect 30828 5182 30830 5234
rect 30882 5182 30996 5234
rect 30828 5180 30996 5182
rect 30828 5170 30884 5180
rect 30492 5070 30494 5122
rect 30546 5070 30548 5122
rect 30492 5058 30548 5070
rect 28140 4900 28196 4910
rect 28140 4806 28196 4844
rect 29708 4900 29764 4910
rect 29708 4806 29764 4844
rect 29820 4898 29876 4910
rect 29820 4846 29822 4898
rect 29874 4846 29876 4898
rect 29820 4788 29876 4846
rect 29820 4722 29876 4732
rect 27580 4338 27860 4340
rect 27580 4286 27582 4338
rect 27634 4286 27860 4338
rect 27580 4284 27860 4286
rect 28028 4452 28084 4462
rect 27580 4274 27636 4284
rect 26908 4172 27524 4228
rect 27468 3666 27524 4172
rect 27468 3614 27470 3666
rect 27522 3614 27524 3666
rect 27468 3602 27524 3614
rect 26236 2380 26404 2436
rect 26236 800 26292 2380
rect 28028 800 28084 4396
rect 30268 4340 30324 4956
rect 31276 5012 31332 5022
rect 30716 4900 30772 4910
rect 30716 4450 30772 4844
rect 30716 4398 30718 4450
rect 30770 4398 30772 4450
rect 30716 4386 30772 4398
rect 31276 4788 31332 4956
rect 31276 4450 31332 4732
rect 31276 4398 31278 4450
rect 31330 4398 31332 4450
rect 31276 4386 31332 4398
rect 28252 4228 28308 4238
rect 30268 4228 30324 4284
rect 31052 4340 31108 4350
rect 31052 4246 31108 4284
rect 30380 4228 30436 4238
rect 30268 4226 30436 4228
rect 30268 4174 30382 4226
rect 30434 4174 30436 4226
rect 30268 4172 30436 4174
rect 28252 4134 28308 4172
rect 30380 4162 30436 4172
rect 31164 4228 31220 4238
rect 31164 4134 31220 4172
rect 30492 3668 30548 3678
rect 30492 3574 30548 3612
rect 31388 3554 31444 6188
rect 31612 5012 31668 7422
rect 31948 7476 32004 8372
rect 32396 8258 32452 8764
rect 32396 8206 32398 8258
rect 32450 8206 32452 8258
rect 32396 8194 32452 8206
rect 32956 8818 33460 8820
rect 32956 8766 33406 8818
rect 33458 8766 33460 8818
rect 32956 8764 33460 8766
rect 32620 8036 32676 8046
rect 31836 6804 31892 6814
rect 31836 5906 31892 6748
rect 31836 5854 31838 5906
rect 31890 5854 31892 5906
rect 31836 5842 31892 5854
rect 31948 5794 32004 7420
rect 32284 8034 32676 8036
rect 32284 7982 32622 8034
rect 32674 7982 32676 8034
rect 32284 7980 32676 7982
rect 32284 7698 32340 7980
rect 32620 7970 32676 7980
rect 32844 8034 32900 8046
rect 32844 7982 32846 8034
rect 32898 7982 32900 8034
rect 32284 7646 32286 7698
rect 32338 7646 32340 7698
rect 32172 7252 32228 7262
rect 32060 7250 32228 7252
rect 32060 7198 32174 7250
rect 32226 7198 32228 7250
rect 32060 7196 32228 7198
rect 32060 6802 32116 7196
rect 32172 7186 32228 7196
rect 32060 6750 32062 6802
rect 32114 6750 32116 6802
rect 32060 6738 32116 6750
rect 32284 6132 32340 7646
rect 32508 7588 32564 7598
rect 32732 7588 32788 7598
rect 32508 7586 32732 7588
rect 32508 7534 32510 7586
rect 32562 7534 32732 7586
rect 32508 7532 32732 7534
rect 32508 7522 32564 7532
rect 32732 7522 32788 7532
rect 32284 6066 32340 6076
rect 31948 5742 31950 5794
rect 32002 5742 32004 5794
rect 31948 5730 32004 5742
rect 32508 5908 32564 5918
rect 32396 5684 32452 5694
rect 32396 5590 32452 5628
rect 31612 4946 31668 4956
rect 32284 4900 32340 4910
rect 32284 4564 32340 4844
rect 32060 4562 32340 4564
rect 32060 4510 32286 4562
rect 32338 4510 32340 4562
rect 32060 4508 32340 4510
rect 31612 4452 31668 4462
rect 31612 4358 31668 4396
rect 31388 3502 31390 3554
rect 31442 3502 31444 3554
rect 31388 3490 31444 3502
rect 31612 3668 31668 3678
rect 29820 3444 29876 3454
rect 28364 3332 28420 3342
rect 28364 3238 28420 3276
rect 29820 800 29876 3388
rect 31612 800 31668 3612
rect 32060 3332 32116 4508
rect 32284 4498 32340 4508
rect 32396 4676 32452 4686
rect 32508 4676 32564 5852
rect 32452 4620 32564 4676
rect 32060 3266 32116 3276
rect 32172 4114 32228 4126
rect 32172 4062 32174 4114
rect 32226 4062 32228 4114
rect 32172 2884 32228 4062
rect 32284 3556 32340 3566
rect 32396 3556 32452 4620
rect 32508 4452 32564 4462
rect 32508 4358 32564 4396
rect 32844 3668 32900 7982
rect 32956 7476 33012 8764
rect 33404 8754 33460 8764
rect 33516 8428 33572 8988
rect 34188 9042 34244 9054
rect 34188 8990 34190 9042
rect 34242 8990 34244 9042
rect 33068 8372 33572 8428
rect 33740 8484 33796 8494
rect 34076 8484 34132 8494
rect 33068 8146 33124 8372
rect 33740 8258 33796 8428
rect 33740 8206 33742 8258
rect 33794 8206 33796 8258
rect 33740 8194 33796 8206
rect 33852 8372 34132 8428
rect 34188 8428 34244 8990
rect 34412 8932 34468 9212
rect 34524 9156 34580 9884
rect 34524 9090 34580 9100
rect 35084 10612 35140 10668
rect 35196 10658 35252 10668
rect 34524 8932 34580 8942
rect 34412 8930 34580 8932
rect 34412 8878 34526 8930
rect 34578 8878 34580 8930
rect 34412 8876 34580 8878
rect 34524 8866 34580 8876
rect 35084 8428 35140 10556
rect 35420 10612 35476 10622
rect 35420 10610 35588 10612
rect 35420 10558 35422 10610
rect 35474 10558 35588 10610
rect 35420 10556 35588 10558
rect 35420 10546 35476 10556
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34188 8372 34356 8428
rect 33068 8094 33070 8146
rect 33122 8094 33124 8146
rect 33068 8082 33124 8094
rect 33180 8148 33236 8158
rect 33180 8054 33236 8092
rect 33292 8036 33348 8046
rect 33180 7588 33236 7598
rect 33180 7494 33236 7532
rect 32956 7382 33012 7420
rect 33292 7474 33348 7980
rect 33628 7588 33684 7598
rect 33628 7494 33684 7532
rect 33292 7422 33294 7474
rect 33346 7422 33348 7474
rect 33292 6804 33348 7422
rect 33852 7364 33908 8372
rect 34076 8148 34132 8158
rect 34076 8146 34244 8148
rect 34076 8094 34078 8146
rect 34130 8094 34244 8146
rect 34076 8092 34244 8094
rect 34076 8082 34132 8092
rect 33964 8036 34020 8046
rect 33964 7942 34020 7980
rect 34076 7586 34132 7598
rect 34076 7534 34078 7586
rect 34130 7534 34132 7586
rect 33964 7364 34020 7374
rect 33852 7362 34020 7364
rect 33852 7310 33966 7362
rect 34018 7310 34020 7362
rect 33852 7308 34020 7310
rect 33964 7298 34020 7308
rect 33292 6738 33348 6748
rect 34076 6580 34132 7534
rect 34188 7588 34244 8092
rect 34188 7028 34244 7532
rect 34300 7476 34356 8372
rect 34972 8372 35140 8428
rect 35532 8428 35588 10556
rect 35644 10610 35700 11228
rect 35756 11218 35812 11228
rect 36428 10948 36484 11342
rect 36988 11394 37044 11406
rect 36988 11342 36990 11394
rect 37042 11342 37044 11394
rect 36988 11060 37044 11342
rect 36988 10994 37044 11004
rect 37100 11396 37156 11406
rect 37324 11396 37380 11406
rect 36428 10882 36484 10892
rect 37100 10834 37156 11340
rect 37100 10782 37102 10834
rect 37154 10782 37156 10834
rect 37100 10770 37156 10782
rect 37212 11340 37324 11396
rect 36652 10724 36708 10734
rect 36652 10630 36708 10668
rect 35644 10558 35646 10610
rect 35698 10558 35700 10610
rect 35644 10276 35700 10558
rect 36092 10610 36148 10622
rect 36092 10558 36094 10610
rect 36146 10558 36148 10610
rect 35756 10500 35812 10510
rect 36092 10500 36148 10558
rect 36316 10612 36372 10622
rect 36316 10518 36372 10556
rect 35756 10498 36148 10500
rect 35756 10446 35758 10498
rect 35810 10446 36148 10498
rect 35756 10444 36148 10446
rect 36540 10498 36596 10510
rect 36540 10446 36542 10498
rect 36594 10446 36596 10498
rect 35756 10434 35812 10444
rect 35644 10220 36148 10276
rect 35644 9940 35700 9950
rect 35644 9846 35700 9884
rect 36092 9714 36148 10220
rect 36428 9828 36484 9838
rect 36428 9734 36484 9772
rect 36092 9662 36094 9714
rect 36146 9662 36148 9714
rect 36092 9650 36148 9662
rect 36540 9156 36596 10446
rect 37212 10164 37268 11340
rect 37324 11330 37380 11340
rect 37548 11396 37604 11406
rect 37548 11302 37604 11340
rect 37548 10948 37604 10958
rect 37548 10612 37604 10892
rect 37100 9940 37156 9950
rect 37100 9826 37156 9884
rect 37100 9774 37102 9826
rect 37154 9774 37156 9826
rect 37100 9762 37156 9774
rect 36652 9156 36708 9166
rect 36540 9154 36708 9156
rect 36540 9102 36654 9154
rect 36706 9102 36708 9154
rect 36540 9100 36708 9102
rect 36652 9090 36708 9100
rect 36988 8484 37044 8494
rect 37212 8484 37268 10108
rect 37436 10610 37604 10612
rect 37436 10558 37550 10610
rect 37602 10558 37604 10610
rect 37436 10556 37604 10558
rect 37436 9042 37492 10556
rect 37548 10546 37604 10556
rect 37548 9940 37604 9950
rect 37660 9940 37716 11564
rect 37548 9938 37716 9940
rect 37548 9886 37550 9938
rect 37602 9886 37716 9938
rect 37548 9884 37716 9886
rect 37548 9874 37604 9884
rect 37436 8990 37438 9042
rect 37490 8990 37492 9042
rect 37436 8978 37492 8990
rect 36988 8482 37268 8484
rect 36988 8430 36990 8482
rect 37042 8430 37268 8482
rect 36988 8428 37268 8430
rect 37660 8428 37716 9884
rect 37884 9828 37940 12686
rect 38220 12740 38276 12750
rect 38220 12646 38276 12684
rect 38332 11396 38388 15820
rect 38500 15820 38612 15876
rect 38668 15876 38724 15886
rect 38444 15810 38500 15820
rect 38668 15782 38724 15820
rect 38556 15652 38612 15662
rect 38556 15426 38612 15596
rect 38668 15540 38724 15550
rect 38780 15540 38836 16604
rect 38892 16098 38948 16940
rect 39116 16548 39172 17390
rect 39116 16482 39172 16492
rect 39452 16884 39508 16894
rect 38892 16046 38894 16098
rect 38946 16046 38948 16098
rect 38892 16034 38948 16046
rect 39452 16098 39508 16828
rect 39452 16046 39454 16098
rect 39506 16046 39508 16098
rect 39452 16034 39508 16046
rect 39564 16770 39620 16782
rect 39564 16718 39566 16770
rect 39618 16718 39620 16770
rect 39116 15986 39172 15998
rect 39116 15934 39118 15986
rect 39170 15934 39172 15986
rect 39116 15876 39172 15934
rect 39564 15876 39620 16718
rect 39116 15820 39508 15876
rect 38668 15538 38836 15540
rect 38668 15486 38670 15538
rect 38722 15486 38836 15538
rect 38668 15484 38836 15486
rect 38892 15540 38948 15550
rect 38668 15474 38724 15484
rect 38892 15446 38948 15484
rect 39340 15540 39396 15550
rect 38556 15374 38558 15426
rect 38610 15374 38612 15426
rect 38556 14980 38612 15374
rect 39228 15428 39284 15466
rect 39228 15362 39284 15372
rect 39340 15426 39396 15484
rect 39340 15374 39342 15426
rect 39394 15374 39396 15426
rect 39340 15362 39396 15374
rect 38780 15316 38836 15326
rect 39452 15316 39508 15820
rect 39564 15810 39620 15820
rect 39676 15764 39732 15774
rect 39676 15426 39732 15708
rect 39900 15652 39956 17836
rect 40236 16212 40292 18060
rect 40348 17780 40404 17790
rect 40572 17780 40628 20748
rect 41020 20690 41076 20702
rect 41020 20638 41022 20690
rect 41074 20638 41076 20690
rect 40348 17778 40628 17780
rect 40348 17726 40350 17778
rect 40402 17726 40628 17778
rect 40348 17724 40628 17726
rect 40684 20580 40740 20590
rect 40348 17714 40404 17724
rect 40572 17556 40628 17566
rect 40684 17556 40740 20524
rect 41020 20356 41076 20638
rect 41020 20290 41076 20300
rect 40908 20244 40964 20254
rect 40908 20018 40964 20188
rect 41244 20242 41300 21420
rect 41356 20580 41412 21534
rect 41356 20514 41412 20524
rect 41468 21364 41524 22316
rect 41580 21476 41636 23492
rect 41692 23492 41748 23502
rect 41692 22482 41748 23436
rect 41804 23380 41860 23390
rect 41804 23286 41860 23324
rect 42028 23378 42084 23548
rect 42028 23326 42030 23378
rect 42082 23326 42084 23378
rect 42028 23314 42084 23326
rect 42140 23044 42196 26238
rect 42252 25172 42308 25182
rect 42252 24610 42308 25116
rect 42252 24558 42254 24610
rect 42306 24558 42308 24610
rect 42252 24546 42308 24558
rect 42140 22988 42308 23044
rect 41692 22430 41694 22482
rect 41746 22430 41748 22482
rect 41692 22418 41748 22430
rect 42140 22372 42196 22382
rect 42140 22278 42196 22316
rect 42252 22148 42308 22988
rect 42140 22092 42308 22148
rect 42028 21588 42084 21598
rect 41804 21476 41860 21486
rect 41580 21474 41860 21476
rect 41580 21422 41806 21474
rect 41858 21422 41860 21474
rect 41580 21420 41860 21422
rect 41244 20190 41246 20242
rect 41298 20190 41300 20242
rect 41244 20178 41300 20190
rect 40908 19966 40910 20018
rect 40962 19966 40964 20018
rect 40908 18450 40964 19966
rect 41132 20020 41188 20030
rect 41132 20018 41300 20020
rect 41132 19966 41134 20018
rect 41186 19966 41300 20018
rect 41132 19964 41300 19966
rect 41132 19954 41188 19964
rect 41020 19796 41076 19806
rect 41020 18674 41076 19740
rect 41020 18622 41022 18674
rect 41074 18622 41076 18674
rect 41020 18610 41076 18622
rect 41244 19460 41300 19964
rect 41356 20018 41412 20030
rect 41356 19966 41358 20018
rect 41410 19966 41412 20018
rect 41356 19796 41412 19966
rect 41356 19730 41412 19740
rect 40908 18398 40910 18450
rect 40962 18398 40964 18450
rect 40908 18386 40964 18398
rect 41132 18450 41188 18462
rect 41132 18398 41134 18450
rect 41186 18398 41188 18450
rect 41132 17892 41188 18398
rect 41132 17826 41188 17836
rect 40628 17500 40740 17556
rect 40348 16884 40404 16894
rect 40348 16790 40404 16828
rect 40236 16156 40516 16212
rect 40236 15988 40292 15998
rect 39676 15374 39678 15426
rect 39730 15374 39732 15426
rect 39676 15362 39732 15374
rect 39788 15596 39956 15652
rect 40012 15986 40292 15988
rect 40012 15934 40238 15986
rect 40290 15934 40292 15986
rect 40012 15932 40292 15934
rect 39788 15316 39844 15596
rect 39452 15260 39620 15316
rect 38780 15148 38836 15260
rect 38556 14914 38612 14924
rect 38668 15092 38836 15148
rect 39340 15204 39396 15214
rect 39228 15092 39284 15102
rect 38556 14532 38612 14542
rect 38556 14438 38612 14476
rect 38668 13634 38724 15092
rect 39228 14998 39284 15036
rect 39004 14868 39060 14878
rect 39060 14812 39172 14868
rect 39004 14802 39060 14812
rect 39004 14532 39060 14542
rect 39004 14438 39060 14476
rect 39116 14530 39172 14812
rect 39116 14478 39118 14530
rect 39170 14478 39172 14530
rect 38892 14420 38948 14430
rect 38892 14326 38948 14364
rect 39116 13972 39172 14478
rect 39340 14084 39396 15148
rect 39564 15148 39620 15260
rect 39788 15250 39844 15260
rect 39900 15428 39956 15438
rect 39564 15092 39732 15148
rect 39564 14530 39620 14542
rect 39564 14478 39566 14530
rect 39618 14478 39620 14530
rect 39564 14420 39620 14478
rect 39564 14354 39620 14364
rect 38668 13582 38670 13634
rect 38722 13582 38724 13634
rect 38668 13570 38724 13582
rect 39004 13916 39172 13972
rect 39228 14028 39396 14084
rect 39676 14084 39732 15092
rect 39900 14532 39956 15372
rect 40012 15202 40068 15932
rect 40236 15922 40292 15932
rect 40012 15150 40014 15202
rect 40066 15150 40068 15202
rect 40012 15138 40068 15150
rect 40348 15876 40404 15886
rect 39900 14476 40180 14532
rect 39788 14308 39844 14318
rect 39788 14214 39844 14252
rect 39900 14306 39956 14318
rect 39900 14254 39902 14306
rect 39954 14254 39956 14306
rect 39900 14084 39956 14254
rect 40012 14308 40068 14318
rect 40012 14214 40068 14252
rect 39676 14028 39956 14084
rect 38668 12964 38724 12974
rect 38668 12870 38724 12908
rect 39004 12852 39060 13916
rect 39116 13746 39172 13758
rect 39116 13694 39118 13746
rect 39170 13694 39172 13746
rect 39116 13300 39172 13694
rect 39116 13234 39172 13244
rect 39004 12786 39060 12796
rect 39228 12628 39284 14028
rect 39340 13860 39396 13870
rect 39676 13860 39732 13870
rect 39340 13858 39676 13860
rect 39340 13806 39342 13858
rect 39394 13806 39676 13858
rect 39340 13804 39676 13806
rect 39340 13794 39396 13804
rect 39676 13766 39732 13804
rect 40012 13860 40068 13870
rect 40124 13860 40180 14476
rect 40236 14420 40292 14430
rect 40236 14306 40292 14364
rect 40236 14254 40238 14306
rect 40290 14254 40292 14306
rect 40236 13972 40292 14254
rect 40348 14196 40404 15820
rect 40348 14130 40404 14140
rect 40460 14308 40516 16156
rect 40348 13972 40404 13982
rect 40236 13916 40348 13972
rect 40012 13858 40180 13860
rect 40012 13806 40014 13858
rect 40066 13806 40180 13858
rect 40012 13804 40180 13806
rect 40012 13794 40068 13804
rect 40236 13748 40292 13758
rect 40236 13654 40292 13692
rect 39788 13634 39844 13646
rect 39788 13582 39790 13634
rect 39842 13582 39844 13634
rect 39788 13300 39844 13582
rect 40348 13524 40404 13916
rect 39452 13244 39844 13300
rect 40236 13468 40404 13524
rect 39452 13074 39508 13244
rect 39452 13022 39454 13074
rect 39506 13022 39508 13074
rect 39452 13010 39508 13022
rect 39004 12572 39284 12628
rect 40012 12740 40068 12750
rect 40236 12740 40292 13468
rect 40068 12684 40292 12740
rect 38332 11330 38388 11340
rect 38780 12180 38836 12190
rect 39004 12180 39060 12572
rect 39116 12404 39172 12414
rect 39172 12348 39284 12404
rect 39116 12338 39172 12348
rect 38780 12178 39060 12180
rect 38780 12126 38782 12178
rect 38834 12126 39060 12178
rect 38780 12124 39060 12126
rect 39228 12178 39284 12348
rect 40012 12402 40068 12684
rect 40012 12350 40014 12402
rect 40066 12350 40068 12402
rect 40012 12338 40068 12350
rect 39564 12180 39620 12190
rect 39228 12126 39230 12178
rect 39282 12126 39284 12178
rect 38108 11282 38164 11294
rect 38108 11230 38110 11282
rect 38162 11230 38164 11282
rect 38108 10948 38164 11230
rect 38108 9828 38164 10892
rect 38220 10498 38276 10510
rect 38220 10446 38222 10498
rect 38274 10446 38276 10498
rect 38220 10052 38276 10446
rect 38220 9986 38276 9996
rect 38332 10164 38388 10174
rect 38220 9828 38276 9838
rect 38108 9826 38276 9828
rect 38108 9774 38222 9826
rect 38274 9774 38276 9826
rect 38108 9772 38276 9774
rect 37884 9042 37940 9772
rect 38220 9762 38276 9772
rect 37884 8990 37886 9042
rect 37938 8990 37940 9042
rect 37884 8978 37940 8990
rect 38332 9042 38388 10108
rect 38668 9940 38724 9950
rect 38780 9940 38836 12124
rect 39228 12114 39284 12126
rect 39452 12124 39564 12180
rect 39116 12068 39172 12078
rect 38332 8990 38334 9042
rect 38386 8990 38388 9042
rect 38332 8978 38388 8990
rect 38444 9884 38668 9940
rect 38724 9884 38836 9940
rect 38892 11956 38948 11966
rect 38444 8932 38500 9884
rect 38668 9846 38724 9884
rect 38892 9268 38948 11900
rect 39004 9716 39060 9726
rect 39004 9622 39060 9660
rect 38556 9212 38948 9268
rect 38556 9044 38612 9212
rect 39116 9156 39172 12012
rect 39340 10052 39396 10062
rect 39340 9266 39396 9996
rect 39340 9214 39342 9266
rect 39394 9214 39396 9266
rect 39340 9202 39396 9214
rect 38780 9100 39172 9156
rect 38780 9044 38836 9100
rect 38556 9042 38836 9044
rect 38556 8990 38782 9042
rect 38834 8990 38836 9042
rect 38556 8988 38836 8990
rect 38444 8866 38500 8876
rect 35532 8372 36036 8428
rect 36988 8418 37044 8428
rect 37660 8372 38164 8428
rect 34524 8258 34580 8270
rect 34524 8206 34526 8258
rect 34578 8206 34580 8258
rect 34524 8036 34580 8206
rect 34524 7970 34580 7980
rect 34748 8034 34804 8046
rect 34748 7982 34750 8034
rect 34802 7982 34804 8034
rect 34748 7812 34804 7982
rect 34748 7746 34804 7756
rect 34972 7586 35028 8372
rect 35980 8306 36036 8316
rect 35308 8260 35364 8270
rect 35084 8148 35140 8158
rect 35084 8054 35140 8092
rect 34972 7534 34974 7586
rect 35026 7534 35028 7586
rect 34748 7476 34804 7486
rect 34860 7476 34916 7486
rect 34300 7474 34860 7476
rect 34300 7422 34750 7474
rect 34802 7422 34860 7474
rect 34300 7420 34860 7422
rect 34748 7410 34804 7420
rect 34300 7252 34356 7262
rect 34300 7158 34356 7196
rect 34188 6972 34356 7028
rect 34300 6916 34356 6972
rect 34748 6916 34804 6926
rect 34300 6914 34804 6916
rect 34300 6862 34750 6914
rect 34802 6862 34804 6914
rect 34300 6860 34804 6862
rect 34188 6804 34244 6814
rect 34300 6804 34356 6860
rect 34748 6850 34804 6860
rect 34188 6802 34356 6804
rect 34188 6750 34190 6802
rect 34242 6750 34356 6802
rect 34188 6748 34356 6750
rect 34188 6738 34244 6748
rect 34524 6692 34580 6702
rect 34524 6598 34580 6636
rect 33852 6524 34132 6580
rect 33740 5794 33796 5806
rect 33740 5742 33742 5794
rect 33794 5742 33796 5794
rect 32956 5124 33012 5134
rect 32956 5030 33012 5068
rect 33740 5122 33796 5742
rect 33740 5070 33742 5122
rect 33794 5070 33796 5122
rect 33740 4676 33796 5070
rect 33852 4900 33908 6524
rect 34860 6468 34916 7420
rect 33852 4834 33908 4844
rect 33964 6412 34916 6468
rect 33740 4610 33796 4620
rect 33964 4562 34020 6412
rect 34300 6132 34356 6142
rect 34076 5684 34132 5694
rect 34076 5346 34132 5628
rect 34076 5294 34078 5346
rect 34130 5294 34132 5346
rect 34076 5282 34132 5294
rect 34188 5124 34244 5134
rect 34300 5124 34356 6076
rect 34412 5124 34468 5134
rect 34748 5124 34804 5134
rect 34300 5122 34748 5124
rect 34300 5070 34414 5122
rect 34466 5070 34748 5122
rect 34300 5068 34748 5070
rect 34972 5124 35028 7534
rect 35308 7362 35364 8204
rect 35868 8260 35924 8270
rect 35868 8166 35924 8204
rect 37100 8260 37156 8270
rect 37100 8166 37156 8204
rect 37548 8258 37604 8270
rect 37548 8206 37550 8258
rect 37602 8206 37604 8258
rect 36316 8148 36372 8158
rect 36316 8054 36372 8092
rect 35420 8036 35476 8046
rect 35980 8036 36036 8046
rect 35420 8034 35812 8036
rect 35420 7982 35422 8034
rect 35474 7982 35812 8034
rect 35420 7980 35812 7982
rect 35420 7970 35476 7980
rect 35308 7310 35310 7362
rect 35362 7310 35364 7362
rect 35308 7298 35364 7310
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35084 6916 35140 6926
rect 35084 6690 35140 6860
rect 35756 6916 35812 7980
rect 35756 6802 35812 6860
rect 35756 6750 35758 6802
rect 35810 6750 35812 6802
rect 35756 6738 35812 6750
rect 35084 6638 35086 6690
rect 35138 6638 35140 6690
rect 35084 6626 35140 6638
rect 35644 6692 35700 6702
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35084 5124 35140 5134
rect 34972 5122 35140 5124
rect 34972 5070 35086 5122
rect 35138 5070 35140 5122
rect 34972 5068 35140 5070
rect 34188 5030 34244 5068
rect 34412 5058 34468 5068
rect 34748 5030 34804 5068
rect 35084 5058 35140 5068
rect 35420 5124 35476 5134
rect 35420 5030 35476 5068
rect 35644 5010 35700 6636
rect 35980 6580 36036 7980
rect 36092 8034 36148 8046
rect 36092 7982 36094 8034
rect 36146 7982 36148 8034
rect 36092 6916 36148 7982
rect 36092 6850 36148 6860
rect 36204 8034 36260 8046
rect 36204 7982 36206 8034
rect 36258 7982 36260 8034
rect 36204 7700 36260 7982
rect 36204 6804 36260 7644
rect 37548 7476 37604 8206
rect 37772 8258 37828 8270
rect 37772 8206 37774 8258
rect 37826 8206 37828 8258
rect 37772 8148 37828 8206
rect 37548 7410 37604 7420
rect 37660 8092 37772 8148
rect 37436 7362 37492 7374
rect 37436 7310 37438 7362
rect 37490 7310 37492 7362
rect 36204 6738 36260 6748
rect 36876 7252 36932 7262
rect 36092 6692 36148 6702
rect 36092 6598 36148 6636
rect 35980 6514 36036 6524
rect 36428 6580 36484 6590
rect 36428 6486 36484 6524
rect 36316 6244 36372 6254
rect 35756 5236 35812 5246
rect 35756 5234 36260 5236
rect 35756 5182 35758 5234
rect 35810 5182 36260 5234
rect 35756 5180 36260 5182
rect 35756 5170 35812 5180
rect 35644 4958 35646 5010
rect 35698 4958 35700 5010
rect 35644 4946 35700 4958
rect 36092 5012 36148 5022
rect 36092 4918 36148 4956
rect 34860 4900 34916 4910
rect 34860 4898 35140 4900
rect 34860 4846 34862 4898
rect 34914 4846 35140 4898
rect 34860 4844 35140 4846
rect 34860 4834 34916 4844
rect 33964 4510 33966 4562
rect 34018 4510 34020 4562
rect 33964 4498 34020 4510
rect 34412 4676 34468 4686
rect 33068 4450 33124 4462
rect 33068 4398 33070 4450
rect 33122 4398 33124 4450
rect 32956 3668 33012 3678
rect 32844 3666 33012 3668
rect 32844 3614 32958 3666
rect 33010 3614 33012 3666
rect 32844 3612 33012 3614
rect 32956 3602 33012 3612
rect 32284 3554 32452 3556
rect 32284 3502 32286 3554
rect 32338 3502 32452 3554
rect 32284 3500 32452 3502
rect 32284 3490 32340 3500
rect 33068 3444 33124 4398
rect 33740 4340 33796 4350
rect 33740 4246 33796 4284
rect 34412 4338 34468 4620
rect 35084 4450 35140 4844
rect 35084 4398 35086 4450
rect 35138 4398 35140 4450
rect 35084 4386 35140 4398
rect 35980 4676 36036 4686
rect 34412 4286 34414 4338
rect 34466 4286 34468 4338
rect 34412 4274 34468 4286
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35196 3780 35252 3790
rect 33068 3378 33124 3388
rect 33404 3668 33460 3678
rect 32172 2818 32228 2828
rect 33404 800 33460 3612
rect 35084 3666 35140 3678
rect 35084 3614 35086 3666
rect 35138 3614 35140 3666
rect 35084 3556 35140 3614
rect 35084 3490 35140 3500
rect 35196 800 35252 3724
rect 35980 3554 36036 4620
rect 36204 4116 36260 5180
rect 36316 5124 36372 6188
rect 36876 6244 36932 7196
rect 36988 6692 37044 6702
rect 36988 6598 37044 6636
rect 36876 6178 36932 6188
rect 37100 6578 37156 6590
rect 37100 6526 37102 6578
rect 37154 6526 37156 6578
rect 36428 5684 36484 5694
rect 36428 5346 36484 5628
rect 36428 5294 36430 5346
rect 36482 5294 36484 5346
rect 36428 5282 36484 5294
rect 36988 5234 37044 5246
rect 36988 5182 36990 5234
rect 37042 5182 37044 5234
rect 36428 5124 36484 5134
rect 36988 5124 37044 5182
rect 36316 5122 37044 5124
rect 36316 5070 36430 5122
rect 36482 5070 37044 5122
rect 36316 5068 37044 5070
rect 36428 5058 36484 5068
rect 37100 4340 37156 6526
rect 37212 4340 37268 4350
rect 37100 4284 37212 4340
rect 37212 4226 37268 4284
rect 37212 4174 37214 4226
rect 37266 4174 37268 4226
rect 37212 4162 37268 4174
rect 36988 4116 37044 4126
rect 36204 4060 36820 4116
rect 36764 3666 36820 4060
rect 36764 3614 36766 3666
rect 36818 3614 36820 3666
rect 36764 3602 36820 3614
rect 35980 3502 35982 3554
rect 36034 3502 36036 3554
rect 35980 3490 36036 3502
rect 36988 800 37044 4060
rect 37436 3220 37492 7310
rect 37548 6804 37604 6814
rect 37548 4338 37604 6748
rect 37660 6802 37716 8092
rect 37772 8082 37828 8092
rect 37884 8036 37940 8046
rect 37884 7942 37940 7980
rect 37884 7588 37940 7598
rect 37660 6750 37662 6802
rect 37714 6750 37716 6802
rect 37660 6738 37716 6750
rect 37772 7476 37828 7486
rect 37772 6690 37828 7420
rect 37772 6638 37774 6690
rect 37826 6638 37828 6690
rect 37772 6626 37828 6638
rect 37884 4452 37940 7532
rect 37884 4386 37940 4396
rect 38108 6132 38164 8372
rect 38556 7586 38612 7598
rect 38556 7534 38558 7586
rect 38610 7534 38612 7586
rect 38220 7474 38276 7486
rect 38220 7422 38222 7474
rect 38274 7422 38276 7474
rect 38220 6804 38276 7422
rect 38556 7364 38612 7534
rect 38220 6738 38276 6748
rect 38444 7308 38556 7364
rect 38332 6578 38388 6590
rect 38332 6526 38334 6578
rect 38386 6526 38388 6578
rect 38332 6468 38388 6526
rect 38108 4452 38164 6076
rect 38220 6412 38332 6468
rect 38220 5124 38276 6412
rect 38332 6402 38388 6412
rect 38332 5908 38388 5918
rect 38444 5908 38500 7308
rect 38556 7298 38612 7308
rect 38668 6132 38724 8988
rect 38780 8978 38836 8988
rect 39228 9042 39284 9054
rect 39228 8990 39230 9042
rect 39282 8990 39284 9042
rect 38892 8932 38948 8942
rect 38780 8258 38836 8270
rect 38780 8206 38782 8258
rect 38834 8206 38836 8258
rect 38780 6916 38836 8206
rect 38892 7698 38948 8876
rect 39228 8820 39284 8990
rect 39452 8820 39508 12124
rect 39564 12086 39620 12124
rect 39788 12178 39844 12190
rect 39788 12126 39790 12178
rect 39842 12126 39844 12178
rect 39676 12066 39732 12078
rect 39676 12014 39678 12066
rect 39730 12014 39732 12066
rect 39564 11844 39620 11854
rect 39564 9154 39620 11788
rect 39564 9102 39566 9154
rect 39618 9102 39620 9154
rect 39564 9090 39620 9102
rect 39676 9042 39732 12014
rect 39788 11844 39844 12126
rect 39788 11778 39844 11788
rect 40348 10498 40404 10510
rect 40348 10446 40350 10498
rect 40402 10446 40404 10498
rect 40348 10388 40404 10446
rect 40348 10322 40404 10332
rect 39788 9716 39844 9726
rect 39844 9660 39956 9716
rect 39788 9650 39844 9660
rect 39676 8990 39678 9042
rect 39730 8990 39732 9042
rect 39676 8978 39732 8990
rect 39228 8764 39732 8820
rect 38892 7646 38894 7698
rect 38946 7646 38948 7698
rect 38892 7634 38948 7646
rect 39228 8036 39284 8046
rect 39452 8036 39508 8046
rect 39228 7474 39284 7980
rect 39228 7422 39230 7474
rect 39282 7422 39284 7474
rect 39228 7410 39284 7422
rect 39340 8034 39508 8036
rect 39340 7982 39454 8034
rect 39506 7982 39508 8034
rect 39340 7980 39508 7982
rect 38780 6860 38948 6916
rect 38668 6066 38724 6076
rect 38780 6692 38836 6702
rect 38668 5908 38724 5918
rect 38444 5906 38724 5908
rect 38444 5854 38670 5906
rect 38722 5854 38724 5906
rect 38444 5852 38724 5854
rect 38332 5814 38388 5852
rect 38668 5842 38724 5852
rect 38780 5796 38836 6636
rect 38780 5730 38836 5740
rect 38892 5684 38948 6860
rect 39116 6130 39172 6142
rect 39116 6078 39118 6130
rect 39170 6078 39172 6130
rect 39004 5908 39060 5918
rect 39004 5814 39060 5852
rect 38892 5628 39060 5684
rect 38220 5058 38276 5068
rect 38108 4386 38164 4396
rect 38780 4900 38836 4910
rect 37548 4286 37550 4338
rect 37602 4286 37604 4338
rect 37548 4274 37604 4286
rect 38556 4116 38612 4126
rect 38556 4022 38612 4060
rect 37436 3154 37492 3164
rect 38780 800 38836 4844
rect 38892 3668 38948 3678
rect 39004 3668 39060 5628
rect 39116 5234 39172 6078
rect 39228 6020 39284 6030
rect 39228 5926 39284 5964
rect 39116 5182 39118 5234
rect 39170 5182 39172 5234
rect 39116 5170 39172 5182
rect 39340 3780 39396 7980
rect 39452 7970 39508 7980
rect 39564 7700 39620 7710
rect 39452 7698 39620 7700
rect 39452 7646 39566 7698
rect 39618 7646 39620 7698
rect 39452 7644 39620 7646
rect 39452 6802 39508 7644
rect 39564 7634 39620 7644
rect 39564 7364 39620 7374
rect 39564 7270 39620 7308
rect 39676 7140 39732 8764
rect 39788 7476 39844 7486
rect 39788 7382 39844 7420
rect 39900 7252 39956 9660
rect 40460 9604 40516 14252
rect 40460 9538 40516 9548
rect 40572 15316 40628 17500
rect 41244 17444 41300 19404
rect 41468 19348 41524 21308
rect 41580 20132 41636 20142
rect 41580 20038 41636 20076
rect 41804 19460 41860 21420
rect 42028 20804 42084 21532
rect 42028 20710 42084 20748
rect 42028 19684 42084 19694
rect 41804 19394 41860 19404
rect 41916 19628 42028 19684
rect 41244 17378 41300 17388
rect 41356 19292 41524 19348
rect 40908 16996 40964 17006
rect 40908 16902 40964 16940
rect 41020 16882 41076 16894
rect 41020 16830 41022 16882
rect 41074 16830 41076 16882
rect 41020 16772 41076 16830
rect 41020 16706 41076 16716
rect 41356 16548 41412 19292
rect 41916 19234 41972 19628
rect 42028 19618 42084 19628
rect 42140 19572 42196 22092
rect 42364 21588 42420 26852
rect 42700 26850 42756 26862
rect 42924 26852 42980 26862
rect 42700 26798 42702 26850
rect 42754 26798 42756 26850
rect 42700 26740 42756 26798
rect 42700 26674 42756 26684
rect 42812 26850 42980 26852
rect 42812 26798 42926 26850
rect 42978 26798 42980 26850
rect 42812 26796 42980 26798
rect 42812 26516 42868 26796
rect 42924 26786 42980 26796
rect 43036 26852 43092 26862
rect 43036 26758 43092 26796
rect 42700 26460 42868 26516
rect 42924 26516 42980 26526
rect 43148 26516 43204 27692
rect 42980 26460 43204 26516
rect 43484 27074 43540 29036
rect 43708 28868 43764 30158
rect 43932 29988 43988 30270
rect 43932 29922 43988 29932
rect 43708 28802 43764 28812
rect 44044 28756 44100 31054
rect 44156 30212 44212 35086
rect 44716 35028 44772 39116
rect 45164 38946 45220 38958
rect 45500 38948 45556 41132
rect 45724 40852 45780 40862
rect 45724 40180 45780 40796
rect 45836 40404 45892 43260
rect 46284 42754 46340 42766
rect 46284 42702 46286 42754
rect 46338 42702 46340 42754
rect 45948 41746 46004 41758
rect 45948 41694 45950 41746
rect 46002 41694 46004 41746
rect 45948 41188 46004 41694
rect 46284 41188 46340 42702
rect 46508 41972 46564 43260
rect 46396 41748 46452 41758
rect 46396 41654 46452 41692
rect 46396 41188 46452 41198
rect 46284 41186 46452 41188
rect 46284 41134 46398 41186
rect 46450 41134 46452 41186
rect 46284 41132 46452 41134
rect 45948 41122 46004 41132
rect 45836 40338 45892 40348
rect 45948 40962 46004 40974
rect 45948 40910 45950 40962
rect 46002 40910 46004 40962
rect 45724 40124 45892 40180
rect 45724 39732 45780 39742
rect 45724 39618 45780 39676
rect 45724 39566 45726 39618
rect 45778 39566 45780 39618
rect 45724 39554 45780 39566
rect 45164 38894 45166 38946
rect 45218 38894 45220 38946
rect 44940 38612 44996 38622
rect 45164 38612 45220 38894
rect 45388 38892 45556 38948
rect 45388 38836 45444 38892
rect 45276 38780 45444 38836
rect 45836 38834 45892 40124
rect 45948 38948 46004 40910
rect 46396 40402 46452 41132
rect 46396 40350 46398 40402
rect 46450 40350 46452 40402
rect 46284 39396 46340 39406
rect 46284 39302 46340 39340
rect 45948 38882 46004 38892
rect 46284 39060 46340 39070
rect 46284 38836 46340 39004
rect 45836 38782 45838 38834
rect 45890 38782 45892 38834
rect 45276 38722 45332 38780
rect 45276 38670 45278 38722
rect 45330 38670 45332 38722
rect 45276 38658 45332 38670
rect 45724 38724 45780 38762
rect 45724 38658 45780 38668
rect 44828 38610 44996 38612
rect 44828 38558 44942 38610
rect 44994 38558 44996 38610
rect 44828 38556 44996 38558
rect 44828 38052 44884 38556
rect 44940 38546 44996 38556
rect 45052 38556 45164 38612
rect 44940 38276 44996 38286
rect 45052 38276 45108 38556
rect 44940 38274 45108 38276
rect 44940 38222 44942 38274
rect 44994 38222 45108 38274
rect 44940 38220 45108 38222
rect 44940 38210 44996 38220
rect 45164 38164 45220 38556
rect 45388 38164 45444 38174
rect 45164 38162 45444 38164
rect 45164 38110 45390 38162
rect 45442 38110 45444 38162
rect 45164 38108 45444 38110
rect 45388 38098 45444 38108
rect 44828 37986 44884 37996
rect 45612 38052 45668 38062
rect 45612 38050 45780 38052
rect 45612 37998 45614 38050
rect 45666 37998 45780 38050
rect 45612 37996 45780 37998
rect 45612 37986 45668 37996
rect 45052 37938 45108 37950
rect 45052 37886 45054 37938
rect 45106 37886 45108 37938
rect 45052 37268 45108 37886
rect 45724 37490 45780 37996
rect 45724 37438 45726 37490
rect 45778 37438 45780 37490
rect 45724 37426 45780 37438
rect 45164 37380 45220 37390
rect 45164 37286 45220 37324
rect 45500 37380 45556 37390
rect 44828 37212 45108 37268
rect 44828 37154 44884 37212
rect 44828 37102 44830 37154
rect 44882 37102 44884 37154
rect 44828 37090 44884 37102
rect 45052 36594 45108 37212
rect 45052 36542 45054 36594
rect 45106 36542 45108 36594
rect 45052 36530 45108 36542
rect 45388 37266 45444 37278
rect 45388 37214 45390 37266
rect 45442 37214 45444 37266
rect 45388 36932 45444 37214
rect 45276 36484 45332 36494
rect 45276 36390 45332 36428
rect 45388 36482 45444 36876
rect 45388 36430 45390 36482
rect 45442 36430 45444 36482
rect 45388 36418 45444 36430
rect 45164 36260 45220 36270
rect 45500 36260 45556 37324
rect 45612 37378 45668 37390
rect 45612 37326 45614 37378
rect 45666 37326 45668 37378
rect 45612 36484 45668 37326
rect 45836 36708 45892 38782
rect 46172 38834 46340 38836
rect 46172 38782 46286 38834
rect 46338 38782 46340 38834
rect 46172 38780 46340 38782
rect 46060 38610 46116 38622
rect 46060 38558 46062 38610
rect 46114 38558 46116 38610
rect 45948 38276 46004 38286
rect 46060 38276 46116 38558
rect 45948 38274 46116 38276
rect 45948 38222 45950 38274
rect 46002 38222 46116 38274
rect 45948 38220 46116 38222
rect 45948 38210 46004 38220
rect 46172 37492 46228 38780
rect 46284 38770 46340 38780
rect 46396 38668 46452 40350
rect 46508 39842 46564 41916
rect 46732 41860 46788 41870
rect 46508 39790 46510 39842
rect 46562 39790 46564 39842
rect 46508 39778 46564 39790
rect 46620 41858 46788 41860
rect 46620 41806 46734 41858
rect 46786 41806 46788 41858
rect 46620 41804 46788 41806
rect 46620 39172 46676 41804
rect 46732 41794 46788 41804
rect 46844 40516 46900 47292
rect 47516 46786 47572 46798
rect 47516 46734 47518 46786
rect 47570 46734 47572 46786
rect 47180 46562 47236 46574
rect 47180 46510 47182 46562
rect 47234 46510 47236 46562
rect 47180 46004 47236 46510
rect 47180 45938 47236 45948
rect 47068 45106 47124 45118
rect 47068 45054 47070 45106
rect 47122 45054 47124 45106
rect 46956 43316 47012 43326
rect 47068 43316 47124 45054
rect 47180 44660 47236 44670
rect 47180 44434 47236 44604
rect 47180 44382 47182 44434
rect 47234 44382 47236 44434
rect 47180 44370 47236 44382
rect 47292 44548 47348 44558
rect 47292 43538 47348 44492
rect 47292 43486 47294 43538
rect 47346 43486 47348 43538
rect 47292 43474 47348 43486
rect 47404 44322 47460 44334
rect 47404 44270 47406 44322
rect 47458 44270 47460 44322
rect 47012 43260 47124 43316
rect 47180 43428 47236 43438
rect 47180 43316 47236 43372
rect 47404 43316 47460 44270
rect 47516 44324 47572 46734
rect 47628 44660 47684 47628
rect 47740 47458 47796 47470
rect 47740 47406 47742 47458
rect 47794 47406 47796 47458
rect 47740 46452 47796 47406
rect 48188 47458 48244 47964
rect 48188 47406 48190 47458
rect 48242 47406 48244 47458
rect 48188 47394 48244 47406
rect 48748 47570 48804 47582
rect 48748 47518 48750 47570
rect 48802 47518 48804 47570
rect 48748 47012 48804 47518
rect 49084 47458 49140 47470
rect 49084 47406 49086 47458
rect 49138 47406 49140 47458
rect 49084 47348 49140 47406
rect 49084 47282 49140 47292
rect 48748 46946 48804 46956
rect 48860 46844 49700 46900
rect 48748 46788 48804 46798
rect 48860 46788 48916 46844
rect 48748 46786 48916 46788
rect 48748 46734 48750 46786
rect 48802 46734 48916 46786
rect 48748 46732 48916 46734
rect 48748 46722 48804 46732
rect 47740 46386 47796 46396
rect 47852 46674 47908 46686
rect 47852 46622 47854 46674
rect 47906 46622 47908 46674
rect 47852 46004 47908 46622
rect 48972 46674 49028 46686
rect 48972 46622 48974 46674
rect 49026 46622 49028 46674
rect 47852 45948 48692 46004
rect 48412 45780 48468 45790
rect 48076 45778 48468 45780
rect 48076 45726 48414 45778
rect 48466 45726 48468 45778
rect 48076 45724 48468 45726
rect 47628 44604 48020 44660
rect 47964 44324 48020 44604
rect 48076 44546 48132 45724
rect 48412 45714 48468 45724
rect 48076 44494 48078 44546
rect 48130 44494 48132 44546
rect 48076 44482 48132 44494
rect 48412 45332 48468 45342
rect 48412 44546 48468 45276
rect 48412 44494 48414 44546
rect 48466 44494 48468 44546
rect 48412 44482 48468 44494
rect 48188 44324 48244 44334
rect 47964 44322 48244 44324
rect 47964 44270 48190 44322
rect 48242 44270 48244 44322
rect 47964 44268 48244 44270
rect 47516 44258 47572 44268
rect 48188 44258 48244 44268
rect 48524 44322 48580 44334
rect 48524 44270 48526 44322
rect 48578 44270 48580 44322
rect 47740 44100 47796 44110
rect 48524 44100 48580 44270
rect 47740 44098 48580 44100
rect 47740 44046 47742 44098
rect 47794 44046 48580 44098
rect 47740 44044 48580 44046
rect 47740 44034 47796 44044
rect 48636 43652 48692 45948
rect 48748 45220 48804 45230
rect 48748 45218 48916 45220
rect 48748 45166 48750 45218
rect 48802 45166 48916 45218
rect 48748 45164 48916 45166
rect 48748 45154 48804 45164
rect 48860 44546 48916 45164
rect 48860 44494 48862 44546
rect 48914 44494 48916 44546
rect 48860 44482 48916 44494
rect 48972 43876 49028 46622
rect 49084 45892 49140 45902
rect 49084 45798 49140 45836
rect 49084 45106 49140 45118
rect 49084 45054 49086 45106
rect 49138 45054 49140 45106
rect 49084 44324 49140 45054
rect 49308 44548 49364 44558
rect 49308 44546 49588 44548
rect 49308 44494 49310 44546
rect 49362 44494 49588 44546
rect 49308 44492 49588 44494
rect 49308 44482 49364 44492
rect 49084 44268 49476 44324
rect 49196 44100 49252 44110
rect 49196 44098 49364 44100
rect 49196 44046 49198 44098
rect 49250 44046 49364 44098
rect 49196 44044 49364 44046
rect 49196 44034 49252 44044
rect 48972 43820 49252 43876
rect 47516 43540 47572 43550
rect 47516 43538 47796 43540
rect 47516 43486 47518 43538
rect 47570 43486 47796 43538
rect 47516 43484 47796 43486
rect 47516 43474 47572 43484
rect 47180 43260 47460 43316
rect 47628 43314 47684 43326
rect 47628 43262 47630 43314
rect 47682 43262 47684 43314
rect 46956 43250 47012 43260
rect 47628 42980 47684 43262
rect 47068 42924 47684 42980
rect 47068 42866 47124 42924
rect 47068 42814 47070 42866
rect 47122 42814 47124 42866
rect 47068 42802 47124 42814
rect 47180 42196 47236 42206
rect 47068 42194 47236 42196
rect 47068 42142 47182 42194
rect 47234 42142 47236 42194
rect 47068 42140 47236 42142
rect 47068 41298 47124 42140
rect 47180 42130 47236 42140
rect 47180 41972 47236 41982
rect 47180 41878 47236 41916
rect 47516 41972 47572 41982
rect 47740 41972 47796 43484
rect 47964 43428 48020 43438
rect 47516 41970 47796 41972
rect 47516 41918 47518 41970
rect 47570 41918 47796 41970
rect 47516 41916 47796 41918
rect 47852 43372 47964 43428
rect 47292 41748 47348 41758
rect 47292 41746 47460 41748
rect 47292 41694 47294 41746
rect 47346 41694 47460 41746
rect 47292 41692 47460 41694
rect 47292 41682 47348 41692
rect 47068 41246 47070 41298
rect 47122 41246 47124 41298
rect 47068 41234 47124 41246
rect 47404 40628 47460 41692
rect 47516 40852 47572 41916
rect 47516 40786 47572 40796
rect 47404 40572 47796 40628
rect 46844 40450 46900 40460
rect 47628 40404 47684 40414
rect 47516 40348 47628 40404
rect 47292 40292 47348 40302
rect 46620 39106 46676 39116
rect 46732 40180 46788 40190
rect 46060 37436 46228 37492
rect 46284 38612 46452 38668
rect 46620 38948 46676 38958
rect 46284 38050 46340 38612
rect 46284 37998 46286 38050
rect 46338 37998 46340 38050
rect 45612 36418 45668 36428
rect 45724 36652 45892 36708
rect 45948 37268 46004 37278
rect 45052 35140 45108 35150
rect 44604 34972 44772 35028
rect 44828 35028 44884 35038
rect 44828 35026 44996 35028
rect 44828 34974 44830 35026
rect 44882 34974 44996 35026
rect 44828 34972 44996 34974
rect 44268 34804 44324 34814
rect 44268 34710 44324 34748
rect 44380 34356 44436 34366
rect 44380 34262 44436 34300
rect 44268 32450 44324 32462
rect 44268 32398 44270 32450
rect 44322 32398 44324 32450
rect 44268 32340 44324 32398
rect 44268 32274 44324 32284
rect 44380 32452 44436 32462
rect 44268 31780 44324 31790
rect 44380 31780 44436 32396
rect 44324 31724 44436 31780
rect 44268 31686 44324 31724
rect 44604 31220 44660 34972
rect 44828 34962 44884 34972
rect 44940 34804 44996 34972
rect 44716 34132 44772 34142
rect 44716 34038 44772 34076
rect 44828 33346 44884 33358
rect 44828 33294 44830 33346
rect 44882 33294 44884 33346
rect 44716 32564 44772 32574
rect 44716 32470 44772 32508
rect 44604 31154 44660 31164
rect 44828 31890 44884 33294
rect 44940 33236 44996 34748
rect 45052 33796 45108 35084
rect 45164 34132 45220 36204
rect 45388 36204 45556 36260
rect 45164 34066 45220 34076
rect 45276 35586 45332 35598
rect 45276 35534 45278 35586
rect 45330 35534 45332 35586
rect 45276 34916 45332 35534
rect 45052 33730 45108 33740
rect 45164 33908 45220 33918
rect 45164 33460 45220 33852
rect 45276 33684 45332 34860
rect 45388 34130 45444 36204
rect 45724 35924 45780 36652
rect 45836 36484 45892 36494
rect 45948 36484 46004 37212
rect 46060 36706 46116 37436
rect 46060 36654 46062 36706
rect 46114 36654 46116 36706
rect 46060 36642 46116 36654
rect 45836 36482 46004 36484
rect 45836 36430 45838 36482
rect 45890 36430 46004 36482
rect 45836 36428 46004 36430
rect 45836 36418 45892 36428
rect 45388 34078 45390 34130
rect 45442 34078 45444 34130
rect 45388 34066 45444 34078
rect 45500 34130 45556 34142
rect 45500 34078 45502 34130
rect 45554 34078 45556 34130
rect 45500 34020 45556 34078
rect 45724 34130 45780 35868
rect 45836 35700 45892 35710
rect 45836 35606 45892 35644
rect 45724 34078 45726 34130
rect 45778 34078 45780 34130
rect 45724 34066 45780 34078
rect 45612 34020 45668 34030
rect 45500 33964 45612 34020
rect 45612 33954 45668 33964
rect 45836 33906 45892 33918
rect 45836 33854 45838 33906
rect 45890 33854 45892 33906
rect 45276 33618 45332 33628
rect 45500 33796 45556 33806
rect 45164 33404 45332 33460
rect 45052 33236 45108 33246
rect 44940 33234 45108 33236
rect 44940 33182 45054 33234
rect 45106 33182 45108 33234
rect 44940 33180 45108 33182
rect 44940 33012 44996 33022
rect 44940 32788 44996 32956
rect 45052 32788 45108 33180
rect 45164 33236 45220 33246
rect 45164 33142 45220 33180
rect 45164 32788 45220 32798
rect 45052 32786 45220 32788
rect 45052 32734 45166 32786
rect 45218 32734 45220 32786
rect 45052 32732 45220 32734
rect 44940 32694 44996 32732
rect 45164 32722 45220 32732
rect 45276 32786 45332 33404
rect 45276 32734 45278 32786
rect 45330 32734 45332 32786
rect 45276 32722 45332 32734
rect 45388 33346 45444 33358
rect 45388 33294 45390 33346
rect 45442 33294 45444 33346
rect 45388 32564 45444 33294
rect 45388 32498 45444 32508
rect 45500 32674 45556 33740
rect 45836 33460 45892 33854
rect 45836 33394 45892 33404
rect 45836 33236 45892 33246
rect 45948 33236 46004 36428
rect 46284 36482 46340 37998
rect 46620 37266 46676 38892
rect 46620 37214 46622 37266
rect 46674 37214 46676 37266
rect 46620 36932 46676 37214
rect 46732 37042 46788 40124
rect 47068 40068 47124 40078
rect 47068 39732 47124 40012
rect 47068 39618 47124 39676
rect 47068 39566 47070 39618
rect 47122 39566 47124 39618
rect 47068 39554 47124 39566
rect 47180 39620 47236 39630
rect 47180 39526 47236 39564
rect 46956 39508 47012 39518
rect 46956 39414 47012 39452
rect 47180 39396 47236 39406
rect 47068 38836 47124 38846
rect 47068 38742 47124 38780
rect 47180 38668 47236 39340
rect 47068 38612 47236 38668
rect 47068 38162 47124 38612
rect 47068 38110 47070 38162
rect 47122 38110 47124 38162
rect 47068 38098 47124 38110
rect 46844 37380 46900 37390
rect 46844 37266 46900 37324
rect 46844 37214 46846 37266
rect 46898 37214 46900 37266
rect 46844 37202 46900 37214
rect 46732 36990 46734 37042
rect 46786 36990 46788 37042
rect 46732 36978 46788 36990
rect 46620 36866 46676 36876
rect 47068 36596 47124 36606
rect 47292 36596 47348 40236
rect 47404 39508 47460 39518
rect 47404 39060 47460 39452
rect 47404 38834 47460 39004
rect 47516 38948 47572 40348
rect 47628 40338 47684 40348
rect 47740 39730 47796 40572
rect 47740 39678 47742 39730
rect 47794 39678 47796 39730
rect 47740 39666 47796 39678
rect 47628 39508 47684 39518
rect 47628 39414 47684 39452
rect 47852 39396 47908 43372
rect 47964 43362 48020 43372
rect 48076 43426 48132 43438
rect 48076 43374 48078 43426
rect 48130 43374 48132 43426
rect 48076 43316 48132 43374
rect 48076 43250 48132 43260
rect 48636 42868 48692 43596
rect 48972 43650 49028 43662
rect 48972 43598 48974 43650
rect 49026 43598 49028 43650
rect 48860 43428 48916 43438
rect 48860 43334 48916 43372
rect 48636 42802 48692 42812
rect 48748 43314 48804 43326
rect 48748 43262 48750 43314
rect 48802 43262 48804 43314
rect 48188 41860 48244 41870
rect 48188 41766 48244 41804
rect 48748 40404 48804 43262
rect 48860 42082 48916 42094
rect 48860 42030 48862 42082
rect 48914 42030 48916 42082
rect 48860 40852 48916 42030
rect 48860 40786 48916 40796
rect 48972 40628 49028 43598
rect 49196 43092 49252 43820
rect 48748 40338 48804 40348
rect 48860 40626 49028 40628
rect 48860 40574 48974 40626
rect 49026 40574 49028 40626
rect 48860 40572 49028 40574
rect 48748 40180 48804 40190
rect 48748 40086 48804 40124
rect 47964 40068 48020 40078
rect 47964 39618 48020 40012
rect 48748 39732 48804 39742
rect 48300 39730 48804 39732
rect 48300 39678 48750 39730
rect 48802 39678 48804 39730
rect 48300 39676 48804 39678
rect 47964 39566 47966 39618
rect 48018 39566 48020 39618
rect 47964 39554 48020 39566
rect 48188 39620 48244 39630
rect 48188 39526 48244 39564
rect 47852 39330 47908 39340
rect 47628 38948 47684 38958
rect 47516 38946 47684 38948
rect 47516 38894 47630 38946
rect 47682 38894 47684 38946
rect 47516 38892 47684 38894
rect 47628 38882 47684 38892
rect 47404 38782 47406 38834
rect 47458 38782 47460 38834
rect 47404 38770 47460 38782
rect 48076 38836 48132 38846
rect 48076 38742 48132 38780
rect 48188 38724 48244 38762
rect 48188 38658 48244 38668
rect 47964 37378 48020 37390
rect 47964 37326 47966 37378
rect 48018 37326 48020 37378
rect 47068 36594 47348 36596
rect 47068 36542 47070 36594
rect 47122 36542 47348 36594
rect 47068 36540 47348 36542
rect 47628 37266 47684 37278
rect 47628 37214 47630 37266
rect 47682 37214 47684 37266
rect 47068 36530 47124 36540
rect 46284 36430 46286 36482
rect 46338 36430 46340 36482
rect 46284 36418 46340 36430
rect 47628 36260 47684 37214
rect 47964 37044 48020 37326
rect 47964 36978 48020 36988
rect 47628 36194 47684 36204
rect 48300 35812 48356 39676
rect 48748 39666 48804 39676
rect 48860 39506 48916 40572
rect 48972 40562 49028 40572
rect 49084 43036 49252 43092
rect 48972 40292 49028 40302
rect 48972 40198 49028 40236
rect 49084 39732 49140 43036
rect 49196 42868 49252 42878
rect 49196 42774 49252 42812
rect 49196 41972 49252 41982
rect 49308 41972 49364 44044
rect 49196 41970 49364 41972
rect 49196 41918 49198 41970
rect 49250 41918 49364 41970
rect 49196 41916 49364 41918
rect 49196 41906 49252 41916
rect 49196 41300 49252 41310
rect 49196 41206 49252 41244
rect 49084 39676 49252 39732
rect 48860 39454 48862 39506
rect 48914 39454 48916 39506
rect 48748 38948 48804 38958
rect 48748 38854 48804 38892
rect 48748 37380 48804 37390
rect 48748 37286 48804 37324
rect 48860 37044 48916 39454
rect 49084 39506 49140 39518
rect 49084 39454 49086 39506
rect 49138 39454 49140 39506
rect 49084 39060 49140 39454
rect 48860 36978 48916 36988
rect 48972 39004 49140 39060
rect 47292 35756 48356 35812
rect 48412 36484 48468 36494
rect 47180 35252 47236 35262
rect 46956 34804 47012 34814
rect 46956 34710 47012 34748
rect 47180 34354 47236 35196
rect 47180 34302 47182 34354
rect 47234 34302 47236 34354
rect 47180 34290 47236 34302
rect 47068 34130 47124 34142
rect 47068 34078 47070 34130
rect 47122 34078 47124 34130
rect 46172 34020 46228 34030
rect 46172 33926 46228 33964
rect 46732 34018 46788 34030
rect 46732 33966 46734 34018
rect 46786 33966 46788 34018
rect 46508 33908 46564 33918
rect 46508 33814 46564 33852
rect 45836 33234 46004 33236
rect 45836 33182 45838 33234
rect 45890 33182 46004 33234
rect 45836 33180 46004 33182
rect 46396 33346 46452 33358
rect 46396 33294 46398 33346
rect 46450 33294 46452 33346
rect 45836 33170 45892 33180
rect 46284 32788 46340 32798
rect 45500 32622 45502 32674
rect 45554 32622 45556 32674
rect 45052 32340 45108 32350
rect 44828 31838 44830 31890
rect 44882 31838 44884 31890
rect 44828 31108 44884 31838
rect 44940 31892 44996 31902
rect 44940 31798 44996 31836
rect 44940 31108 44996 31118
rect 44828 31052 44940 31108
rect 44940 31042 44996 31052
rect 45052 30772 45108 32284
rect 45500 32228 45556 32622
rect 45948 32786 46340 32788
rect 45948 32734 46286 32786
rect 46338 32734 46340 32786
rect 45948 32732 46340 32734
rect 45724 32452 45780 32462
rect 45724 32358 45780 32396
rect 45500 32162 45556 32172
rect 45724 32004 45780 32014
rect 45724 31892 45780 31948
rect 45500 31836 45780 31892
rect 44940 30716 45108 30772
rect 45164 31778 45220 31790
rect 45500 31780 45556 31836
rect 45164 31726 45166 31778
rect 45218 31726 45220 31778
rect 44156 30146 44212 30156
rect 44828 30210 44884 30222
rect 44828 30158 44830 30210
rect 44882 30158 44884 30210
rect 44044 28690 44100 28700
rect 44380 29986 44436 29998
rect 44380 29934 44382 29986
rect 44434 29934 44436 29986
rect 44380 28644 44436 29934
rect 44380 28578 44436 28588
rect 44716 29428 44772 29438
rect 44044 28530 44100 28542
rect 44044 28478 44046 28530
rect 44098 28478 44100 28530
rect 44044 27186 44100 28478
rect 44156 28420 44212 28430
rect 44156 28418 44660 28420
rect 44156 28366 44158 28418
rect 44210 28366 44660 28418
rect 44156 28364 44660 28366
rect 44156 28354 44212 28364
rect 44156 27748 44212 27758
rect 44156 27654 44212 27692
rect 44044 27134 44046 27186
rect 44098 27134 44100 27186
rect 44044 27122 44100 27134
rect 43484 27022 43486 27074
rect 43538 27022 43540 27074
rect 42476 26180 42532 26190
rect 42476 26086 42532 26124
rect 42588 24724 42644 24734
rect 42364 21522 42420 21532
rect 42476 24668 42588 24724
rect 42476 21586 42532 24668
rect 42588 24658 42644 24668
rect 42588 23044 42644 23054
rect 42588 22950 42644 22988
rect 42476 21534 42478 21586
rect 42530 21534 42532 21586
rect 42476 21522 42532 21534
rect 42588 22484 42644 22494
rect 42700 22484 42756 26460
rect 42924 26450 42980 26460
rect 43484 26180 43540 27022
rect 43708 26962 43764 26974
rect 43708 26910 43710 26962
rect 43762 26910 43764 26962
rect 43708 26908 43764 26910
rect 43484 26114 43540 26124
rect 43596 26852 43764 26908
rect 43932 26962 43988 26974
rect 43932 26910 43934 26962
rect 43986 26910 43988 26962
rect 43596 26740 43652 26852
rect 42924 25732 42980 25742
rect 42980 25676 43092 25732
rect 42924 25666 42980 25676
rect 42924 25506 42980 25518
rect 42924 25454 42926 25506
rect 42978 25454 42980 25506
rect 42924 25284 42980 25454
rect 42924 25218 42980 25228
rect 43036 24388 43092 25676
rect 43596 25620 43652 26684
rect 43932 25732 43988 26910
rect 43484 25564 43652 25620
rect 43708 25676 43988 25732
rect 44044 26852 44100 26862
rect 43036 24322 43092 24332
rect 43148 25282 43204 25294
rect 43148 25230 43150 25282
rect 43202 25230 43204 25282
rect 42812 23826 42868 23838
rect 42812 23774 42814 23826
rect 42866 23774 42868 23826
rect 42812 23268 42868 23774
rect 43148 23604 43204 25230
rect 43148 23538 43204 23548
rect 43260 25282 43316 25294
rect 43260 25230 43262 25282
rect 43314 25230 43316 25282
rect 42812 23212 43204 23268
rect 42588 22482 42756 22484
rect 42588 22430 42590 22482
rect 42642 22430 42756 22482
rect 42588 22428 42756 22430
rect 42812 23044 42868 23054
rect 42588 22372 42644 22428
rect 42588 21364 42644 22316
rect 42252 21308 42644 21364
rect 42252 20578 42308 21308
rect 42588 20804 42644 20814
rect 42364 20692 42420 20702
rect 42364 20598 42420 20636
rect 42252 20526 42254 20578
rect 42306 20526 42308 20578
rect 42252 20244 42308 20526
rect 42252 20178 42308 20188
rect 42476 20578 42532 20590
rect 42476 20526 42478 20578
rect 42530 20526 42532 20578
rect 42252 19906 42308 19918
rect 42252 19854 42254 19906
rect 42306 19854 42308 19906
rect 42252 19796 42308 19854
rect 42476 19908 42532 20526
rect 42476 19842 42532 19852
rect 42252 19730 42308 19740
rect 42140 19516 42308 19572
rect 41916 19182 41918 19234
rect 41970 19182 41972 19234
rect 41916 18564 41972 19182
rect 41916 18498 41972 18508
rect 42028 18452 42084 18462
rect 42252 18452 42308 19516
rect 42588 19460 42644 20748
rect 42700 20690 42756 20702
rect 42700 20638 42702 20690
rect 42754 20638 42756 20690
rect 42700 19796 42756 20638
rect 42812 20468 42868 22988
rect 43036 22820 43092 22830
rect 42812 20402 42868 20412
rect 42924 22764 43036 22820
rect 42700 19730 42756 19740
rect 42924 19684 42980 22764
rect 43036 22754 43092 22764
rect 43148 22260 43204 23212
rect 43260 22484 43316 25230
rect 43372 25284 43428 25294
rect 43484 25284 43540 25564
rect 43596 25396 43652 25406
rect 43596 25302 43652 25340
rect 43372 25282 43540 25284
rect 43372 25230 43374 25282
rect 43426 25230 43540 25282
rect 43372 25228 43540 25230
rect 43372 24612 43428 25228
rect 43708 24948 43764 25676
rect 43820 25508 43876 25518
rect 43820 25060 43876 25452
rect 43932 25284 43988 25294
rect 44044 25284 44100 26796
rect 44604 26402 44660 28364
rect 44716 27860 44772 29372
rect 44716 27766 44772 27804
rect 44828 28866 44884 30158
rect 44940 30100 44996 30716
rect 45052 30548 45108 30558
rect 45052 30322 45108 30492
rect 45052 30270 45054 30322
rect 45106 30270 45108 30322
rect 45052 30258 45108 30270
rect 45164 30324 45220 31726
rect 45388 31724 45556 31780
rect 45724 31778 45780 31836
rect 45724 31726 45726 31778
rect 45778 31726 45780 31778
rect 45164 30258 45220 30268
rect 45276 30772 45332 30782
rect 45276 30210 45332 30716
rect 45276 30158 45278 30210
rect 45330 30158 45332 30210
rect 45276 30146 45332 30158
rect 45052 30100 45108 30110
rect 44940 30098 45108 30100
rect 44940 30046 45054 30098
rect 45106 30046 45108 30098
rect 44940 30044 45108 30046
rect 44828 28814 44830 28866
rect 44882 28814 44884 28866
rect 44828 27300 44884 28814
rect 45052 28644 45108 30044
rect 45164 28868 45220 28878
rect 45388 28868 45444 31724
rect 45724 31714 45780 31726
rect 45836 31780 45892 31790
rect 45612 31668 45668 31678
rect 45612 31574 45668 31612
rect 45500 31554 45556 31566
rect 45500 31502 45502 31554
rect 45554 31502 45556 31554
rect 45500 30324 45556 31502
rect 45612 31220 45668 31230
rect 45612 31126 45668 31164
rect 45836 31218 45892 31724
rect 45836 31166 45838 31218
rect 45890 31166 45892 31218
rect 45836 31154 45892 31166
rect 45836 30882 45892 30894
rect 45836 30830 45838 30882
rect 45890 30830 45892 30882
rect 45500 30268 45668 30324
rect 45500 30098 45556 30110
rect 45500 30046 45502 30098
rect 45554 30046 45556 30098
rect 45500 29876 45556 30046
rect 45500 29810 45556 29820
rect 45612 29764 45668 30268
rect 45724 29988 45780 29998
rect 45724 29894 45780 29932
rect 45612 29698 45668 29708
rect 45836 29316 45892 30830
rect 45948 30212 46004 32732
rect 46284 32722 46340 32732
rect 46396 32564 46452 33294
rect 46172 32508 46452 32564
rect 46620 32564 46676 32574
rect 46172 31780 46228 32508
rect 46620 32470 46676 32508
rect 46284 32338 46340 32350
rect 46284 32286 46286 32338
rect 46338 32286 46340 32338
rect 46284 32004 46340 32286
rect 46284 31938 46340 31948
rect 46396 32338 46452 32350
rect 46396 32286 46398 32338
rect 46450 32286 46452 32338
rect 46284 31780 46340 31790
rect 46172 31778 46340 31780
rect 46172 31726 46286 31778
rect 46338 31726 46340 31778
rect 46172 31724 46340 31726
rect 46060 30996 46116 31006
rect 46060 30902 46116 30940
rect 46060 30212 46116 30222
rect 45948 30210 46116 30212
rect 45948 30158 46062 30210
rect 46114 30158 46116 30210
rect 45948 30156 46116 30158
rect 46060 30146 46116 30156
rect 45948 29988 46004 29998
rect 45948 29894 46004 29932
rect 46172 29540 46228 31724
rect 46284 31714 46340 31724
rect 46284 30884 46340 30894
rect 46284 30790 46340 30828
rect 46396 30436 46452 32286
rect 46732 31892 46788 33966
rect 47068 33908 47124 34078
rect 47068 33842 47124 33852
rect 47068 33460 47124 33470
rect 47068 33366 47124 33404
rect 47292 33012 47348 35756
rect 48188 35588 48244 35598
rect 48188 35586 48356 35588
rect 48188 35534 48190 35586
rect 48242 35534 48356 35586
rect 48188 35532 48356 35534
rect 48188 35522 48244 35532
rect 47628 35476 47684 35486
rect 47516 35474 47684 35476
rect 47516 35422 47630 35474
rect 47682 35422 47684 35474
rect 47516 35420 47684 35422
rect 47404 34356 47460 34366
rect 47404 34262 47460 34300
rect 47180 32956 47348 33012
rect 47068 32562 47124 32574
rect 47068 32510 47070 32562
rect 47122 32510 47124 32562
rect 47068 32116 47124 32510
rect 46508 31780 46564 31790
rect 46508 31556 46564 31724
rect 46508 30994 46564 31500
rect 46508 30942 46510 30994
rect 46562 30942 46564 30994
rect 46508 30930 46564 30942
rect 46620 31668 46676 31678
rect 46508 30548 46564 30558
rect 46620 30548 46676 31612
rect 46564 30492 46676 30548
rect 46508 30482 46564 30492
rect 46396 30370 46452 30380
rect 46620 30324 46676 30334
rect 46396 30212 46452 30222
rect 46396 30118 46452 30156
rect 46620 29986 46676 30268
rect 46732 30212 46788 31836
rect 46844 32060 47124 32116
rect 46844 31668 46900 32060
rect 47068 31892 47124 31902
rect 47180 31892 47236 32956
rect 47068 31890 47236 31892
rect 47068 31838 47070 31890
rect 47122 31838 47236 31890
rect 47068 31836 47236 31838
rect 47292 32786 47348 32798
rect 47292 32734 47294 32786
rect 47346 32734 47348 32786
rect 47068 31826 47124 31836
rect 46844 31612 47012 31668
rect 46956 31556 47012 31612
rect 46956 31500 47236 31556
rect 46844 31444 46900 31454
rect 46900 31388 47012 31444
rect 46844 31378 46900 31388
rect 46956 31106 47012 31388
rect 46956 31054 46958 31106
rect 47010 31054 47012 31106
rect 46956 31042 47012 31054
rect 46844 30772 46900 30782
rect 46844 30678 46900 30716
rect 46844 30212 46900 30222
rect 46732 30210 46900 30212
rect 46732 30158 46846 30210
rect 46898 30158 46900 30210
rect 46732 30156 46900 30158
rect 46844 30146 46900 30156
rect 47068 30210 47124 30222
rect 47068 30158 47070 30210
rect 47122 30158 47124 30210
rect 46620 29934 46622 29986
rect 46674 29934 46676 29986
rect 46172 29538 46340 29540
rect 46172 29486 46174 29538
rect 46226 29486 46340 29538
rect 46172 29484 46340 29486
rect 46172 29474 46228 29484
rect 45836 29260 46228 29316
rect 45164 28866 45444 28868
rect 45164 28814 45166 28866
rect 45218 28814 45444 28866
rect 45164 28812 45444 28814
rect 45164 28802 45220 28812
rect 45500 28756 45556 28766
rect 45164 28644 45220 28654
rect 45052 28642 45220 28644
rect 45052 28590 45166 28642
rect 45218 28590 45220 28642
rect 45052 28588 45220 28590
rect 45164 28578 45220 28588
rect 45500 28642 45556 28700
rect 45500 28590 45502 28642
rect 45554 28590 45556 28642
rect 45500 28578 45556 28590
rect 46060 28644 46116 28654
rect 46060 28550 46116 28588
rect 45388 28532 45444 28542
rect 45052 27748 45108 27758
rect 44940 27300 44996 27310
rect 44828 27298 44996 27300
rect 44828 27246 44942 27298
rect 44994 27246 44996 27298
rect 44828 27244 44996 27246
rect 44940 27234 44996 27244
rect 44604 26350 44606 26402
rect 44658 26350 44660 26402
rect 44604 26338 44660 26350
rect 44828 26962 44884 26974
rect 44828 26910 44830 26962
rect 44882 26910 44884 26962
rect 44268 26292 44324 26302
rect 44268 25620 44324 26236
rect 44268 25506 44324 25564
rect 44268 25454 44270 25506
rect 44322 25454 44324 25506
rect 44268 25442 44324 25454
rect 43988 25228 44100 25284
rect 43932 25190 43988 25228
rect 44828 25172 44884 26910
rect 44828 25106 44884 25116
rect 43820 25004 44100 25060
rect 43372 24546 43428 24556
rect 43484 24724 43540 24734
rect 43484 23940 43540 24668
rect 43484 23846 43540 23884
rect 43372 23492 43428 23502
rect 43428 23436 43540 23492
rect 43372 23426 43428 23436
rect 43372 23154 43428 23166
rect 43372 23102 43374 23154
rect 43426 23102 43428 23154
rect 43372 22820 43428 23102
rect 43372 22754 43428 22764
rect 43372 22484 43428 22494
rect 43260 22482 43428 22484
rect 43260 22430 43374 22482
rect 43426 22430 43428 22482
rect 43260 22428 43428 22430
rect 43372 22418 43428 22428
rect 43260 22260 43316 22270
rect 43148 22258 43316 22260
rect 43148 22206 43262 22258
rect 43314 22206 43316 22258
rect 43148 22204 43316 22206
rect 43260 22194 43316 22204
rect 43036 21588 43092 21598
rect 43036 20580 43092 21532
rect 43260 21476 43316 21486
rect 43148 21474 43316 21476
rect 43148 21422 43262 21474
rect 43314 21422 43316 21474
rect 43148 21420 43316 21422
rect 43148 20804 43204 21420
rect 43260 21410 43316 21420
rect 43484 20804 43540 23436
rect 43596 23044 43652 23054
rect 43708 23044 43764 24892
rect 43932 24612 43988 24622
rect 43932 23826 43988 24556
rect 43932 23774 43934 23826
rect 43986 23774 43988 23826
rect 43932 23762 43988 23774
rect 43652 22988 43764 23044
rect 43596 22978 43652 22988
rect 43820 22372 43876 22382
rect 44044 22372 44100 25004
rect 45052 24722 45108 27692
rect 45388 27186 45444 28476
rect 46172 28530 46228 29260
rect 46172 28478 46174 28530
rect 46226 28478 46228 28530
rect 46172 28466 46228 28478
rect 45388 27134 45390 27186
rect 45442 27134 45444 27186
rect 45388 27122 45444 27134
rect 45836 27860 45892 27870
rect 45836 27186 45892 27804
rect 45836 27134 45838 27186
rect 45890 27134 45892 27186
rect 45836 27122 45892 27134
rect 46284 27074 46340 29484
rect 46620 28980 46676 29934
rect 46732 29988 46788 29998
rect 46732 29894 46788 29932
rect 46844 29764 46900 29774
rect 46900 29708 47012 29764
rect 46844 29698 46900 29708
rect 46284 27022 46286 27074
rect 46338 27022 46340 27074
rect 45276 26516 45332 26526
rect 45276 25506 45332 26460
rect 46060 26516 46116 26526
rect 46060 26422 46116 26460
rect 45388 26290 45444 26302
rect 45388 26238 45390 26290
rect 45442 26238 45444 26290
rect 45388 26068 45444 26238
rect 45724 26292 45780 26302
rect 45724 26198 45780 26236
rect 46284 26068 46340 27022
rect 45388 26012 46340 26068
rect 45276 25454 45278 25506
rect 45330 25454 45332 25506
rect 45276 25442 45332 25454
rect 45500 25508 45556 25518
rect 45500 25506 45780 25508
rect 45500 25454 45502 25506
rect 45554 25454 45780 25506
rect 45500 25452 45780 25454
rect 45500 25442 45556 25452
rect 45052 24670 45054 24722
rect 45106 24670 45108 24722
rect 45052 24658 45108 24670
rect 45388 25282 45444 25294
rect 45388 25230 45390 25282
rect 45442 25230 45444 25282
rect 44380 24612 44436 24622
rect 44380 24518 44436 24556
rect 44156 23938 44212 23950
rect 44156 23886 44158 23938
rect 44210 23886 44212 23938
rect 44156 23716 44212 23886
rect 44828 23940 44884 23950
rect 44884 23884 44996 23940
rect 44828 23846 44884 23884
rect 44156 23650 44212 23660
rect 44940 23604 44996 23884
rect 44940 23266 44996 23548
rect 44940 23214 44942 23266
rect 44994 23214 44996 23266
rect 44940 23202 44996 23214
rect 44604 22708 44660 22718
rect 43820 22370 44100 22372
rect 43820 22318 43822 22370
rect 43874 22318 44100 22370
rect 43820 22316 44100 22318
rect 44156 22596 44212 22606
rect 44156 22482 44212 22540
rect 44156 22430 44158 22482
rect 44210 22430 44212 22482
rect 43484 20748 43652 20804
rect 43148 20710 43204 20748
rect 43036 20524 43204 20580
rect 42924 19618 42980 19628
rect 43036 20020 43092 20030
rect 42476 19404 42644 19460
rect 42476 19012 42532 19404
rect 42924 19348 42980 19358
rect 42476 18946 42532 18956
rect 42588 19346 42980 19348
rect 42588 19294 42926 19346
rect 42978 19294 42980 19346
rect 42588 19292 42980 19294
rect 42588 18562 42644 19292
rect 42924 19282 42980 19292
rect 43036 19348 43092 19964
rect 43036 19234 43092 19292
rect 43036 19182 43038 19234
rect 43090 19182 43092 19234
rect 42924 19012 42980 19022
rect 42924 18918 42980 18956
rect 43036 18788 43092 19182
rect 42588 18510 42590 18562
rect 42642 18510 42644 18562
rect 42588 18498 42644 18510
rect 42924 18732 43092 18788
rect 42364 18452 42420 18462
rect 42252 18396 42364 18452
rect 42028 18358 42084 18396
rect 42364 18386 42420 18396
rect 42812 18452 42868 18462
rect 42140 18340 42196 18350
rect 42140 18228 42196 18284
rect 42028 18172 42196 18228
rect 42476 18338 42532 18350
rect 42476 18286 42478 18338
rect 42530 18286 42532 18338
rect 41468 16884 41524 16894
rect 41468 16790 41524 16828
rect 41916 16660 41972 16670
rect 42028 16660 42084 18172
rect 42476 18004 42532 18286
rect 42140 17948 42532 18004
rect 42588 18228 42644 18238
rect 42140 16994 42196 17948
rect 42476 17780 42532 17790
rect 42588 17780 42644 18172
rect 42476 17778 42644 17780
rect 42476 17726 42478 17778
rect 42530 17726 42644 17778
rect 42476 17724 42644 17726
rect 42476 17714 42532 17724
rect 42140 16942 42142 16994
rect 42194 16942 42196 16994
rect 42140 16930 42196 16942
rect 41972 16604 42084 16660
rect 41916 16594 41972 16604
rect 40460 9268 40516 9278
rect 40572 9268 40628 15260
rect 40908 16492 41412 16548
rect 40796 14980 40852 14990
rect 40796 14642 40852 14924
rect 40796 14590 40798 14642
rect 40850 14590 40852 14642
rect 40796 14578 40852 14590
rect 40908 10164 40964 16492
rect 42364 16212 42420 16222
rect 41916 16210 42420 16212
rect 41916 16158 42366 16210
rect 42418 16158 42420 16210
rect 41916 16156 42420 16158
rect 41468 15540 41524 15550
rect 41916 15540 41972 16156
rect 42364 16146 42420 16156
rect 42700 16100 42756 16110
rect 41468 15538 41972 15540
rect 41468 15486 41470 15538
rect 41522 15486 41972 15538
rect 41468 15484 41972 15486
rect 41468 15474 41524 15484
rect 41132 15428 41188 15438
rect 41188 15372 41300 15428
rect 41132 15334 41188 15372
rect 41020 13972 41076 13982
rect 41020 13878 41076 13916
rect 41244 13972 41300 15372
rect 41916 15426 41972 15484
rect 41916 15374 41918 15426
rect 41970 15374 41972 15426
rect 41692 15092 41748 15102
rect 41356 14644 41412 14654
rect 41356 14550 41412 14588
rect 41244 13878 41300 13916
rect 41468 13972 41524 13982
rect 41692 13972 41748 15036
rect 41916 14980 41972 15374
rect 42476 16098 42756 16100
rect 42476 16046 42702 16098
rect 42754 16046 42756 16098
rect 42476 16044 42756 16046
rect 42028 15314 42084 15326
rect 42028 15262 42030 15314
rect 42082 15262 42084 15314
rect 42028 15148 42084 15262
rect 42140 15316 42196 15326
rect 42140 15314 42308 15316
rect 42140 15262 42142 15314
rect 42194 15262 42308 15314
rect 42140 15260 42308 15262
rect 42140 15250 42196 15260
rect 42028 15082 42084 15092
rect 41916 14924 42084 14980
rect 41468 13970 41748 13972
rect 41468 13918 41470 13970
rect 41522 13918 41748 13970
rect 41468 13916 41748 13918
rect 41468 13860 41524 13916
rect 41468 13794 41524 13804
rect 41356 13748 41412 13758
rect 41356 13654 41412 13692
rect 41692 13746 41748 13916
rect 42028 13860 42084 14924
rect 42252 14644 42308 15260
rect 42028 13794 42084 13804
rect 42140 13972 42196 13982
rect 41692 13694 41694 13746
rect 41746 13694 41748 13746
rect 41692 13682 41748 13694
rect 42140 13746 42196 13916
rect 42140 13694 42142 13746
rect 42194 13694 42196 13746
rect 42140 13682 42196 13694
rect 42252 13746 42308 14588
rect 42252 13694 42254 13746
rect 42306 13694 42308 13746
rect 41916 13634 41972 13646
rect 41916 13582 41918 13634
rect 41970 13582 41972 13634
rect 41804 13524 41860 13534
rect 41580 13300 41636 13310
rect 41580 13074 41636 13244
rect 41580 13022 41582 13074
rect 41634 13022 41636 13074
rect 41580 13010 41636 13022
rect 41244 12628 41300 12638
rect 41244 12180 41300 12572
rect 41244 12086 41300 12124
rect 41468 12180 41524 12190
rect 41468 12086 41524 12124
rect 41692 12178 41748 12190
rect 41692 12126 41694 12178
rect 41746 12126 41748 12178
rect 41020 12068 41076 12078
rect 41020 11974 41076 12012
rect 41692 11844 41748 12126
rect 41692 11778 41748 11788
rect 41244 10724 41300 10734
rect 41244 10630 41300 10668
rect 41468 10388 41524 10398
rect 41468 10294 41524 10332
rect 41692 10386 41748 10398
rect 41692 10334 41694 10386
rect 41746 10334 41748 10386
rect 41244 10276 41300 10286
rect 41244 10164 41300 10220
rect 40908 10108 41300 10164
rect 41132 9940 41188 9950
rect 41132 9846 41188 9884
rect 40460 9266 40628 9268
rect 40460 9214 40462 9266
rect 40514 9214 40628 9266
rect 40460 9212 40628 9214
rect 41244 9266 41300 10108
rect 41692 9940 41748 10334
rect 41804 10164 41860 13468
rect 41916 12740 41972 13582
rect 42252 13524 42308 13694
rect 42476 13636 42532 16044
rect 42700 16034 42756 16044
rect 42812 15874 42868 18396
rect 42924 17778 42980 18732
rect 42924 17726 42926 17778
rect 42978 17726 42980 17778
rect 42924 17714 42980 17726
rect 43036 18564 43092 18574
rect 42924 15988 42980 15998
rect 42924 15894 42980 15932
rect 42812 15822 42814 15874
rect 42866 15822 42868 15874
rect 42812 15810 42868 15822
rect 43036 15314 43092 18508
rect 43036 15262 43038 15314
rect 43090 15262 43092 15314
rect 43036 15148 43092 15262
rect 42588 15090 42644 15102
rect 42588 15038 42590 15090
rect 42642 15038 42644 15090
rect 42588 13748 42644 15038
rect 42924 15092 43092 15148
rect 42812 13972 42868 13982
rect 42812 13878 42868 13916
rect 42588 13692 42868 13748
rect 42028 13468 42308 13524
rect 42364 13580 42532 13636
rect 42588 13580 42756 13636
rect 42028 13074 42084 13468
rect 42364 13412 42420 13580
rect 42588 13524 42644 13580
rect 42588 13458 42644 13468
rect 42700 13522 42756 13580
rect 42700 13470 42702 13522
rect 42754 13470 42756 13522
rect 42700 13458 42756 13470
rect 42812 13524 42868 13692
rect 42812 13458 42868 13468
rect 42028 13022 42030 13074
rect 42082 13022 42084 13074
rect 42028 13010 42084 13022
rect 42140 13356 42420 13412
rect 41916 12674 41972 12684
rect 42028 12852 42084 12862
rect 41916 12178 41972 12190
rect 41916 12126 41918 12178
rect 41970 12126 41972 12178
rect 41916 10610 41972 12126
rect 41916 10558 41918 10610
rect 41970 10558 41972 10610
rect 41916 10500 41972 10558
rect 41916 10434 41972 10444
rect 41804 10098 41860 10108
rect 42028 10052 42084 12796
rect 42140 11732 42196 13356
rect 42700 13300 42756 13310
rect 42756 13244 42868 13300
rect 42700 13234 42756 13244
rect 42364 13076 42420 13086
rect 42364 12962 42420 13020
rect 42364 12910 42366 12962
rect 42418 12910 42420 12962
rect 42364 12898 42420 12910
rect 42812 12962 42868 13244
rect 42812 12910 42814 12962
rect 42866 12910 42868 12962
rect 42812 12898 42868 12910
rect 42476 12740 42532 12750
rect 42476 12178 42532 12684
rect 42588 12404 42644 12414
rect 42812 12404 42868 12414
rect 42644 12348 42756 12404
rect 42588 12338 42644 12348
rect 42476 12126 42478 12178
rect 42530 12126 42532 12178
rect 42476 12114 42532 12126
rect 42700 12292 42756 12348
rect 42700 12178 42756 12236
rect 42812 12290 42868 12348
rect 42812 12238 42814 12290
rect 42866 12238 42868 12290
rect 42812 12226 42868 12238
rect 42700 12126 42702 12178
rect 42754 12126 42756 12178
rect 42700 12114 42756 12126
rect 42924 12068 42980 15092
rect 42364 11956 42420 11966
rect 42476 11956 42532 11966
rect 42364 11954 42476 11956
rect 42364 11902 42366 11954
rect 42418 11902 42476 11954
rect 42364 11900 42476 11902
rect 42364 11890 42420 11900
rect 42140 11676 42420 11732
rect 42364 10834 42420 11676
rect 42364 10782 42366 10834
rect 42418 10782 42420 10834
rect 42364 10770 42420 10782
rect 42476 10612 42532 11900
rect 42924 11396 42980 12012
rect 43036 13522 43092 13534
rect 43036 13470 43038 13522
rect 43090 13470 43092 13522
rect 43036 11508 43092 13470
rect 43148 13074 43204 20524
rect 43260 20578 43316 20590
rect 43260 20526 43262 20578
rect 43314 20526 43316 20578
rect 43260 20468 43316 20526
rect 43372 20580 43428 20590
rect 43372 20486 43428 20524
rect 43484 20578 43540 20590
rect 43484 20526 43486 20578
rect 43538 20526 43540 20578
rect 43260 20402 43316 20412
rect 43260 19908 43316 19918
rect 43484 19908 43540 20526
rect 43596 20020 43652 20748
rect 43596 19954 43652 19964
rect 43708 20690 43764 20702
rect 43708 20638 43710 20690
rect 43762 20638 43764 20690
rect 43316 19852 43540 19908
rect 43260 19234 43316 19852
rect 43708 19572 43764 20638
rect 43260 19182 43262 19234
rect 43314 19182 43316 19234
rect 43260 19170 43316 19182
rect 43596 19516 43764 19572
rect 43596 19236 43652 19516
rect 43484 19122 43540 19134
rect 43484 19070 43486 19122
rect 43538 19070 43540 19122
rect 43484 18564 43540 19070
rect 43484 18498 43540 18508
rect 43260 18340 43316 18350
rect 43596 18340 43652 19180
rect 43260 18338 43652 18340
rect 43260 18286 43262 18338
rect 43314 18286 43652 18338
rect 43260 18284 43652 18286
rect 43260 18274 43316 18284
rect 43372 18004 43428 18014
rect 43372 17778 43428 17948
rect 43372 17726 43374 17778
rect 43426 17726 43428 17778
rect 43372 17714 43428 17726
rect 43820 17778 43876 22316
rect 44156 22260 44212 22430
rect 43932 22204 44212 22260
rect 43932 18900 43988 22204
rect 44044 20692 44100 20702
rect 44044 20598 44100 20636
rect 44156 20580 44212 20590
rect 44156 20578 44436 20580
rect 44156 20526 44158 20578
rect 44210 20526 44436 20578
rect 44156 20524 44436 20526
rect 44156 20514 44212 20524
rect 44380 20130 44436 20524
rect 44380 20078 44382 20130
rect 44434 20078 44436 20130
rect 44380 20066 44436 20078
rect 44044 19908 44100 19918
rect 44044 19234 44100 19852
rect 44044 19182 44046 19234
rect 44098 19182 44100 19234
rect 44044 19170 44100 19182
rect 44268 19572 44324 19582
rect 44268 19124 44324 19516
rect 43932 18834 43988 18844
rect 44156 19010 44212 19022
rect 44156 18958 44158 19010
rect 44210 18958 44212 19010
rect 44156 18900 44212 18958
rect 44156 18834 44212 18844
rect 44268 18676 44324 19068
rect 44380 19012 44436 19022
rect 44380 19010 44548 19012
rect 44380 18958 44382 19010
rect 44434 18958 44548 19010
rect 44380 18956 44548 18958
rect 44380 18946 44436 18956
rect 43820 17726 43822 17778
rect 43874 17726 43876 17778
rect 43820 17714 43876 17726
rect 44156 18620 44324 18676
rect 44156 17666 44212 18620
rect 44268 18452 44324 18462
rect 44324 18396 44436 18452
rect 44268 18386 44324 18396
rect 44156 17614 44158 17666
rect 44210 17614 44212 17666
rect 44156 17602 44212 17614
rect 44156 17444 44212 17454
rect 44156 16212 44212 17388
rect 44268 16772 44324 16782
rect 44380 16772 44436 18396
rect 44268 16770 44436 16772
rect 44268 16718 44270 16770
rect 44322 16718 44436 16770
rect 44268 16716 44436 16718
rect 44268 16706 44324 16716
rect 44492 16548 44548 18956
rect 44604 16660 44660 22652
rect 45388 22596 45444 25230
rect 45612 25282 45668 25294
rect 45612 25230 45614 25282
rect 45666 25230 45668 25282
rect 45612 24836 45668 25230
rect 45724 25060 45780 25452
rect 46284 25506 46340 26012
rect 46284 25454 46286 25506
rect 46338 25454 46340 25506
rect 46284 25442 46340 25454
rect 46396 28924 46676 28980
rect 45836 25394 45892 25406
rect 45836 25342 45838 25394
rect 45890 25342 45892 25394
rect 45836 25284 45892 25342
rect 45836 25218 45892 25228
rect 46396 25284 46452 28924
rect 46508 28754 46564 28766
rect 46508 28702 46510 28754
rect 46562 28702 46564 28754
rect 46508 27972 46564 28702
rect 46956 28530 47012 29708
rect 47068 29540 47124 30158
rect 47068 29474 47124 29484
rect 47068 28756 47124 28766
rect 47180 28756 47236 31500
rect 47292 30996 47348 32734
rect 47404 32562 47460 32574
rect 47404 32510 47406 32562
rect 47458 32510 47460 32562
rect 47404 31220 47460 32510
rect 47516 31780 47572 35420
rect 47628 35410 47684 35420
rect 47964 35476 48020 35486
rect 47964 35474 48132 35476
rect 47964 35422 47966 35474
rect 48018 35422 48132 35474
rect 47964 35420 48132 35422
rect 47964 35410 48020 35420
rect 47628 34916 47684 34926
rect 47628 34822 47684 34860
rect 47740 34692 47796 34702
rect 47628 34020 47684 34030
rect 47628 33926 47684 33964
rect 47628 32564 47684 32574
rect 47628 32470 47684 32508
rect 47740 31892 47796 34636
rect 48076 32900 48132 35420
rect 48188 35028 48244 35038
rect 48188 34934 48244 34972
rect 48188 34692 48244 34702
rect 48188 34354 48244 34636
rect 48188 34302 48190 34354
rect 48242 34302 48244 34354
rect 48188 34290 48244 34302
rect 48076 32834 48132 32844
rect 48076 32676 48132 32686
rect 48076 32582 48132 32620
rect 47964 32562 48020 32574
rect 47964 32510 47966 32562
rect 48018 32510 48020 32562
rect 47852 32452 47908 32462
rect 47964 32452 48020 32510
rect 47908 32396 48020 32452
rect 48076 32452 48132 32462
rect 47852 32386 47908 32396
rect 48076 32338 48132 32396
rect 48076 32286 48078 32338
rect 48130 32286 48132 32338
rect 48076 32274 48132 32286
rect 47740 31826 47796 31836
rect 48300 31892 48356 35532
rect 48412 34916 48468 36428
rect 48748 35924 48804 35934
rect 48748 35830 48804 35868
rect 48972 35028 49028 39004
rect 49084 38834 49140 38846
rect 49084 38782 49086 38834
rect 49138 38782 49140 38834
rect 49084 37492 49140 38782
rect 49196 38724 49252 39676
rect 49196 38162 49252 38668
rect 49196 38110 49198 38162
rect 49250 38110 49252 38162
rect 49196 38098 49252 38110
rect 49084 37436 49252 37492
rect 49084 37268 49140 37278
rect 49084 37174 49140 37212
rect 49084 37044 49140 37054
rect 49084 36372 49140 36988
rect 49196 36596 49252 37436
rect 49196 36502 49252 36540
rect 49084 36316 49252 36372
rect 49084 36148 49140 36158
rect 49084 35922 49140 36092
rect 49084 35870 49086 35922
rect 49138 35870 49140 35922
rect 49084 35858 49140 35870
rect 49084 35028 49140 35038
rect 48972 35026 49140 35028
rect 48972 34974 49086 35026
rect 49138 34974 49140 35026
rect 48972 34972 49140 34974
rect 49084 34962 49140 34972
rect 48412 34914 48692 34916
rect 48412 34862 48414 34914
rect 48466 34862 48692 34914
rect 48412 34860 48692 34862
rect 48412 34850 48468 34860
rect 48412 34244 48468 34254
rect 48468 34188 48580 34244
rect 48412 34178 48468 34188
rect 48300 31826 48356 31836
rect 48412 32564 48468 32574
rect 47516 31714 47572 31724
rect 48412 31668 48468 32508
rect 48524 32452 48580 34188
rect 48524 32386 48580 32396
rect 48300 31612 48468 31668
rect 47404 31164 47908 31220
rect 47292 30930 47348 30940
rect 47628 30996 47684 31006
rect 47628 30902 47684 30940
rect 47740 30994 47796 31006
rect 47740 30942 47742 30994
rect 47794 30942 47796 30994
rect 47404 30436 47460 30446
rect 47068 28754 47236 28756
rect 47068 28702 47070 28754
rect 47122 28702 47236 28754
rect 47068 28700 47236 28702
rect 47292 30380 47404 30436
rect 47068 28690 47124 28700
rect 46956 28478 46958 28530
rect 47010 28478 47012 28530
rect 46956 28466 47012 28478
rect 47180 28532 47236 28542
rect 47292 28532 47348 30380
rect 47404 30342 47460 30380
rect 47516 30324 47572 30334
rect 47740 30324 47796 30942
rect 47572 30268 47684 30324
rect 47516 30258 47572 30268
rect 47404 30212 47460 30250
rect 47404 30146 47460 30156
rect 47628 30100 47684 30268
rect 47740 30258 47796 30268
rect 47852 30882 47908 31164
rect 47852 30830 47854 30882
rect 47906 30830 47908 30882
rect 47740 30100 47796 30110
rect 47628 30098 47796 30100
rect 47628 30046 47742 30098
rect 47794 30046 47796 30098
rect 47628 30044 47796 30046
rect 47740 30034 47796 30044
rect 47180 28530 47348 28532
rect 47180 28478 47182 28530
rect 47234 28478 47348 28530
rect 47180 28476 47348 28478
rect 47404 29988 47460 29998
rect 47404 28644 47460 29932
rect 47740 28868 47796 28878
rect 47740 28774 47796 28812
rect 47404 28530 47460 28588
rect 47404 28478 47406 28530
rect 47458 28478 47460 28530
rect 47180 28466 47236 28476
rect 47404 28466 47460 28478
rect 47852 28530 47908 30830
rect 47964 30994 48020 31006
rect 47964 30942 47966 30994
rect 48018 30942 48020 30994
rect 47964 30436 48020 30942
rect 48076 30994 48132 31006
rect 48076 30942 48078 30994
rect 48130 30942 48132 30994
rect 48076 30660 48132 30942
rect 48076 30594 48132 30604
rect 47964 30370 48020 30380
rect 48300 30322 48356 31612
rect 48636 31220 48692 34860
rect 48748 34804 48804 34814
rect 48748 34580 48804 34748
rect 48748 34524 48916 34580
rect 48748 34356 48804 34366
rect 48748 34242 48804 34300
rect 48860 34354 48916 34524
rect 48860 34302 48862 34354
rect 48914 34302 48916 34354
rect 48860 34290 48916 34302
rect 48748 34190 48750 34242
rect 48802 34190 48804 34242
rect 48748 34178 48804 34190
rect 49084 34132 49140 34142
rect 49196 34132 49252 36316
rect 49308 36148 49364 41916
rect 49420 41300 49476 44268
rect 49420 41234 49476 41244
rect 49308 36082 49364 36092
rect 49420 40852 49476 40862
rect 49084 34130 49252 34132
rect 49084 34078 49086 34130
rect 49138 34078 49252 34130
rect 49084 34076 49252 34078
rect 49084 34066 49140 34076
rect 48860 34020 48916 34030
rect 48916 33964 49028 34020
rect 48860 33954 48916 33964
rect 48748 32676 48804 32686
rect 48748 32582 48804 32620
rect 48748 31220 48804 31230
rect 48300 30270 48302 30322
rect 48354 30270 48356 30322
rect 48300 30258 48356 30270
rect 48412 31218 48804 31220
rect 48412 31166 48750 31218
rect 48802 31166 48804 31218
rect 48412 31164 48804 31166
rect 48188 30212 48244 30222
rect 48076 28644 48132 28654
rect 48076 28550 48132 28588
rect 47852 28478 47854 28530
rect 47906 28478 47908 28530
rect 47852 28466 47908 28478
rect 48076 28084 48132 28094
rect 48188 28084 48244 30156
rect 48412 30210 48468 31164
rect 48748 31154 48804 31164
rect 48412 30158 48414 30210
rect 48466 30158 48468 30210
rect 48412 30146 48468 30158
rect 48524 30660 48580 30670
rect 48524 30210 48580 30604
rect 48524 30158 48526 30210
rect 48578 30158 48580 30210
rect 48524 29652 48580 30158
rect 48076 28082 48244 28084
rect 48076 28030 48078 28082
rect 48130 28030 48244 28082
rect 48076 28028 48244 28030
rect 48300 29596 48580 29652
rect 48636 30548 48692 30558
rect 48076 28018 48132 28028
rect 46508 27916 46900 27972
rect 46844 27858 46900 27916
rect 46844 27806 46846 27858
rect 46898 27806 46900 27858
rect 46620 27748 46676 27758
rect 46508 27636 46564 27646
rect 46508 27542 46564 27580
rect 46508 26516 46564 26526
rect 46508 26422 46564 26460
rect 46620 26404 46676 27692
rect 46844 26908 46900 27806
rect 47068 27748 47124 27758
rect 47068 27746 47348 27748
rect 47068 27694 47070 27746
rect 47122 27694 47348 27746
rect 47068 27692 47348 27694
rect 47068 27682 47124 27692
rect 47068 26964 47124 26974
rect 46844 26852 47012 26908
rect 47068 26870 47124 26908
rect 46620 26310 46676 26348
rect 46844 26404 46900 26414
rect 46844 26310 46900 26348
rect 46732 26180 46788 26190
rect 46732 26086 46788 26124
rect 46956 26068 47012 26852
rect 47068 26292 47124 26302
rect 47068 26198 47124 26236
rect 46396 25218 46452 25228
rect 46844 26012 47012 26068
rect 45724 25004 46788 25060
rect 45836 24836 45892 24846
rect 45612 24834 45892 24836
rect 45612 24782 45838 24834
rect 45890 24782 45892 24834
rect 45612 24780 45892 24782
rect 45500 24722 45556 24734
rect 45500 24670 45502 24722
rect 45554 24670 45556 24722
rect 45500 23716 45556 24670
rect 45836 24724 45892 24780
rect 46284 24836 46340 24846
rect 46284 24742 46340 24780
rect 46732 24834 46788 25004
rect 46732 24782 46734 24834
rect 46786 24782 46788 24834
rect 46732 24770 46788 24782
rect 45836 24658 45892 24668
rect 46172 24612 46228 24622
rect 46172 24518 46228 24556
rect 46620 24500 46676 24510
rect 46396 24498 46676 24500
rect 46396 24446 46622 24498
rect 46674 24446 46676 24498
rect 46396 24444 46676 24446
rect 46396 24164 46452 24444
rect 46620 24434 46676 24444
rect 45612 24108 46452 24164
rect 45612 24050 45668 24108
rect 45612 23998 45614 24050
rect 45666 23998 45668 24050
rect 45612 23986 45668 23998
rect 45500 23650 45556 23660
rect 46060 23492 46116 23502
rect 46116 23436 46340 23492
rect 46060 23426 46116 23436
rect 45388 22530 45444 22540
rect 44940 22484 44996 22494
rect 44940 22390 44996 22428
rect 45164 22372 45220 22382
rect 45948 22372 46004 22382
rect 46284 22372 46340 23436
rect 46844 23156 46900 26012
rect 46956 25732 47012 25742
rect 46956 25618 47012 25676
rect 46956 25566 46958 25618
rect 47010 25566 47012 25618
rect 46956 25554 47012 25566
rect 47180 24948 47236 24958
rect 47180 24854 47236 24892
rect 47068 24500 47124 24510
rect 46844 23100 47012 23156
rect 45164 22370 45332 22372
rect 45164 22318 45166 22370
rect 45218 22318 45332 22370
rect 45164 22316 45332 22318
rect 45164 22306 45220 22316
rect 45276 21476 45332 22316
rect 45948 22278 46004 22316
rect 46060 22370 46340 22372
rect 46060 22318 46286 22370
rect 46338 22318 46340 22370
rect 46060 22316 46340 22318
rect 45500 22148 45556 22158
rect 45500 21588 45556 22092
rect 46060 21924 46116 22316
rect 46284 22306 46340 22316
rect 45948 21868 46116 21924
rect 45836 21588 45892 21598
rect 45500 21586 45892 21588
rect 45500 21534 45838 21586
rect 45890 21534 45892 21586
rect 45500 21532 45892 21534
rect 45388 21476 45444 21486
rect 45276 21474 45444 21476
rect 45276 21422 45390 21474
rect 45442 21422 45444 21474
rect 45276 21420 45444 21422
rect 45388 21410 45444 21420
rect 45836 21140 45892 21532
rect 45948 21476 46004 21868
rect 46844 21812 46900 21822
rect 46844 21718 46900 21756
rect 46956 21812 47012 23100
rect 47068 22482 47124 24444
rect 47068 22430 47070 22482
rect 47122 22430 47124 22482
rect 47068 22418 47124 22430
rect 47292 22148 47348 27692
rect 47628 27746 47684 27758
rect 47628 27694 47630 27746
rect 47682 27694 47684 27746
rect 47516 27634 47572 27646
rect 47516 27582 47518 27634
rect 47570 27582 47572 27634
rect 47516 26964 47572 27582
rect 47516 26898 47572 26908
rect 47628 26908 47684 27694
rect 48188 27746 48244 27758
rect 48188 27694 48190 27746
rect 48242 27694 48244 27746
rect 48076 27188 48132 27198
rect 47628 26852 47796 26908
rect 47628 26628 47684 26638
rect 47516 26516 47572 26526
rect 47516 26290 47572 26460
rect 47628 26514 47684 26572
rect 47628 26462 47630 26514
rect 47682 26462 47684 26514
rect 47628 26450 47684 26462
rect 47740 26514 47796 26852
rect 47740 26462 47742 26514
rect 47794 26462 47796 26514
rect 47740 26450 47796 26462
rect 47516 26238 47518 26290
rect 47570 26238 47572 26290
rect 47516 25396 47572 26238
rect 47516 25330 47572 25340
rect 47852 26404 47908 26414
rect 47852 26290 47908 26348
rect 48076 26402 48132 27132
rect 48076 26350 48078 26402
rect 48130 26350 48132 26402
rect 48076 26338 48132 26350
rect 47852 26238 47854 26290
rect 47906 26238 47908 26290
rect 47740 25172 47796 25182
rect 47628 24610 47684 24622
rect 47628 24558 47630 24610
rect 47682 24558 47684 24610
rect 47628 24388 47684 24558
rect 47628 24322 47684 24332
rect 47740 24050 47796 25116
rect 47740 23998 47742 24050
rect 47794 23998 47796 24050
rect 47740 23986 47796 23998
rect 47852 24724 47908 26238
rect 48188 26292 48244 27694
rect 48300 27636 48356 29596
rect 48412 28644 48468 28654
rect 48636 28644 48692 30492
rect 48860 30436 48916 30446
rect 48860 30342 48916 30380
rect 48748 30324 48804 30334
rect 48748 29650 48804 30268
rect 48748 29598 48750 29650
rect 48802 29598 48804 29650
rect 48748 29586 48804 29598
rect 48860 29540 48916 29550
rect 48860 29446 48916 29484
rect 48412 28642 48692 28644
rect 48412 28590 48414 28642
rect 48466 28590 48692 28642
rect 48412 28588 48692 28590
rect 48748 28754 48804 28766
rect 48748 28702 48750 28754
rect 48802 28702 48804 28754
rect 48412 28578 48468 28588
rect 48748 27860 48804 28702
rect 48636 27804 48804 27860
rect 48412 27636 48468 27646
rect 48300 27580 48412 27636
rect 48412 27570 48468 27580
rect 48636 27412 48692 27804
rect 48860 27746 48916 27758
rect 48860 27694 48862 27746
rect 48914 27694 48916 27746
rect 48748 27636 48804 27646
rect 48748 27542 48804 27580
rect 48636 27356 48804 27412
rect 48748 26628 48804 27356
rect 48860 27188 48916 27694
rect 48972 27748 49028 33964
rect 49196 33460 49252 33470
rect 49196 33458 49364 33460
rect 49196 33406 49198 33458
rect 49250 33406 49364 33458
rect 49196 33404 49364 33406
rect 49196 33394 49252 33404
rect 49084 32562 49140 32574
rect 49084 32510 49086 32562
rect 49138 32510 49140 32562
rect 49084 32340 49140 32510
rect 49084 32274 49140 32284
rect 49196 31892 49252 31902
rect 49084 31836 49196 31892
rect 49084 31218 49140 31836
rect 49196 31798 49252 31836
rect 49084 31166 49086 31218
rect 49138 31166 49140 31218
rect 49084 31154 49140 31166
rect 49308 30996 49364 33404
rect 49308 30930 49364 30940
rect 49084 30100 49140 30110
rect 49140 30044 49252 30100
rect 49084 30034 49140 30044
rect 48972 27682 49028 27692
rect 49084 29540 49140 29550
rect 48860 27122 48916 27132
rect 49084 26908 49140 29484
rect 49196 28642 49252 30044
rect 49196 28590 49198 28642
rect 49250 28590 49252 28642
rect 49196 27636 49252 28590
rect 49196 27570 49252 27580
rect 49196 27188 49252 27198
rect 49196 27094 49252 27132
rect 49420 26908 49476 40796
rect 49532 39620 49588 44492
rect 49644 40068 49700 46844
rect 49644 40002 49700 40012
rect 49532 39554 49588 39564
rect 49532 36596 49588 36606
rect 49532 30436 49588 36540
rect 49532 30370 49588 30380
rect 48748 26562 48804 26572
rect 48972 26852 49140 26908
rect 49308 26852 49476 26908
rect 48188 25620 48244 26236
rect 48860 26180 48916 26190
rect 48860 26086 48916 26124
rect 48748 26066 48804 26078
rect 48748 26014 48750 26066
rect 48802 26014 48804 26066
rect 48748 25732 48804 26014
rect 48748 25666 48804 25676
rect 48188 25554 48244 25564
rect 48188 25396 48244 25406
rect 47852 23828 47908 24668
rect 47852 23762 47908 23772
rect 48076 24724 48132 24734
rect 48076 23380 48132 24668
rect 48188 23938 48244 25340
rect 48860 24610 48916 24622
rect 48860 24558 48862 24610
rect 48914 24558 48916 24610
rect 48748 24500 48804 24510
rect 48748 24406 48804 24444
rect 48188 23886 48190 23938
rect 48242 23886 48244 23938
rect 48188 23874 48244 23886
rect 48300 24388 48356 24398
rect 48300 23938 48356 24332
rect 48412 24052 48468 24062
rect 48860 24052 48916 24558
rect 48412 24050 48916 24052
rect 48412 23998 48414 24050
rect 48466 23998 48916 24050
rect 48412 23996 48916 23998
rect 48412 23986 48468 23996
rect 48300 23886 48302 23938
rect 48354 23886 48356 23938
rect 48300 23874 48356 23886
rect 48524 23828 48580 23838
rect 48524 23734 48580 23772
rect 48748 23828 48804 23838
rect 48972 23828 49028 26852
rect 49084 25620 49140 25630
rect 49084 25526 49140 25564
rect 49196 24052 49252 24062
rect 49196 23958 49252 23996
rect 48748 23826 49028 23828
rect 48748 23774 48750 23826
rect 48802 23774 49028 23826
rect 48748 23772 49028 23774
rect 48748 23762 48804 23772
rect 48076 23314 48132 23324
rect 48972 23156 49028 23772
rect 49308 23548 49364 26852
rect 49308 23492 49476 23548
rect 48972 23100 49252 23156
rect 48860 23044 48916 23054
rect 48860 23042 49140 23044
rect 48860 22990 48862 23042
rect 48914 22990 49140 23042
rect 48860 22988 49140 22990
rect 48860 22978 48916 22988
rect 47292 22082 47348 22092
rect 48748 22930 48804 22942
rect 48748 22878 48750 22930
rect 48802 22878 48804 22930
rect 48748 21924 48804 22878
rect 49084 21924 49140 22988
rect 49196 22482 49252 23100
rect 49196 22430 49198 22482
rect 49250 22430 49252 22482
rect 49196 22418 49252 22430
rect 48748 21868 49028 21924
rect 49084 21868 49252 21924
rect 47292 21812 47348 21822
rect 46956 21810 47348 21812
rect 46956 21758 47294 21810
rect 47346 21758 47348 21810
rect 46956 21756 47348 21758
rect 46060 21698 46116 21710
rect 46060 21646 46062 21698
rect 46114 21646 46116 21698
rect 46060 21588 46116 21646
rect 46956 21698 47012 21756
rect 47292 21746 47348 21756
rect 47740 21812 47796 21822
rect 47740 21718 47796 21756
rect 46956 21646 46958 21698
rect 47010 21646 47012 21698
rect 46956 21634 47012 21646
rect 46396 21588 46452 21598
rect 46060 21586 46452 21588
rect 46060 21534 46398 21586
rect 46450 21534 46452 21586
rect 46060 21532 46452 21534
rect 45948 21420 46340 21476
rect 45836 21084 46116 21140
rect 45724 20804 45780 20814
rect 45724 20710 45780 20748
rect 44940 20690 44996 20702
rect 45948 20692 46004 20702
rect 44940 20638 44942 20690
rect 44994 20638 44996 20690
rect 44828 20580 44884 20590
rect 44828 17778 44884 20524
rect 44940 20132 44996 20638
rect 45836 20690 46004 20692
rect 45836 20638 45950 20690
rect 46002 20638 46004 20690
rect 45836 20636 46004 20638
rect 44940 20066 44996 20076
rect 45052 20578 45108 20590
rect 45052 20526 45054 20578
rect 45106 20526 45108 20578
rect 45052 20020 45108 20526
rect 45388 20578 45444 20590
rect 45388 20526 45390 20578
rect 45442 20526 45444 20578
rect 45052 19954 45108 19964
rect 45164 20132 45220 20142
rect 45164 20018 45220 20076
rect 45164 19966 45166 20018
rect 45218 19966 45220 20018
rect 45164 19954 45220 19966
rect 45052 19796 45108 19806
rect 45052 19346 45108 19740
rect 45052 19294 45054 19346
rect 45106 19294 45108 19346
rect 45052 19282 45108 19294
rect 45388 19012 45444 20526
rect 45500 20018 45556 20030
rect 45500 19966 45502 20018
rect 45554 19966 45556 20018
rect 45500 19236 45556 19966
rect 45724 20020 45780 20030
rect 45724 19926 45780 19964
rect 45612 19908 45668 19918
rect 45612 19814 45668 19852
rect 45500 19142 45556 19180
rect 45388 18956 45556 19012
rect 45388 18340 45444 18350
rect 44940 18338 45444 18340
rect 44940 18286 45390 18338
rect 45442 18286 45444 18338
rect 44940 18284 45444 18286
rect 44940 17890 44996 18284
rect 45388 18274 45444 18284
rect 44940 17838 44942 17890
rect 44994 17838 44996 17890
rect 44940 17826 44996 17838
rect 44828 17726 44830 17778
rect 44882 17726 44884 17778
rect 44828 17714 44884 17726
rect 44604 16594 44660 16604
rect 44716 17668 44772 17678
rect 44716 16884 44772 17612
rect 45500 17666 45556 18956
rect 45500 17614 45502 17666
rect 45554 17614 45556 17666
rect 45500 17602 45556 17614
rect 45724 18340 45780 18350
rect 45724 17666 45780 18284
rect 45724 17614 45726 17666
rect 45778 17614 45780 17666
rect 45724 17602 45780 17614
rect 45836 17668 45892 20636
rect 45948 20626 46004 20636
rect 46060 19908 46116 21084
rect 46284 20802 46340 21420
rect 46284 20750 46286 20802
rect 46338 20750 46340 20802
rect 46284 20132 46340 20750
rect 45948 19122 46004 19134
rect 45948 19070 45950 19122
rect 46002 19070 46004 19122
rect 45948 18564 46004 19070
rect 45948 18498 46004 18508
rect 45836 17612 46004 17668
rect 45276 17556 45332 17566
rect 44492 16482 44548 16492
rect 44268 16212 44324 16222
rect 44156 16210 44324 16212
rect 44156 16158 44270 16210
rect 44322 16158 44324 16210
rect 44156 16156 44324 16158
rect 44268 16146 44324 16156
rect 43596 15986 43652 15998
rect 43596 15934 43598 15986
rect 43650 15934 43652 15986
rect 43484 14420 43540 14430
rect 43148 13022 43150 13074
rect 43202 13022 43204 13074
rect 43148 13010 43204 13022
rect 43372 14418 43540 14420
rect 43372 14366 43486 14418
rect 43538 14366 43540 14418
rect 43372 14364 43540 14366
rect 43372 12404 43428 14364
rect 43484 14354 43540 14364
rect 43484 13746 43540 13758
rect 43484 13694 43486 13746
rect 43538 13694 43540 13746
rect 43484 13636 43540 13694
rect 43484 13570 43540 13580
rect 43596 12852 43652 15934
rect 43820 15988 43876 15998
rect 43596 12786 43652 12796
rect 43708 13412 43764 13422
rect 43372 12338 43428 12348
rect 43260 12292 43316 12302
rect 43260 12178 43316 12236
rect 43260 12126 43262 12178
rect 43314 12126 43316 12178
rect 43260 12114 43316 12126
rect 43484 12180 43540 12190
rect 43484 12086 43540 12124
rect 43148 11954 43204 11966
rect 43148 11902 43150 11954
rect 43202 11902 43204 11954
rect 43148 11732 43204 11902
rect 43596 11954 43652 11966
rect 43596 11902 43598 11954
rect 43650 11902 43652 11954
rect 43148 11666 43204 11676
rect 43484 11844 43540 11854
rect 43036 11452 43316 11508
rect 42924 11394 43092 11396
rect 42924 11342 42926 11394
rect 42978 11342 43092 11394
rect 42924 11340 43092 11342
rect 42924 11330 42980 11340
rect 42028 9986 42084 9996
rect 42252 10556 42532 10612
rect 42924 10724 42980 10734
rect 41748 9884 41860 9940
rect 41692 9874 41748 9884
rect 41468 9826 41524 9838
rect 41468 9774 41470 9826
rect 41522 9774 41524 9826
rect 41244 9214 41246 9266
rect 41298 9214 41300 9266
rect 40460 9202 40516 9212
rect 41244 9202 41300 9214
rect 41356 9380 41412 9390
rect 41356 9042 41412 9324
rect 41356 8990 41358 9042
rect 41410 8990 41412 9042
rect 41356 8978 41412 8990
rect 41468 9044 41524 9774
rect 41804 9266 41860 9884
rect 41804 9214 41806 9266
rect 41858 9214 41860 9266
rect 41804 9202 41860 9214
rect 42028 9828 42084 9838
rect 42028 9266 42084 9772
rect 42028 9214 42030 9266
rect 42082 9214 42084 9266
rect 42028 9202 42084 9214
rect 42140 9380 42196 9390
rect 41468 8708 41524 8988
rect 41244 8652 41524 8708
rect 41916 8930 41972 8942
rect 41916 8878 41918 8930
rect 41970 8878 41972 8930
rect 40908 8372 40964 8382
rect 40012 7812 40068 7822
rect 40012 7586 40068 7756
rect 40012 7534 40014 7586
rect 40066 7534 40068 7586
rect 40012 7522 40068 7534
rect 40124 7700 40180 7710
rect 39900 7196 40068 7252
rect 39676 7084 39956 7140
rect 39452 6750 39454 6802
rect 39506 6750 39508 6802
rect 39452 6738 39508 6750
rect 39788 6916 39844 6926
rect 39452 6580 39508 6590
rect 39452 6018 39508 6524
rect 39452 5966 39454 6018
rect 39506 5966 39508 6018
rect 39452 5954 39508 5966
rect 39788 4900 39844 6860
rect 39900 6130 39956 7084
rect 39900 6078 39902 6130
rect 39954 6078 39956 6130
rect 39900 6066 39956 6078
rect 40012 6130 40068 7196
rect 40012 6078 40014 6130
rect 40066 6078 40068 6130
rect 40012 6066 40068 6078
rect 40124 6018 40180 7644
rect 40908 7586 40964 8316
rect 40908 7534 40910 7586
rect 40962 7534 40964 7586
rect 40908 7522 40964 7534
rect 41244 7474 41300 8652
rect 41356 8484 41412 8494
rect 41412 8428 41524 8484
rect 41356 8418 41412 8428
rect 41244 7422 41246 7474
rect 41298 7422 41300 7474
rect 41244 7410 41300 7422
rect 41356 8258 41412 8270
rect 41356 8206 41358 8258
rect 41410 8206 41412 8258
rect 41132 7364 41188 7374
rect 41132 7270 41188 7308
rect 40124 5966 40126 6018
rect 40178 5966 40180 6018
rect 40124 5954 40180 5966
rect 41244 7252 41300 7262
rect 41244 5906 41300 7196
rect 41244 5854 41246 5906
rect 41298 5854 41300 5906
rect 41244 5842 41300 5854
rect 40348 5796 40404 5806
rect 39900 5124 39956 5134
rect 40348 5124 40404 5740
rect 41020 5796 41076 5806
rect 41020 5684 41076 5740
rect 41356 5796 41412 8206
rect 41468 6356 41524 8428
rect 41916 7700 41972 8878
rect 42140 8596 42196 9324
rect 41916 7634 41972 7644
rect 42028 8540 42196 8596
rect 41580 7476 41636 7486
rect 41580 7382 41636 7420
rect 42028 7474 42084 8540
rect 42140 8148 42196 8158
rect 42140 8054 42196 8092
rect 42028 7422 42030 7474
rect 42082 7422 42084 7474
rect 42028 7410 42084 7422
rect 42252 7476 42308 10556
rect 42588 10500 42644 10510
rect 42588 10406 42644 10444
rect 42588 10052 42644 10062
rect 42476 9602 42532 9614
rect 42476 9550 42478 9602
rect 42530 9550 42532 9602
rect 42476 9492 42532 9550
rect 42476 9426 42532 9436
rect 42476 9268 42532 9278
rect 42364 8818 42420 8830
rect 42364 8766 42366 8818
rect 42418 8766 42420 8818
rect 42364 7698 42420 8766
rect 42364 7646 42366 7698
rect 42418 7646 42420 7698
rect 42364 7634 42420 7646
rect 42476 7698 42532 9212
rect 42588 8932 42644 9996
rect 42588 8838 42644 8876
rect 42924 8930 42980 10668
rect 42924 8878 42926 8930
rect 42978 8878 42980 8930
rect 42700 8820 42756 8830
rect 42924 8820 42980 8878
rect 42700 8818 42980 8820
rect 42700 8766 42702 8818
rect 42754 8766 42980 8818
rect 42700 8764 42980 8766
rect 42700 8754 42756 8764
rect 42812 8036 42868 8046
rect 42588 7812 42644 7822
rect 42644 7756 42756 7812
rect 42588 7746 42644 7756
rect 42476 7646 42478 7698
rect 42530 7646 42532 7698
rect 42476 7634 42532 7646
rect 42588 7476 42644 7486
rect 42252 7474 42644 7476
rect 42252 7422 42590 7474
rect 42642 7422 42644 7474
rect 42252 7420 42644 7422
rect 42588 7410 42644 7420
rect 41692 7362 41748 7374
rect 41692 7310 41694 7362
rect 41746 7310 41748 7362
rect 41580 6804 41636 6814
rect 41692 6804 41748 7310
rect 42476 6804 42532 6814
rect 41580 6802 41972 6804
rect 41580 6750 41582 6802
rect 41634 6750 41972 6802
rect 41580 6748 41972 6750
rect 41580 6738 41636 6748
rect 41916 6690 41972 6748
rect 42476 6710 42532 6748
rect 41916 6638 41918 6690
rect 41970 6638 41972 6690
rect 41916 6626 41972 6638
rect 42588 6692 42644 6702
rect 42700 6692 42756 7756
rect 42588 6690 42756 6692
rect 42588 6638 42590 6690
rect 42642 6638 42756 6690
rect 42588 6636 42756 6638
rect 42588 6626 42644 6636
rect 42140 6580 42196 6590
rect 42140 6486 42196 6524
rect 42700 6578 42756 6636
rect 42700 6526 42702 6578
rect 42754 6526 42756 6578
rect 42700 6514 42756 6526
rect 42364 6468 42420 6478
rect 42364 6374 42420 6412
rect 41468 6300 41748 6356
rect 41356 5730 41412 5740
rect 39900 5122 40404 5124
rect 39900 5070 39902 5122
rect 39954 5070 40350 5122
rect 40402 5070 40404 5122
rect 39900 5068 40404 5070
rect 39900 5058 39956 5068
rect 40348 5058 40404 5068
rect 40908 5628 41076 5684
rect 39788 4834 39844 4844
rect 39340 3714 39396 3724
rect 40572 4564 40628 4574
rect 38892 3666 39060 3668
rect 38892 3614 38894 3666
rect 38946 3614 39060 3666
rect 38892 3612 39060 3614
rect 38892 3602 38948 3612
rect 39788 3556 39844 3566
rect 39788 3462 39844 3500
rect 40572 800 40628 4508
rect 40908 4338 40964 5628
rect 41020 5012 41076 5022
rect 41020 4918 41076 4956
rect 41692 4450 41748 6300
rect 41692 4398 41694 4450
rect 41746 4398 41748 4450
rect 41692 4386 41748 4398
rect 40908 4286 40910 4338
rect 40962 4286 40964 4338
rect 40908 4274 40964 4286
rect 40796 3668 40852 3678
rect 40796 3574 40852 3612
rect 42812 3554 42868 7980
rect 43036 7474 43092 11340
rect 43036 7422 43038 7474
rect 43090 7422 43092 7474
rect 43036 7252 43092 7422
rect 43260 7252 43316 11452
rect 43484 11394 43540 11788
rect 43596 11620 43652 11902
rect 43708 11956 43764 13356
rect 43820 12962 43876 15932
rect 44716 15148 44772 16828
rect 45164 17554 45332 17556
rect 45164 17502 45278 17554
rect 45330 17502 45332 17554
rect 45164 17500 45332 17502
rect 44940 16548 44996 16558
rect 44716 15092 44884 15148
rect 44828 14980 44884 15092
rect 44268 14530 44324 14542
rect 44268 14478 44270 14530
rect 44322 14478 44324 14530
rect 44156 13634 44212 13646
rect 44156 13582 44158 13634
rect 44210 13582 44212 13634
rect 44156 13524 44212 13582
rect 44268 13636 44324 14478
rect 44492 13860 44548 13870
rect 44268 13570 44324 13580
rect 44380 13804 44492 13860
rect 44156 13458 44212 13468
rect 43820 12910 43822 12962
rect 43874 12910 43876 12962
rect 43820 12898 43876 12910
rect 44044 12962 44100 12974
rect 44044 12910 44046 12962
rect 44098 12910 44100 12962
rect 44044 12852 44100 12910
rect 44044 12786 44100 12796
rect 43708 11890 43764 11900
rect 44044 12066 44100 12078
rect 44044 12014 44046 12066
rect 44098 12014 44100 12066
rect 43596 11554 43652 11564
rect 43484 11342 43486 11394
rect 43538 11342 43540 11394
rect 43484 11284 43540 11342
rect 43484 11218 43540 11228
rect 43708 11282 43764 11294
rect 43708 11230 43710 11282
rect 43762 11230 43764 11282
rect 43708 10500 43764 11230
rect 43820 11284 43876 11294
rect 43820 11190 43876 11228
rect 44044 10724 44100 12014
rect 44268 11956 44324 11966
rect 44268 11862 44324 11900
rect 44268 11620 44324 11630
rect 44268 11526 44324 11564
rect 44044 10658 44100 10668
rect 43708 10434 43764 10444
rect 43372 10388 43428 10398
rect 43372 8036 43428 10332
rect 43372 7970 43428 7980
rect 44268 8370 44324 8382
rect 44268 8318 44270 8370
rect 44322 8318 44324 8370
rect 43260 7196 43428 7252
rect 43036 7186 43092 7196
rect 43036 6916 43092 6926
rect 43372 6916 43428 7196
rect 43036 6692 43092 6860
rect 43260 6860 43428 6916
rect 43484 6916 43540 6926
rect 43540 6860 43652 6916
rect 43260 6802 43316 6860
rect 43484 6850 43540 6860
rect 43260 6750 43262 6802
rect 43314 6750 43316 6802
rect 43260 6738 43316 6750
rect 42924 6690 43092 6692
rect 42924 6638 43038 6690
rect 43090 6638 43092 6690
rect 42924 6636 43092 6638
rect 42924 6578 42980 6636
rect 43036 6626 43092 6636
rect 42924 6526 42926 6578
rect 42978 6526 42980 6578
rect 42924 6514 42980 6526
rect 43484 6580 43540 6590
rect 43036 6468 43092 6478
rect 42924 5796 42980 5806
rect 42924 5702 42980 5740
rect 43036 5236 43092 6412
rect 43260 6468 43316 6478
rect 43260 6374 43316 6412
rect 43484 6466 43540 6524
rect 43484 6414 43486 6466
rect 43538 6414 43540 6466
rect 43148 5236 43204 5246
rect 43036 5180 43148 5236
rect 43148 5142 43204 5180
rect 43484 4788 43540 6414
rect 43596 5122 43652 6860
rect 43596 5070 43598 5122
rect 43650 5070 43652 5122
rect 43596 5058 43652 5070
rect 43708 6578 43764 6590
rect 43708 6526 43710 6578
rect 43762 6526 43764 6578
rect 43708 5122 43764 6526
rect 44156 6580 44212 6590
rect 44268 6580 44324 8318
rect 44156 6578 44324 6580
rect 44156 6526 44158 6578
rect 44210 6526 44324 6578
rect 44156 6524 44324 6526
rect 44156 6514 44212 6524
rect 44044 6466 44100 6478
rect 44044 6414 44046 6466
rect 44098 6414 44100 6466
rect 43708 5070 43710 5122
rect 43762 5070 43764 5122
rect 43484 4722 43540 4732
rect 43708 4228 43764 5070
rect 43820 6244 43876 6254
rect 43820 5122 43876 6188
rect 44044 6020 44100 6414
rect 44044 5954 44100 5964
rect 44268 6020 44324 6524
rect 44268 5954 44324 5964
rect 43820 5070 43822 5122
rect 43874 5070 43876 5122
rect 43820 5058 43876 5070
rect 44044 5236 44100 5246
rect 44044 5122 44100 5180
rect 44380 5236 44436 13804
rect 44492 13794 44548 13804
rect 44828 13636 44884 14924
rect 44940 14642 44996 16492
rect 45052 15876 45108 15886
rect 45052 15782 45108 15820
rect 45164 14980 45220 17500
rect 45276 17490 45332 17500
rect 45612 17442 45668 17454
rect 45612 17390 45614 17442
rect 45666 17390 45668 17442
rect 45388 16996 45444 17006
rect 45612 16996 45668 17390
rect 45836 17444 45892 17454
rect 45836 17350 45892 17388
rect 45388 16994 45668 16996
rect 45388 16942 45390 16994
rect 45442 16942 45668 16994
rect 45388 16940 45668 16942
rect 45388 16930 45444 16940
rect 45948 16772 46004 17612
rect 45948 16212 46004 16716
rect 45836 16210 46004 16212
rect 45836 16158 45950 16210
rect 46002 16158 46004 16210
rect 45836 16156 46004 16158
rect 45164 14924 45556 14980
rect 44940 14590 44942 14642
rect 44994 14590 44996 14642
rect 44940 14578 44996 14590
rect 45500 14642 45556 14924
rect 45500 14590 45502 14642
rect 45554 14590 45556 14642
rect 45500 14578 45556 14590
rect 45388 14532 45444 14542
rect 45388 14438 45444 14476
rect 45724 14532 45780 14542
rect 45836 14532 45892 16156
rect 45948 16146 46004 16156
rect 46060 15988 46116 19852
rect 46172 20018 46228 20030
rect 46172 19966 46174 20018
rect 46226 19966 46228 20018
rect 46172 19012 46228 19966
rect 46284 19234 46340 20076
rect 46284 19182 46286 19234
rect 46338 19182 46340 19234
rect 46284 19170 46340 19182
rect 46172 18946 46228 18956
rect 46172 18452 46228 18462
rect 46172 18450 46340 18452
rect 46172 18398 46174 18450
rect 46226 18398 46340 18450
rect 46172 18396 46340 18398
rect 46172 18386 46228 18396
rect 46284 17668 46340 18396
rect 46284 17574 46340 17612
rect 46396 17108 46452 21532
rect 46732 21588 46788 21598
rect 46732 21494 46788 21532
rect 47516 21588 47572 21598
rect 47516 21494 47572 21532
rect 48636 21588 48692 21598
rect 48748 21588 48804 21598
rect 48692 21586 48804 21588
rect 48692 21534 48750 21586
rect 48802 21534 48804 21586
rect 48692 21532 48804 21534
rect 47404 21474 47460 21486
rect 47404 21422 47406 21474
rect 47458 21422 47460 21474
rect 47404 21028 47460 21422
rect 47068 20972 47460 21028
rect 47068 20914 47124 20972
rect 47068 20862 47070 20914
rect 47122 20862 47124 20914
rect 47068 20850 47124 20862
rect 46844 20804 46900 20814
rect 46732 20130 46788 20142
rect 46732 20078 46734 20130
rect 46786 20078 46788 20130
rect 46620 20018 46676 20030
rect 46620 19966 46622 20018
rect 46674 19966 46676 20018
rect 46508 18564 46564 18574
rect 46508 18470 46564 18508
rect 46620 18340 46676 19966
rect 46732 20020 46788 20078
rect 46732 18450 46788 19964
rect 46732 18398 46734 18450
rect 46786 18398 46788 18450
rect 46732 18386 46788 18398
rect 46620 18274 46676 18284
rect 46844 18116 46900 20748
rect 47068 20244 47124 20254
rect 47068 19346 47124 20188
rect 47404 20132 47460 20142
rect 47404 20130 47572 20132
rect 47404 20078 47406 20130
rect 47458 20078 47572 20130
rect 47404 20076 47572 20078
rect 47404 20066 47460 20076
rect 47068 19294 47070 19346
rect 47122 19294 47124 19346
rect 47068 19282 47124 19294
rect 47516 18562 47572 20076
rect 47852 20018 47908 20030
rect 47852 19966 47854 20018
rect 47906 19966 47908 20018
rect 47852 19348 47908 19966
rect 47852 19282 47908 19292
rect 48188 20018 48244 20030
rect 48188 19966 48190 20018
rect 48242 19966 48244 20018
rect 47516 18510 47518 18562
rect 47570 18510 47572 18562
rect 47516 18498 47572 18510
rect 47852 19012 47908 19022
rect 47068 18228 47124 18238
rect 46956 18226 47124 18228
rect 46956 18174 47070 18226
rect 47122 18174 47124 18226
rect 46956 18172 47124 18174
rect 46956 18116 47012 18172
rect 47068 18162 47124 18172
rect 46396 17042 46452 17052
rect 46732 18060 47012 18116
rect 45724 14530 45892 14532
rect 45724 14478 45726 14530
rect 45778 14478 45892 14530
rect 45724 14476 45892 14478
rect 45948 15932 46116 15988
rect 46284 16098 46340 16110
rect 46284 16046 46286 16098
rect 46338 16046 46340 16098
rect 45948 14530 46004 15932
rect 46060 15202 46116 15214
rect 46060 15150 46062 15202
rect 46114 15150 46116 15202
rect 46060 14980 46116 15150
rect 46284 15148 46340 16046
rect 46284 15092 46452 15148
rect 46116 14924 46340 14980
rect 46060 14914 46116 14924
rect 45948 14478 45950 14530
rect 46002 14478 46004 14530
rect 45724 14466 45780 14476
rect 45948 14466 46004 14478
rect 46284 14530 46340 14924
rect 46284 14478 46286 14530
rect 46338 14478 46340 14530
rect 46284 14466 46340 14478
rect 45052 14308 45108 14318
rect 45836 14308 45892 14318
rect 45052 14306 45220 14308
rect 45052 14254 45054 14306
rect 45106 14254 45220 14306
rect 45052 14252 45220 14254
rect 45052 14242 45108 14252
rect 44604 11954 44660 11966
rect 44604 11902 44606 11954
rect 44658 11902 44660 11954
rect 44604 10724 44660 11902
rect 44492 10164 44548 10174
rect 44492 5908 44548 10108
rect 44604 9828 44660 10668
rect 44716 11732 44772 11742
rect 44716 10722 44772 11676
rect 44828 11394 44884 13580
rect 44940 13524 44996 13534
rect 44996 13468 45108 13524
rect 44940 13458 44996 13468
rect 45052 13186 45108 13468
rect 45052 13134 45054 13186
rect 45106 13134 45108 13186
rect 45052 13122 45108 13134
rect 45164 13076 45220 14252
rect 45500 13188 45556 13198
rect 45164 13010 45220 13020
rect 45388 13132 45500 13188
rect 45388 13074 45444 13132
rect 45500 13122 45556 13132
rect 45836 13186 45892 14252
rect 46396 13972 46452 15092
rect 46732 14532 46788 18060
rect 47852 17892 47908 18956
rect 48188 18676 48244 19966
rect 48636 18676 48692 21532
rect 48748 21522 48804 21532
rect 48748 21362 48804 21374
rect 48748 21310 48750 21362
rect 48802 21310 48804 21362
rect 48748 20244 48804 21310
rect 48748 20178 48804 20188
rect 48748 20018 48804 20030
rect 48748 19966 48750 20018
rect 48802 19966 48804 20018
rect 48748 19908 48804 19966
rect 48748 19842 48804 19852
rect 48748 18900 48804 18910
rect 48804 18844 48916 18900
rect 48748 18834 48804 18844
rect 48748 18676 48804 18686
rect 48188 18674 48804 18676
rect 48188 18622 48750 18674
rect 48802 18622 48804 18674
rect 48188 18620 48804 18622
rect 48748 18610 48804 18620
rect 47964 18452 48020 18462
rect 47964 18450 48132 18452
rect 47964 18398 47966 18450
rect 48018 18398 48132 18450
rect 47964 18396 48132 18398
rect 47964 18386 48020 18396
rect 47852 17826 47908 17836
rect 47068 17556 47124 17566
rect 47068 17554 47908 17556
rect 47068 17502 47070 17554
rect 47122 17502 47908 17554
rect 47068 17500 47908 17502
rect 47068 17490 47124 17500
rect 47516 16772 47572 16782
rect 47516 16678 47572 16716
rect 47852 16770 47908 17500
rect 47964 17108 48020 17118
rect 47964 17014 48020 17052
rect 47852 16718 47854 16770
rect 47906 16718 47908 16770
rect 47852 16706 47908 16718
rect 47068 16548 47124 16558
rect 47068 16212 47124 16492
rect 48076 16324 48132 18396
rect 48636 17892 48692 17902
rect 48524 17836 48636 17892
rect 48188 16660 48244 16670
rect 48188 16658 48356 16660
rect 48188 16606 48190 16658
rect 48242 16606 48356 16658
rect 48188 16604 48356 16606
rect 48188 16594 48244 16604
rect 48188 16324 48244 16334
rect 48076 16322 48244 16324
rect 48076 16270 48190 16322
rect 48242 16270 48244 16322
rect 48076 16268 48244 16270
rect 47068 16098 47124 16156
rect 47068 16046 47070 16098
rect 47122 16046 47124 16098
rect 47068 16034 47124 16046
rect 47292 16098 47348 16110
rect 47292 16046 47294 16098
rect 47346 16046 47348 16098
rect 46732 14466 46788 14476
rect 46844 15986 46900 15998
rect 46844 15934 46846 15986
rect 46898 15934 46900 15986
rect 46620 13972 46676 13982
rect 46396 13970 46676 13972
rect 46396 13918 46622 13970
rect 46674 13918 46676 13970
rect 46396 13916 46676 13918
rect 46284 13636 46340 13646
rect 46396 13636 46452 13916
rect 46620 13906 46676 13916
rect 46732 13972 46788 13982
rect 46284 13634 46452 13636
rect 46284 13582 46286 13634
rect 46338 13582 46452 13634
rect 46284 13580 46452 13582
rect 46284 13570 46340 13580
rect 45836 13134 45838 13186
rect 45890 13134 45892 13186
rect 45836 13122 45892 13134
rect 45388 13022 45390 13074
rect 45442 13022 45444 13074
rect 45388 13010 45444 13022
rect 46060 12964 46116 12974
rect 46060 12870 46116 12908
rect 46284 12962 46340 12974
rect 46284 12910 46286 12962
rect 46338 12910 46340 12962
rect 45164 12738 45220 12750
rect 45164 12686 45166 12738
rect 45218 12686 45220 12738
rect 45164 12516 45220 12686
rect 46172 12740 46228 12750
rect 46172 12646 46228 12684
rect 45388 12628 45444 12638
rect 45444 12572 45556 12628
rect 45388 12562 45444 12572
rect 45164 12450 45220 12460
rect 45276 12292 45332 12302
rect 45052 12290 45332 12292
rect 45052 12238 45278 12290
rect 45330 12238 45332 12290
rect 45052 12236 45332 12238
rect 44828 11342 44830 11394
rect 44882 11342 44884 11394
rect 44828 11330 44884 11342
rect 44940 12178 44996 12190
rect 44940 12126 44942 12178
rect 44994 12126 44996 12178
rect 44716 10670 44718 10722
rect 44770 10670 44772 10722
rect 44716 10658 44772 10670
rect 44940 10164 44996 12126
rect 44604 9762 44660 9772
rect 44716 10108 44996 10164
rect 44716 6132 44772 10108
rect 45052 10052 45108 12236
rect 45276 12226 45332 12236
rect 45388 11284 45444 11294
rect 45388 10612 45444 11228
rect 45500 10836 45556 12572
rect 46284 12404 46340 12910
rect 46620 12850 46676 12862
rect 46620 12798 46622 12850
rect 46674 12798 46676 12850
rect 46284 12338 46340 12348
rect 46508 12516 46564 12526
rect 46508 12402 46564 12460
rect 46508 12350 46510 12402
rect 46562 12350 46564 12402
rect 46508 12338 46564 12350
rect 45836 12290 45892 12302
rect 45836 12238 45838 12290
rect 45890 12238 45892 12290
rect 45836 12180 45892 12238
rect 46620 12292 46676 12798
rect 46732 12516 46788 13916
rect 46844 13188 46900 15934
rect 47292 15148 47348 16046
rect 46956 15092 47348 15148
rect 46956 13858 47012 15092
rect 47740 14644 47796 14654
rect 46956 13806 46958 13858
rect 47010 13806 47012 13858
rect 46956 13748 47012 13806
rect 46956 13682 47012 13692
rect 47068 14418 47124 14430
rect 47068 14366 47070 14418
rect 47122 14366 47124 14418
rect 46844 13122 46900 13132
rect 47068 12740 47124 14366
rect 47740 13860 47796 14588
rect 48188 13972 48244 16268
rect 48300 15764 48356 16604
rect 48412 16212 48468 16222
rect 48412 16118 48468 16156
rect 48524 15988 48580 17836
rect 48636 17826 48692 17836
rect 48860 17332 48916 18844
rect 48748 17276 48916 17332
rect 48972 18450 49028 21868
rect 49084 21362 49140 21374
rect 49084 21310 49086 21362
rect 49138 21310 49140 21362
rect 49084 20132 49140 21310
rect 49196 20914 49252 21868
rect 49196 20862 49198 20914
rect 49250 20862 49252 20914
rect 49196 20850 49252 20862
rect 49420 21700 49476 23492
rect 49084 20038 49140 20076
rect 49196 19348 49252 19358
rect 49196 18788 49252 19292
rect 48972 18398 48974 18450
rect 49026 18398 49028 18450
rect 48748 16772 48804 17276
rect 48860 17108 48916 17118
rect 48972 17108 49028 18398
rect 48860 17106 49028 17108
rect 48860 17054 48862 17106
rect 48914 17054 49028 17106
rect 48860 17052 49028 17054
rect 49084 18732 49252 18788
rect 48860 17042 48916 17052
rect 49084 16994 49140 18732
rect 49196 17892 49252 17902
rect 49196 17778 49252 17836
rect 49196 17726 49198 17778
rect 49250 17726 49252 17778
rect 49196 17714 49252 17726
rect 49084 16942 49086 16994
rect 49138 16942 49140 16994
rect 49084 16930 49140 16942
rect 48748 16770 48916 16772
rect 48748 16718 48750 16770
rect 48802 16718 48916 16770
rect 48748 16716 48916 16718
rect 48748 16706 48804 16716
rect 48860 16098 48916 16716
rect 48860 16046 48862 16098
rect 48914 16046 48916 16098
rect 48860 16034 48916 16046
rect 49084 16660 49140 16670
rect 48636 15988 48692 15998
rect 48524 15986 48692 15988
rect 48524 15934 48638 15986
rect 48690 15934 48692 15986
rect 48524 15932 48692 15934
rect 48636 15922 48692 15932
rect 48748 15874 48804 15886
rect 48748 15822 48750 15874
rect 48802 15822 48804 15874
rect 48748 15764 48804 15822
rect 48300 15708 48804 15764
rect 48860 15426 48916 15438
rect 48860 15374 48862 15426
rect 48914 15374 48916 15426
rect 48860 15316 48916 15374
rect 48860 15250 48916 15260
rect 49084 15314 49140 16604
rect 49084 15262 49086 15314
rect 49138 15262 49140 15314
rect 49084 14868 49140 15262
rect 49084 14802 49140 14812
rect 49196 14644 49252 14654
rect 49196 14550 49252 14588
rect 48300 13972 48356 13982
rect 48188 13970 48356 13972
rect 48188 13918 48302 13970
rect 48354 13918 48356 13970
rect 48188 13916 48356 13918
rect 48300 13906 48356 13916
rect 48860 13860 48916 13870
rect 47740 13858 48020 13860
rect 47740 13806 47742 13858
rect 47794 13806 48020 13858
rect 47740 13804 48020 13806
rect 47740 13794 47796 13804
rect 47516 13748 47572 13758
rect 47516 13746 47684 13748
rect 47516 13694 47518 13746
rect 47570 13694 47684 13746
rect 47516 13692 47684 13694
rect 47516 13682 47572 13692
rect 47292 13634 47348 13646
rect 47292 13582 47294 13634
rect 47346 13582 47348 13634
rect 47292 12964 47348 13582
rect 47628 13076 47684 13692
rect 47964 13524 48020 13804
rect 48860 13766 48916 13804
rect 48972 13858 49028 13870
rect 48972 13806 48974 13858
rect 49026 13806 49028 13858
rect 48076 13748 48132 13758
rect 48748 13748 48804 13758
rect 48132 13692 48244 13748
rect 48076 13654 48132 13692
rect 47964 13188 48020 13468
rect 47964 13132 48132 13188
rect 47852 13076 47908 13086
rect 47628 13020 47796 13076
rect 47516 12964 47572 12974
rect 47292 12962 47460 12964
rect 47292 12910 47294 12962
rect 47346 12910 47460 12962
rect 47292 12908 47460 12910
rect 47292 12898 47348 12908
rect 47068 12674 47124 12684
rect 46732 12460 47012 12516
rect 46732 12292 46788 12302
rect 46620 12290 46788 12292
rect 46620 12238 46734 12290
rect 46786 12238 46788 12290
rect 46620 12236 46788 12238
rect 46732 12226 46788 12236
rect 45836 12114 45892 12124
rect 46060 12180 46116 12190
rect 46060 12178 46676 12180
rect 46060 12126 46062 12178
rect 46114 12126 46676 12178
rect 46060 12124 46676 12126
rect 46060 12114 46116 12124
rect 45948 12068 46004 12078
rect 45948 11974 46004 12012
rect 46396 11956 46452 11966
rect 46060 11954 46452 11956
rect 46060 11902 46398 11954
rect 46450 11902 46452 11954
rect 46060 11900 46452 11902
rect 46060 11620 46116 11900
rect 46396 11890 46452 11900
rect 45612 11564 46116 11620
rect 45612 11506 45668 11564
rect 45612 11454 45614 11506
rect 45666 11454 45668 11506
rect 45612 11442 45668 11454
rect 45836 10836 45892 10846
rect 45500 10834 45892 10836
rect 45500 10782 45838 10834
rect 45890 10782 45892 10834
rect 45500 10780 45892 10782
rect 45836 10770 45892 10780
rect 45276 10388 45332 10398
rect 44940 9996 45108 10052
rect 45164 10332 45276 10388
rect 44828 9940 44884 9950
rect 44828 9846 44884 9884
rect 44940 8820 44996 9996
rect 45052 9828 45108 9838
rect 45052 9734 45108 9772
rect 45052 9156 45108 9166
rect 45164 9156 45220 10332
rect 45276 10322 45332 10332
rect 45388 10050 45444 10556
rect 45388 9998 45390 10050
rect 45442 9998 45444 10050
rect 45388 9986 45444 9998
rect 45500 10610 45556 10622
rect 45500 10558 45502 10610
rect 45554 10558 45556 10610
rect 45052 9154 45220 9156
rect 45052 9102 45054 9154
rect 45106 9102 45220 9154
rect 45052 9100 45220 9102
rect 45052 9090 45108 9100
rect 45500 9044 45556 10558
rect 46060 10612 46116 10622
rect 46060 10518 46116 10556
rect 46508 10386 46564 10398
rect 46508 10334 46510 10386
rect 46562 10334 46564 10386
rect 46284 9826 46340 9838
rect 46284 9774 46286 9826
rect 46338 9774 46340 9826
rect 45836 9604 45892 9614
rect 45892 9548 46004 9604
rect 45836 9510 45892 9548
rect 45836 9044 45892 9054
rect 45500 9042 45892 9044
rect 45500 8990 45838 9042
rect 45890 8990 45892 9042
rect 45500 8988 45892 8990
rect 45500 8820 45556 8830
rect 44940 8764 45500 8820
rect 45500 8258 45556 8764
rect 45500 8206 45502 8258
rect 45554 8206 45556 8258
rect 45500 8194 45556 8206
rect 45276 8148 45332 8158
rect 45164 8146 45332 8148
rect 45164 8094 45278 8146
rect 45330 8094 45332 8146
rect 45164 8092 45332 8094
rect 44940 8036 44996 8046
rect 44940 8034 45108 8036
rect 44940 7982 44942 8034
rect 44994 7982 45108 8034
rect 44940 7980 45108 7982
rect 44940 7970 44996 7980
rect 44828 6692 44884 6702
rect 44828 6244 44884 6636
rect 44828 6178 44884 6188
rect 44940 6466 44996 6478
rect 44940 6414 44942 6466
rect 44994 6414 44996 6466
rect 44716 6066 44772 6076
rect 44492 5852 44772 5908
rect 44380 5170 44436 5180
rect 44044 5070 44046 5122
rect 44098 5070 44100 5122
rect 44044 5058 44100 5070
rect 43932 4898 43988 4910
rect 43932 4846 43934 4898
rect 43986 4846 43988 4898
rect 43932 4788 43988 4846
rect 43932 4722 43988 4732
rect 44156 4900 44212 4910
rect 44156 4450 44212 4844
rect 44156 4398 44158 4450
rect 44210 4398 44212 4450
rect 44156 4386 44212 4398
rect 44380 4452 44436 4462
rect 44380 4358 44436 4396
rect 43820 4228 43876 4238
rect 43708 4226 43876 4228
rect 43708 4174 43822 4226
rect 43874 4174 43876 4226
rect 43708 4172 43876 4174
rect 43820 4162 43876 4172
rect 44268 4226 44324 4238
rect 44268 4174 44270 4226
rect 44322 4174 44324 4226
rect 44268 3780 44324 4174
rect 42812 3502 42814 3554
rect 42866 3502 42868 3554
rect 42812 3490 42868 3502
rect 43932 3724 44324 3780
rect 44492 3892 44548 3902
rect 43036 3444 43092 3454
rect 43036 3350 43092 3388
rect 42364 3332 42420 3342
rect 42364 800 42420 3276
rect 43932 3220 43988 3724
rect 44044 3556 44100 3566
rect 44044 3462 44100 3500
rect 44492 3388 44548 3836
rect 44716 3666 44772 5852
rect 44828 4898 44884 4910
rect 44828 4846 44830 4898
rect 44882 4846 44884 4898
rect 44828 4564 44884 4846
rect 44940 4900 44996 6414
rect 45052 5684 45108 7980
rect 45164 6468 45220 8092
rect 45276 8082 45332 8092
rect 45612 8034 45668 8046
rect 45612 7982 45614 8034
rect 45666 7982 45668 8034
rect 45612 7588 45668 7982
rect 45724 8036 45780 8046
rect 45724 7942 45780 7980
rect 45612 7522 45668 7532
rect 45724 7364 45780 7374
rect 45836 7364 45892 8988
rect 45948 8932 46004 9548
rect 45948 8866 46004 8876
rect 45948 8484 46004 8494
rect 45948 8258 46004 8428
rect 45948 8206 45950 8258
rect 46002 8206 46004 8258
rect 45948 8194 46004 8206
rect 46284 8258 46340 9774
rect 46508 9268 46564 10334
rect 46620 9268 46676 12124
rect 46732 10724 46788 10734
rect 46732 10630 46788 10668
rect 46956 10500 47012 12460
rect 47068 12068 47124 12078
rect 47124 12012 47236 12068
rect 47068 12002 47124 12012
rect 46956 10434 47012 10444
rect 46844 10388 46900 10398
rect 46844 10294 46900 10332
rect 47068 9940 47124 9950
rect 47068 9846 47124 9884
rect 46732 9268 46788 9278
rect 47180 9268 47236 12012
rect 47404 11508 47460 12908
rect 47516 12962 47684 12964
rect 47516 12910 47518 12962
rect 47570 12910 47684 12962
rect 47516 12908 47684 12910
rect 47516 12898 47572 12908
rect 47516 12404 47572 12414
rect 47516 12066 47572 12348
rect 47516 12014 47518 12066
rect 47570 12014 47572 12066
rect 47516 12002 47572 12014
rect 47628 11732 47684 12908
rect 47740 12292 47796 13020
rect 47740 12178 47796 12236
rect 47740 12126 47742 12178
rect 47794 12126 47796 12178
rect 47740 12114 47796 12126
rect 47628 11666 47684 11676
rect 47740 11508 47796 11518
rect 47404 11506 47796 11508
rect 47404 11454 47742 11506
rect 47794 11454 47796 11506
rect 47404 11452 47796 11454
rect 47740 11442 47796 11452
rect 47292 11396 47348 11406
rect 47852 11396 47908 13020
rect 47964 12964 48020 12974
rect 47964 12292 48020 12908
rect 48076 12962 48132 13132
rect 48076 12910 48078 12962
rect 48130 12910 48132 12962
rect 48076 12898 48132 12910
rect 48188 12850 48244 13692
rect 48412 13746 48804 13748
rect 48412 13694 48750 13746
rect 48802 13694 48804 13746
rect 48412 13692 48804 13694
rect 48300 13076 48356 13086
rect 48300 12962 48356 13020
rect 48300 12910 48302 12962
rect 48354 12910 48356 12962
rect 48300 12898 48356 12910
rect 48188 12798 48190 12850
rect 48242 12798 48244 12850
rect 48188 12628 48244 12798
rect 48188 12572 48356 12628
rect 47964 12236 48132 12292
rect 47964 11954 48020 11966
rect 47964 11902 47966 11954
rect 48018 11902 48020 11954
rect 47964 11620 48020 11902
rect 47964 11554 48020 11564
rect 48076 11508 48132 12236
rect 48188 11508 48244 11518
rect 48076 11506 48244 11508
rect 48076 11454 48190 11506
rect 48242 11454 48244 11506
rect 48076 11452 48244 11454
rect 48188 11442 48244 11452
rect 47964 11396 48020 11406
rect 47348 11340 47460 11396
rect 47852 11394 48020 11396
rect 47852 11342 47966 11394
rect 48018 11342 48020 11394
rect 47852 11340 48020 11342
rect 47292 11330 47348 11340
rect 47292 10722 47348 10734
rect 47292 10670 47294 10722
rect 47346 10670 47348 10722
rect 47292 10276 47348 10670
rect 47292 10210 47348 10220
rect 47404 9268 47460 11340
rect 47964 11330 48020 11340
rect 48300 11394 48356 12572
rect 48300 11342 48302 11394
rect 48354 11342 48356 11394
rect 48300 11330 48356 11342
rect 48076 10836 48132 10846
rect 48076 10610 48132 10780
rect 48076 10558 48078 10610
rect 48130 10558 48132 10610
rect 48076 10546 48132 10558
rect 47628 10498 47684 10510
rect 47628 10446 47630 10498
rect 47682 10446 47684 10498
rect 47628 10388 47684 10446
rect 47628 10322 47684 10332
rect 47852 9380 47908 9390
rect 46620 9266 46788 9268
rect 46620 9214 46734 9266
rect 46786 9214 46788 9266
rect 46620 9212 46788 9214
rect 46508 9202 46564 9212
rect 46732 9202 46788 9212
rect 46956 9212 47236 9268
rect 47292 9212 47460 9268
rect 47740 9324 47852 9380
rect 47740 9266 47796 9324
rect 47852 9314 47908 9324
rect 47740 9214 47742 9266
rect 47794 9214 47796 9266
rect 46396 9156 46452 9166
rect 46396 9042 46452 9100
rect 46396 8990 46398 9042
rect 46450 8990 46452 9042
rect 46396 8484 46452 8990
rect 46620 9042 46676 9054
rect 46620 8990 46622 9042
rect 46674 8990 46676 9042
rect 46452 8428 46564 8484
rect 46396 8418 46452 8428
rect 46284 8206 46286 8258
rect 46338 8206 46340 8258
rect 45724 7362 45892 7364
rect 45724 7310 45726 7362
rect 45778 7310 45892 7362
rect 45724 7308 45892 7310
rect 45948 7700 46004 7710
rect 45388 7252 45444 7262
rect 45388 6802 45444 7196
rect 45388 6750 45390 6802
rect 45442 6750 45444 6802
rect 45388 6738 45444 6750
rect 45724 6692 45780 7308
rect 45612 6636 45780 6692
rect 45164 5908 45220 6412
rect 45164 5842 45220 5852
rect 45276 6580 45332 6590
rect 45052 5618 45108 5628
rect 44940 4834 44996 4844
rect 45276 5122 45332 6524
rect 45500 6578 45556 6590
rect 45500 6526 45502 6578
rect 45554 6526 45556 6578
rect 45388 6468 45444 6478
rect 45388 6244 45444 6412
rect 45388 6178 45444 6188
rect 45500 6020 45556 6526
rect 45612 6580 45668 6636
rect 45612 6514 45668 6524
rect 45948 6578 46004 7644
rect 45948 6526 45950 6578
rect 46002 6526 46004 6578
rect 45948 6514 46004 6526
rect 46284 6690 46340 8206
rect 46284 6638 46286 6690
rect 46338 6638 46340 6690
rect 46284 6580 46340 6638
rect 46284 6514 46340 6524
rect 46396 8036 46452 8046
rect 45724 6466 45780 6478
rect 45724 6414 45726 6466
rect 45778 6414 45780 6466
rect 45724 6132 45780 6414
rect 45724 6066 45780 6076
rect 46396 6020 46452 7980
rect 46508 6692 46564 8428
rect 46620 7700 46676 8990
rect 46844 9042 46900 9054
rect 46844 8990 46846 9042
rect 46898 8990 46900 9042
rect 46844 8820 46900 8990
rect 46620 7634 46676 7644
rect 46732 8764 46844 8820
rect 46508 6626 46564 6636
rect 46732 6130 46788 8764
rect 46844 8754 46900 8764
rect 46956 7924 47012 9212
rect 47068 9044 47124 9054
rect 47068 8950 47124 8988
rect 47292 8820 47348 9212
rect 47740 9202 47796 9214
rect 48076 9156 48132 9166
rect 47068 8764 47348 8820
rect 47404 9042 47460 9054
rect 47404 8990 47406 9042
rect 47458 8990 47460 9042
rect 47068 8370 47124 8764
rect 47068 8318 47070 8370
rect 47122 8318 47124 8370
rect 47068 8306 47124 8318
rect 46956 7868 47124 7924
rect 46956 7588 47012 7598
rect 46732 6078 46734 6130
rect 46786 6078 46788 6130
rect 46732 6066 46788 6078
rect 46844 7532 46956 7588
rect 46844 6130 46900 7532
rect 46956 7522 47012 7532
rect 47068 6690 47124 7868
rect 47404 7028 47460 8990
rect 47628 9042 47684 9054
rect 47628 8990 47630 9042
rect 47682 8990 47684 9042
rect 47628 8820 47684 8990
rect 47852 9044 47908 9054
rect 47852 8950 47908 8988
rect 48076 9042 48132 9100
rect 48076 8990 48078 9042
rect 48130 8990 48132 9042
rect 48076 8978 48132 8990
rect 47628 8754 47684 8764
rect 48412 7588 48468 13692
rect 48748 13682 48804 13692
rect 48524 13524 48580 13534
rect 48580 13468 48692 13524
rect 48524 13458 48580 13468
rect 48636 11394 48692 13468
rect 48748 12738 48804 12750
rect 48748 12686 48750 12738
rect 48802 12686 48804 12738
rect 48748 12404 48804 12686
rect 48804 12348 48916 12404
rect 48748 12338 48804 12348
rect 48860 12068 48916 12348
rect 48972 12180 49028 13806
rect 49196 12964 49252 12974
rect 49420 12964 49476 21644
rect 49196 12962 49476 12964
rect 49196 12910 49198 12962
rect 49250 12910 49476 12962
rect 49196 12908 49476 12910
rect 49644 20132 49700 20142
rect 49196 12898 49252 12908
rect 49084 12852 49140 12862
rect 49084 12758 49140 12796
rect 49644 12516 49700 20076
rect 49196 12292 49252 12302
rect 49252 12236 49364 12292
rect 49196 12226 49252 12236
rect 49084 12180 49140 12218
rect 48972 12124 49084 12180
rect 49084 12114 49140 12124
rect 48860 12012 49028 12068
rect 48748 11956 48804 11966
rect 48748 11954 48916 11956
rect 48748 11902 48750 11954
rect 48802 11902 48916 11954
rect 48748 11900 48916 11902
rect 48748 11890 48804 11900
rect 48636 11342 48638 11394
rect 48690 11342 48692 11394
rect 48636 11330 48692 11342
rect 48748 11620 48804 11630
rect 48748 10722 48804 11564
rect 48860 10948 48916 11900
rect 48972 11394 49028 12012
rect 49084 11956 49140 11966
rect 49084 11954 49252 11956
rect 49084 11902 49086 11954
rect 49138 11902 49252 11954
rect 49084 11900 49252 11902
rect 49084 11890 49140 11900
rect 49084 11732 49140 11742
rect 49084 11618 49140 11676
rect 49084 11566 49086 11618
rect 49138 11566 49140 11618
rect 49084 11554 49140 11566
rect 48972 11342 48974 11394
rect 49026 11342 49028 11394
rect 48972 11330 49028 11342
rect 49196 11396 49252 11900
rect 49196 11330 49252 11340
rect 49084 11172 49140 11182
rect 49308 11172 49364 12236
rect 49084 11170 49364 11172
rect 49084 11118 49086 11170
rect 49138 11118 49364 11170
rect 49084 11116 49364 11118
rect 49420 12180 49476 12190
rect 49084 11106 49140 11116
rect 48860 10892 49140 10948
rect 48748 10670 48750 10722
rect 48802 10670 48804 10722
rect 48748 10658 48804 10670
rect 48972 10724 49028 10734
rect 48972 10630 49028 10668
rect 48524 10500 48580 10510
rect 48580 10444 48692 10500
rect 48524 10434 48580 10444
rect 48412 7522 48468 7532
rect 47068 6638 47070 6690
rect 47122 6638 47124 6690
rect 47068 6626 47124 6638
rect 47180 6972 47460 7028
rect 47516 7476 47572 7486
rect 47180 6468 47236 6972
rect 47404 6804 47460 6814
rect 46844 6078 46846 6130
rect 46898 6078 46900 6130
rect 46844 6066 46900 6078
rect 46956 6412 47236 6468
rect 47292 6692 47348 6702
rect 46956 6130 47012 6412
rect 46956 6078 46958 6130
rect 47010 6078 47012 6130
rect 46508 6020 46564 6030
rect 46396 6018 46564 6020
rect 46396 5966 46510 6018
rect 46562 5966 46564 6018
rect 46396 5964 46564 5966
rect 45500 5954 45556 5964
rect 46060 5236 46116 5246
rect 46060 5142 46116 5180
rect 45276 5070 45278 5122
rect 45330 5070 45332 5122
rect 44828 4498 44884 4508
rect 44716 3614 44718 3666
rect 44770 3614 44772 3666
rect 44716 3602 44772 3614
rect 44828 4340 44884 4350
rect 45276 4340 45332 5070
rect 44828 4338 45332 4340
rect 44828 4286 44830 4338
rect 44882 4286 45332 4338
rect 44828 4284 45332 4286
rect 45948 4900 46004 4910
rect 44828 3556 44884 4284
rect 44828 3490 44884 3500
rect 45612 4226 45668 4238
rect 45612 4174 45614 4226
rect 45666 4174 45668 4226
rect 43932 3154 43988 3164
rect 44156 3332 44548 3388
rect 44156 800 44212 3332
rect 45612 2884 45668 4174
rect 45612 2818 45668 2828
rect 45948 800 46004 4844
rect 46508 4228 46564 5964
rect 46956 6020 47012 6078
rect 46956 5954 47012 5964
rect 46508 4162 46564 4172
rect 46844 5908 46900 5918
rect 46844 3666 46900 5852
rect 47180 5908 47236 5918
rect 47292 5908 47348 6636
rect 47180 5906 47348 5908
rect 47180 5854 47182 5906
rect 47234 5854 47348 5906
rect 47180 5852 47348 5854
rect 47180 5842 47236 5852
rect 47404 3778 47460 6748
rect 47516 6130 47572 7420
rect 47516 6078 47518 6130
rect 47570 6078 47572 6130
rect 47516 6066 47572 6078
rect 47740 6244 47796 6254
rect 47740 5906 47796 6188
rect 48636 6132 48692 10444
rect 48860 10498 48916 10510
rect 48860 10446 48862 10498
rect 48914 10446 48916 10498
rect 48860 9940 48916 10446
rect 48860 9874 48916 9884
rect 49084 9380 49140 10892
rect 49196 9938 49252 11116
rect 49196 9886 49198 9938
rect 49250 9886 49252 9938
rect 49196 9874 49252 9886
rect 49084 9314 49140 9324
rect 48748 9156 48804 9166
rect 48748 9062 48804 9100
rect 49084 9042 49140 9054
rect 49084 8990 49086 9042
rect 49138 8990 49140 9042
rect 48748 8932 48804 8942
rect 48748 7476 48804 8876
rect 48860 8148 48916 8158
rect 48860 7698 48916 8092
rect 48860 7646 48862 7698
rect 48914 7646 48916 7698
rect 48860 7634 48916 7646
rect 48972 7586 49028 7598
rect 48972 7534 48974 7586
rect 49026 7534 49028 7586
rect 48972 7476 49028 7534
rect 48748 7420 48916 7476
rect 48748 7252 48804 7262
rect 48748 7158 48804 7196
rect 48748 6132 48804 6142
rect 48636 6130 48804 6132
rect 48636 6078 48750 6130
rect 48802 6078 48804 6130
rect 48636 6076 48804 6078
rect 47740 5854 47742 5906
rect 47794 5854 47796 5906
rect 47740 5842 47796 5854
rect 48188 6020 48244 6030
rect 47628 5684 47684 5694
rect 47404 3726 47406 3778
rect 47458 3726 47460 3778
rect 47404 3714 47460 3726
rect 47516 5012 47572 5022
rect 46844 3614 46846 3666
rect 46898 3614 46900 3666
rect 46844 3602 46900 3614
rect 47516 3666 47572 4956
rect 47628 4004 47684 5628
rect 48188 5234 48244 5964
rect 48188 5182 48190 5234
rect 48242 5182 48244 5234
rect 48188 5170 48244 5182
rect 48076 4450 48132 4462
rect 48076 4398 48078 4450
rect 48130 4398 48132 4450
rect 47740 4228 47796 4238
rect 47740 4134 47796 4172
rect 47628 3948 47796 4004
rect 47516 3614 47518 3666
rect 47570 3614 47572 3666
rect 47516 3602 47572 3614
rect 47628 3780 47684 3790
rect 47628 3442 47684 3724
rect 47628 3390 47630 3442
rect 47682 3390 47684 3442
rect 47628 3378 47684 3390
rect 47740 800 47796 3948
rect 48076 3892 48132 4398
rect 48076 3826 48132 3836
rect 48636 3780 48692 6076
rect 48748 6066 48804 6076
rect 48748 5236 48804 5246
rect 48860 5236 48916 7420
rect 48972 7410 49028 7420
rect 48972 6468 49028 6478
rect 49084 6468 49140 8990
rect 49196 9044 49252 9054
rect 49196 8370 49252 8988
rect 49196 8318 49198 8370
rect 49250 8318 49252 8370
rect 49196 8306 49252 8318
rect 49196 7700 49252 7710
rect 49196 6802 49252 7644
rect 49308 7476 49364 7486
rect 49420 7476 49476 12124
rect 49644 10724 49700 12460
rect 49644 10658 49700 10668
rect 49364 7420 49476 7476
rect 49532 10276 49588 10286
rect 49308 7410 49364 7420
rect 49196 6750 49198 6802
rect 49250 6750 49252 6802
rect 49196 6738 49252 6750
rect 49028 6412 49140 6468
rect 48972 6402 49028 6412
rect 49196 6356 49252 6366
rect 48972 6244 49028 6254
rect 48972 5906 49028 6188
rect 48972 5854 48974 5906
rect 49026 5854 49028 5906
rect 48972 5842 49028 5854
rect 48748 5234 48916 5236
rect 48748 5182 48750 5234
rect 48802 5182 48916 5234
rect 48748 5180 48916 5182
rect 48748 5170 48804 5180
rect 49196 5124 49252 6300
rect 48972 5122 49252 5124
rect 48972 5070 49198 5122
rect 49250 5070 49252 5122
rect 48972 5068 49252 5070
rect 48748 4788 48804 4798
rect 48748 4562 48804 4732
rect 48748 4510 48750 4562
rect 48802 4510 48804 4562
rect 48748 4498 48804 4510
rect 48636 3714 48692 3724
rect 48748 3668 48804 3678
rect 48748 3574 48804 3612
rect 48076 3332 48132 3342
rect 48076 3238 48132 3276
rect 48972 2772 49028 5068
rect 49196 5058 49252 5068
rect 49308 6132 49364 6142
rect 49308 4900 49364 6076
rect 49084 4844 49364 4900
rect 49084 4562 49140 4844
rect 49084 4510 49086 4562
rect 49138 4510 49140 4562
rect 49084 4498 49140 4510
rect 49196 4676 49252 4686
rect 48972 2706 49028 2716
rect 49196 3554 49252 4620
rect 49196 3502 49198 3554
rect 49250 3502 49252 3554
rect 49196 2324 49252 3502
rect 49196 2258 49252 2268
rect 49532 800 49588 10220
rect 21196 700 21588 756
rect 22624 0 22736 800
rect 24416 0 24528 800
rect 26208 0 26320 800
rect 28000 0 28112 800
rect 29792 0 29904 800
rect 31584 0 31696 800
rect 33376 0 33488 800
rect 35168 0 35280 800
rect 36960 0 37072 800
rect 38752 0 38864 800
rect 40544 0 40656 800
rect 42336 0 42448 800
rect 44128 0 44240 800
rect 45920 0 46032 800
rect 47712 0 47824 800
rect 49504 0 49616 800
<< via2 >>
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 48188 48860 48244 48916
rect 33740 47964 33796 48020
rect 6300 46844 6356 46900
rect 15820 47292 15876 47348
rect 11900 46844 11956 46900
rect 6636 46732 6692 46788
rect 8428 46786 8484 46788
rect 8428 46734 8430 46786
rect 8430 46734 8482 46786
rect 8482 46734 8484 46786
rect 8428 46732 8484 46734
rect 3388 46562 3444 46564
rect 3388 46510 3390 46562
rect 3390 46510 3442 46562
rect 3442 46510 3444 46562
rect 3388 46508 3444 46510
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 3052 45724 3108 45780
rect 4396 45778 4452 45780
rect 4396 45726 4398 45778
rect 4398 45726 4450 45778
rect 4450 45726 4452 45778
rect 4396 45724 4452 45726
rect 3500 43596 3556 43652
rect 3052 43538 3108 43540
rect 3052 43486 3054 43538
rect 3054 43486 3106 43538
rect 3106 43486 3108 43538
rect 3052 43484 3108 43486
rect 3948 43484 4004 43540
rect 3276 43426 3332 43428
rect 3276 43374 3278 43426
rect 3278 43374 3330 43426
rect 3330 43374 3332 43426
rect 3276 43372 3332 43374
rect 2492 43260 2548 43316
rect 3836 43314 3892 43316
rect 3836 43262 3838 43314
rect 3838 43262 3890 43314
rect 3890 43262 3892 43314
rect 3836 43260 3892 43262
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4620 44268 4676 44324
rect 9548 46732 9604 46788
rect 7084 46508 7140 46564
rect 4956 45724 5012 45780
rect 5180 44994 5236 44996
rect 5180 44942 5182 44994
rect 5182 44942 5234 44994
rect 5234 44942 5236 44994
rect 5180 44940 5236 44942
rect 5852 44940 5908 44996
rect 6300 45836 6356 45892
rect 6076 45666 6132 45668
rect 6076 45614 6078 45666
rect 6078 45614 6130 45666
rect 6130 45614 6132 45666
rect 6076 45612 6132 45614
rect 5740 44322 5796 44324
rect 5740 44270 5742 44322
rect 5742 44270 5794 44322
rect 5794 44270 5796 44322
rect 5740 44268 5796 44270
rect 6748 44940 6804 44996
rect 5852 43932 5908 43988
rect 5740 43708 5796 43764
rect 4844 43596 4900 43652
rect 5628 43650 5684 43652
rect 5628 43598 5630 43650
rect 5630 43598 5682 43650
rect 5682 43598 5684 43650
rect 5628 43596 5684 43598
rect 2940 40348 2996 40404
rect 3724 40402 3780 40404
rect 3724 40350 3726 40402
rect 3726 40350 3778 40402
rect 3778 40350 3780 40402
rect 3724 40348 3780 40350
rect 2940 39340 2996 39396
rect 2940 38668 2996 38724
rect 4172 43314 4228 43316
rect 4172 43262 4174 43314
rect 4174 43262 4226 43314
rect 4226 43262 4228 43314
rect 4172 43260 4228 43262
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4956 43148 5012 43204
rect 6188 43932 6244 43988
rect 6076 43820 6132 43876
rect 6412 43932 6468 43988
rect 7308 46562 7364 46564
rect 7308 46510 7310 46562
rect 7310 46510 7362 46562
rect 7362 46510 7364 46562
rect 7308 46508 7364 46510
rect 7196 45778 7252 45780
rect 7196 45726 7198 45778
rect 7198 45726 7250 45778
rect 7250 45726 7252 45778
rect 7196 45724 7252 45726
rect 8092 46508 8148 46564
rect 7308 45612 7364 45668
rect 7756 45890 7812 45892
rect 7756 45838 7758 45890
rect 7758 45838 7810 45890
rect 7810 45838 7812 45890
rect 7756 45836 7812 45838
rect 7084 43932 7140 43988
rect 7196 45052 7252 45108
rect 5292 43148 5348 43204
rect 6300 43036 6356 43092
rect 5068 42812 5124 42868
rect 6076 42866 6132 42868
rect 6076 42814 6078 42866
rect 6078 42814 6130 42866
rect 6130 42814 6132 42866
rect 6076 42812 6132 42814
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4508 40460 4564 40516
rect 6412 42978 6468 42980
rect 6412 42926 6414 42978
rect 6414 42926 6466 42978
rect 6466 42926 6468 42978
rect 6412 42924 6468 42926
rect 7084 43484 7140 43540
rect 6860 42924 6916 42980
rect 7756 45052 7812 45108
rect 8988 45106 9044 45108
rect 8988 45054 8990 45106
rect 8990 45054 9042 45106
rect 9042 45054 9044 45106
rect 8988 45052 9044 45054
rect 7644 43762 7700 43764
rect 7644 43710 7646 43762
rect 7646 43710 7698 43762
rect 7698 43710 7700 43762
rect 7644 43708 7700 43710
rect 7420 43650 7476 43652
rect 7420 43598 7422 43650
rect 7422 43598 7474 43650
rect 7474 43598 7476 43650
rect 7420 43596 7476 43598
rect 7532 43426 7588 43428
rect 7532 43374 7534 43426
rect 7534 43374 7586 43426
rect 7586 43374 7588 43426
rect 7532 43372 7588 43374
rect 8092 43314 8148 43316
rect 8092 43262 8094 43314
rect 8094 43262 8146 43314
rect 8146 43262 8148 43314
rect 8092 43260 8148 43262
rect 8540 43484 8596 43540
rect 8876 43484 8932 43540
rect 8204 43148 8260 43204
rect 8428 43314 8484 43316
rect 8428 43262 8430 43314
rect 8430 43262 8482 43314
rect 8482 43262 8484 43314
rect 8428 43260 8484 43262
rect 8428 42812 8484 42868
rect 8876 42700 8932 42756
rect 6636 41970 6692 41972
rect 6636 41918 6638 41970
rect 6638 41918 6690 41970
rect 6690 41918 6692 41970
rect 6636 41916 6692 41918
rect 8204 42588 8260 42644
rect 7980 42194 8036 42196
rect 7980 42142 7982 42194
rect 7982 42142 8034 42194
rect 8034 42142 8036 42194
rect 7980 42140 8036 42142
rect 8316 42140 8372 42196
rect 4620 40402 4676 40404
rect 4620 40350 4622 40402
rect 4622 40350 4674 40402
rect 4674 40350 4676 40402
rect 4620 40348 4676 40350
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 9772 43426 9828 43428
rect 9772 43374 9774 43426
rect 9774 43374 9826 43426
rect 9826 43374 9828 43426
rect 9772 43372 9828 43374
rect 10444 43538 10500 43540
rect 10444 43486 10446 43538
rect 10446 43486 10498 43538
rect 10498 43486 10500 43538
rect 10444 43484 10500 43486
rect 11228 43538 11284 43540
rect 11228 43486 11230 43538
rect 11230 43486 11282 43538
rect 11282 43486 11284 43538
rect 11228 43484 11284 43486
rect 10780 43372 10836 43428
rect 10444 43260 10500 43316
rect 9884 42866 9940 42868
rect 9884 42814 9886 42866
rect 9886 42814 9938 42866
rect 9938 42814 9940 42866
rect 9884 42812 9940 42814
rect 10332 42754 10388 42756
rect 10332 42702 10334 42754
rect 10334 42702 10386 42754
rect 10386 42702 10388 42754
rect 10332 42700 10388 42702
rect 10220 42642 10276 42644
rect 10220 42590 10222 42642
rect 10222 42590 10274 42642
rect 10274 42590 10276 42642
rect 10220 42588 10276 42590
rect 9660 42140 9716 42196
rect 8652 41970 8708 41972
rect 8652 41918 8654 41970
rect 8654 41918 8706 41970
rect 8706 41918 8708 41970
rect 8652 41916 8708 41918
rect 6188 40572 6244 40628
rect 5068 40460 5124 40516
rect 5404 40460 5460 40516
rect 5068 40012 5124 40068
rect 6076 40012 6132 40068
rect 4956 39564 5012 39620
rect 6300 40402 6356 40404
rect 6300 40350 6302 40402
rect 6302 40350 6354 40402
rect 6354 40350 6356 40402
rect 6300 40348 6356 40350
rect 6748 40012 6804 40068
rect 5852 39452 5908 39508
rect 5740 39394 5796 39396
rect 5740 39342 5742 39394
rect 5742 39342 5794 39394
rect 5794 39342 5796 39394
rect 5740 39340 5796 39342
rect 5292 38722 5348 38724
rect 5292 38670 5294 38722
rect 5294 38670 5346 38722
rect 5346 38670 5348 38722
rect 5292 38668 5348 38670
rect 5964 38892 6020 38948
rect 2716 37996 2772 38052
rect 2268 36652 2324 36708
rect 2828 36652 2884 36708
rect 1932 35196 1988 35252
rect 2268 34690 2324 34692
rect 2268 34638 2270 34690
rect 2270 34638 2322 34690
rect 2322 34638 2324 34690
rect 2268 34636 2324 34638
rect 2268 34300 2324 34356
rect 2044 34130 2100 34132
rect 2044 34078 2046 34130
rect 2046 34078 2098 34130
rect 2098 34078 2100 34130
rect 2044 34076 2100 34078
rect 1932 32396 1988 32452
rect 1820 31948 1876 32004
rect 2492 35084 2548 35140
rect 2716 34748 2772 34804
rect 2716 34300 2772 34356
rect 3052 35196 3108 35252
rect 3164 35026 3220 35028
rect 3164 34974 3166 35026
rect 3166 34974 3218 35026
rect 3218 34974 3220 35026
rect 3164 34972 3220 34974
rect 2940 34636 2996 34692
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 5628 37996 5684 38052
rect 3500 35196 3556 35252
rect 3612 35026 3668 35028
rect 3612 34974 3614 35026
rect 3614 34974 3666 35026
rect 3666 34974 3668 35026
rect 3612 34972 3668 34974
rect 3388 34860 3444 34916
rect 3836 34748 3892 34804
rect 3724 34690 3780 34692
rect 3724 34638 3726 34690
rect 3726 34638 3778 34690
rect 3778 34638 3780 34690
rect 3724 34636 3780 34638
rect 4956 37266 5012 37268
rect 4956 37214 4958 37266
rect 4958 37214 5010 37266
rect 5010 37214 5012 37266
rect 4956 37212 5012 37214
rect 7756 40572 7812 40628
rect 7644 40460 7700 40516
rect 7532 39618 7588 39620
rect 7532 39566 7534 39618
rect 7534 39566 7586 39618
rect 7586 39566 7588 39618
rect 7532 39564 7588 39566
rect 8316 40572 8372 40628
rect 7756 39618 7812 39620
rect 7756 39566 7758 39618
rect 7758 39566 7810 39618
rect 7810 39566 7812 39618
rect 7756 39564 7812 39566
rect 6972 38780 7028 38836
rect 7084 38892 7140 38948
rect 8204 40460 8260 40516
rect 8092 39452 8148 39508
rect 8540 39676 8596 39732
rect 8540 39506 8596 39508
rect 8540 39454 8542 39506
rect 8542 39454 8594 39506
rect 8594 39454 8596 39506
rect 8540 39452 8596 39454
rect 6412 37378 6468 37380
rect 6412 37326 6414 37378
rect 6414 37326 6466 37378
rect 6466 37326 6468 37378
rect 6412 37324 6468 37326
rect 8876 40178 8932 40180
rect 8876 40126 8878 40178
rect 8878 40126 8930 40178
rect 8930 40126 8932 40178
rect 8876 40124 8932 40126
rect 8988 39004 9044 39060
rect 9996 41132 10052 41188
rect 9548 40460 9604 40516
rect 9884 41020 9940 41076
rect 9436 40124 9492 40180
rect 9324 39564 9380 39620
rect 9548 38834 9604 38836
rect 9548 38782 9550 38834
rect 9550 38782 9602 38834
rect 9602 38782 9604 38834
rect 9548 38780 9604 38782
rect 9884 39004 9940 39060
rect 10220 39452 10276 39508
rect 6076 37266 6132 37268
rect 6076 37214 6078 37266
rect 6078 37214 6130 37266
rect 6130 37214 6132 37266
rect 6076 37212 6132 37214
rect 4060 34412 4116 34468
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4620 36594 4676 36596
rect 4620 36542 4622 36594
rect 4622 36542 4674 36594
rect 4674 36542 4676 36594
rect 4620 36540 4676 36542
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 3164 34076 3220 34132
rect 2940 33852 2996 33908
rect 2156 31948 2212 32004
rect 4732 34636 4788 34692
rect 4508 34300 4564 34356
rect 4284 33852 4340 33908
rect 4844 34524 4900 34580
rect 5068 35026 5124 35028
rect 5068 34974 5070 35026
rect 5070 34974 5122 35026
rect 5122 34974 5124 35026
rect 5068 34972 5124 34974
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5068 33458 5124 33460
rect 5068 33406 5070 33458
rect 5070 33406 5122 33458
rect 5122 33406 5124 33458
rect 5068 33404 5124 33406
rect 3052 32450 3108 32452
rect 3052 32398 3054 32450
rect 3054 32398 3106 32450
rect 3106 32398 3108 32450
rect 3052 32396 3108 32398
rect 2268 31836 2324 31892
rect 2604 30994 2660 30996
rect 2604 30942 2606 30994
rect 2606 30942 2658 30994
rect 2658 30942 2660 30994
rect 2604 30940 2660 30942
rect 3500 30994 3556 30996
rect 3500 30942 3502 30994
rect 3502 30942 3554 30994
rect 3554 30942 3556 30994
rect 3500 30940 3556 30942
rect 3052 30380 3108 30436
rect 3276 28700 3332 28756
rect 2604 28588 2660 28644
rect 2492 26908 2548 26964
rect 3388 28642 3444 28644
rect 3388 28590 3390 28642
rect 3390 28590 3442 28642
rect 3442 28590 3444 28642
rect 3388 28588 3444 28590
rect 3612 28588 3668 28644
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4620 31890 4676 31892
rect 4620 31838 4622 31890
rect 4622 31838 4674 31890
rect 4674 31838 4676 31890
rect 4620 31836 4676 31838
rect 4956 31836 5012 31892
rect 4060 30994 4116 30996
rect 4060 30942 4062 30994
rect 4062 30942 4114 30994
rect 4114 30942 4116 30994
rect 4060 30940 4116 30942
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4956 30044 5012 30100
rect 6524 36988 6580 37044
rect 6300 35532 6356 35588
rect 7420 35698 7476 35700
rect 7420 35646 7422 35698
rect 7422 35646 7474 35698
rect 7474 35646 7476 35698
rect 7420 35644 7476 35646
rect 6636 35532 6692 35588
rect 7196 35586 7252 35588
rect 7196 35534 7198 35586
rect 7198 35534 7250 35586
rect 7250 35534 7252 35586
rect 7196 35532 7252 35534
rect 6188 34972 6244 35028
rect 5628 34914 5684 34916
rect 5628 34862 5630 34914
rect 5630 34862 5682 34914
rect 5682 34862 5684 34914
rect 5628 34860 5684 34862
rect 5740 34748 5796 34804
rect 5852 34636 5908 34692
rect 7308 34972 7364 35028
rect 6300 34300 6356 34356
rect 8764 38610 8820 38612
rect 8764 38558 8766 38610
rect 8766 38558 8818 38610
rect 8818 38558 8820 38610
rect 8764 38556 8820 38558
rect 8540 37324 8596 37380
rect 10780 42754 10836 42756
rect 10780 42702 10782 42754
rect 10782 42702 10834 42754
rect 10834 42702 10836 42754
rect 10780 42700 10836 42702
rect 10556 40908 10612 40964
rect 11564 42978 11620 42980
rect 11564 42926 11566 42978
rect 11566 42926 11618 42978
rect 11618 42926 11620 42978
rect 11564 42924 11620 42926
rect 11452 42700 11508 42756
rect 11676 41074 11732 41076
rect 11676 41022 11678 41074
rect 11678 41022 11730 41074
rect 11730 41022 11732 41074
rect 11676 41020 11732 41022
rect 11452 39506 11508 39508
rect 11452 39454 11454 39506
rect 11454 39454 11506 39506
rect 11506 39454 11508 39506
rect 11452 39452 11508 39454
rect 12012 43484 12068 43540
rect 12124 42754 12180 42756
rect 12124 42702 12126 42754
rect 12126 42702 12178 42754
rect 12178 42702 12180 42754
rect 12124 42700 12180 42702
rect 12684 41916 12740 41972
rect 12460 41186 12516 41188
rect 12460 41134 12462 41186
rect 12462 41134 12514 41186
rect 12514 41134 12516 41186
rect 12460 41132 12516 41134
rect 12796 40962 12852 40964
rect 12796 40910 12798 40962
rect 12798 40910 12850 40962
rect 12850 40910 12852 40962
rect 12796 40908 12852 40910
rect 15148 42642 15204 42644
rect 15148 42590 15150 42642
rect 15150 42590 15202 42642
rect 15202 42590 15204 42642
rect 15148 42588 15204 42590
rect 13580 41186 13636 41188
rect 13580 41134 13582 41186
rect 13582 41134 13634 41186
rect 13634 41134 13636 41186
rect 13580 41132 13636 41134
rect 8316 37042 8372 37044
rect 8316 36990 8318 37042
rect 8318 36990 8370 37042
rect 8370 36990 8372 37042
rect 8316 36988 8372 36990
rect 8092 36540 8148 36596
rect 9996 38610 10052 38612
rect 9996 38558 9998 38610
rect 9998 38558 10050 38610
rect 10050 38558 10052 38610
rect 9996 38556 10052 38558
rect 10556 38050 10612 38052
rect 10556 37998 10558 38050
rect 10558 37998 10610 38050
rect 10610 37998 10612 38050
rect 10556 37996 10612 37998
rect 10780 37826 10836 37828
rect 10780 37774 10782 37826
rect 10782 37774 10834 37826
rect 10834 37774 10836 37826
rect 10780 37772 10836 37774
rect 8316 35698 8372 35700
rect 8316 35646 8318 35698
rect 8318 35646 8370 35698
rect 8370 35646 8372 35698
rect 8316 35644 8372 35646
rect 8652 35698 8708 35700
rect 8652 35646 8654 35698
rect 8654 35646 8706 35698
rect 8706 35646 8708 35698
rect 8652 35644 8708 35646
rect 7980 35084 8036 35140
rect 8540 35026 8596 35028
rect 8540 34974 8542 35026
rect 8542 34974 8594 35026
rect 8594 34974 8596 35026
rect 8540 34972 8596 34974
rect 7868 34300 7924 34356
rect 5964 33404 6020 33460
rect 5516 31948 5572 32004
rect 5628 31836 5684 31892
rect 5964 31948 6020 32004
rect 5292 30044 5348 30100
rect 4620 29426 4676 29428
rect 4620 29374 4622 29426
rect 4622 29374 4674 29426
rect 4674 29374 4676 29426
rect 4620 29372 4676 29374
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 3724 28476 3780 28532
rect 4732 28812 4788 28868
rect 3276 27244 3332 27300
rect 4396 28700 4452 28756
rect 3836 27244 3892 27300
rect 4508 28642 4564 28644
rect 4508 28590 4510 28642
rect 4510 28590 4562 28642
rect 4562 28590 4564 28642
rect 4508 28588 4564 28590
rect 6300 31106 6356 31108
rect 6300 31054 6302 31106
rect 6302 31054 6354 31106
rect 6354 31054 6356 31106
rect 6300 31052 6356 31054
rect 5964 30716 6020 30772
rect 5292 28588 5348 28644
rect 5516 29426 5572 29428
rect 5516 29374 5518 29426
rect 5518 29374 5570 29426
rect 5570 29374 5572 29426
rect 5516 29372 5572 29374
rect 4844 28476 4900 28532
rect 3612 26962 3668 26964
rect 3612 26910 3614 26962
rect 3614 26910 3666 26962
rect 3666 26910 3668 26962
rect 3612 26908 3668 26910
rect 1820 26290 1876 26292
rect 1820 26238 1822 26290
rect 1822 26238 1874 26290
rect 1874 26238 1876 26290
rect 1820 26236 1876 26238
rect 4620 27804 4676 27860
rect 5628 28812 5684 28868
rect 6972 32956 7028 33012
rect 6412 30716 6468 30772
rect 6412 28754 6468 28756
rect 6412 28702 6414 28754
rect 6414 28702 6466 28754
rect 6466 28702 6468 28754
rect 6412 28700 6468 28702
rect 5964 28588 6020 28644
rect 5516 27858 5572 27860
rect 5516 27806 5518 27858
rect 5518 27806 5570 27858
rect 5570 27806 5572 27858
rect 5516 27804 5572 27806
rect 6860 30882 6916 30884
rect 6860 30830 6862 30882
rect 6862 30830 6914 30882
rect 6914 30830 6916 30882
rect 6860 30828 6916 30830
rect 7308 33180 7364 33236
rect 7196 30770 7252 30772
rect 7196 30718 7198 30770
rect 7198 30718 7250 30770
rect 7250 30718 7252 30770
rect 7196 30716 7252 30718
rect 7196 30492 7252 30548
rect 7756 33234 7812 33236
rect 7756 33182 7758 33234
rect 7758 33182 7810 33234
rect 7810 33182 7812 33234
rect 7756 33180 7812 33182
rect 9212 36482 9268 36484
rect 9212 36430 9214 36482
rect 9214 36430 9266 36482
rect 9266 36430 9268 36482
rect 9212 36428 9268 36430
rect 11788 37772 11844 37828
rect 10220 36594 10276 36596
rect 10220 36542 10222 36594
rect 10222 36542 10274 36594
rect 10274 36542 10276 36594
rect 10220 36540 10276 36542
rect 11228 36540 11284 36596
rect 8876 36316 8932 36372
rect 9660 36316 9716 36372
rect 9212 36204 9268 36260
rect 8988 35196 9044 35252
rect 9324 35138 9380 35140
rect 9324 35086 9326 35138
rect 9326 35086 9378 35138
rect 9378 35086 9380 35138
rect 9324 35084 9380 35086
rect 9324 34690 9380 34692
rect 9324 34638 9326 34690
rect 9326 34638 9378 34690
rect 9378 34638 9380 34690
rect 9324 34636 9380 34638
rect 9884 36428 9940 36484
rect 9660 35644 9716 35700
rect 10556 36482 10612 36484
rect 10556 36430 10558 36482
rect 10558 36430 10610 36482
rect 10610 36430 10612 36482
rect 10556 36428 10612 36430
rect 11564 36482 11620 36484
rect 11564 36430 11566 36482
rect 11566 36430 11618 36482
rect 11618 36430 11620 36482
rect 11564 36428 11620 36430
rect 11452 36258 11508 36260
rect 11452 36206 11454 36258
rect 11454 36206 11506 36258
rect 11506 36206 11508 36258
rect 11452 36204 11508 36206
rect 9772 35084 9828 35140
rect 7532 30882 7588 30884
rect 7532 30830 7534 30882
rect 7534 30830 7586 30882
rect 7586 30830 7588 30882
rect 7532 30828 7588 30830
rect 8316 33180 8372 33236
rect 9100 33346 9156 33348
rect 9100 33294 9102 33346
rect 9102 33294 9154 33346
rect 9154 33294 9156 33346
rect 9100 33292 9156 33294
rect 8876 33068 8932 33124
rect 8764 31948 8820 32004
rect 9212 31724 9268 31780
rect 9436 33234 9492 33236
rect 9436 33182 9438 33234
rect 9438 33182 9490 33234
rect 9490 33182 9492 33234
rect 9436 33180 9492 33182
rect 10444 35196 10500 35252
rect 10108 34354 10164 34356
rect 10108 34302 10110 34354
rect 10110 34302 10162 34354
rect 10162 34302 10164 34354
rect 10108 34300 10164 34302
rect 14028 39618 14084 39620
rect 14028 39566 14030 39618
rect 14030 39566 14082 39618
rect 14082 39566 14084 39618
rect 14028 39564 14084 39566
rect 13916 38668 13972 38724
rect 12684 38220 12740 38276
rect 13580 38274 13636 38276
rect 13580 38222 13582 38274
rect 13582 38222 13634 38274
rect 13634 38222 13636 38274
rect 13580 38220 13636 38222
rect 15036 39618 15092 39620
rect 15036 39566 15038 39618
rect 15038 39566 15090 39618
rect 15090 39566 15092 39618
rect 15036 39564 15092 39566
rect 14924 39506 14980 39508
rect 14924 39454 14926 39506
rect 14926 39454 14978 39506
rect 14978 39454 14980 39506
rect 14924 39452 14980 39454
rect 12684 36316 12740 36372
rect 13804 36370 13860 36372
rect 13804 36318 13806 36370
rect 13806 36318 13858 36370
rect 13858 36318 13860 36370
rect 13804 36316 13860 36318
rect 11788 35196 11844 35252
rect 12684 35196 12740 35252
rect 10556 34636 10612 34692
rect 11228 33964 11284 34020
rect 11004 33292 11060 33348
rect 10556 33234 10612 33236
rect 10556 33182 10558 33234
rect 10558 33182 10610 33234
rect 10610 33182 10612 33234
rect 10556 33180 10612 33182
rect 10892 33068 10948 33124
rect 10108 32674 10164 32676
rect 10108 32622 10110 32674
rect 10110 32622 10162 32674
rect 10162 32622 10164 32674
rect 10108 32620 10164 32622
rect 10780 32620 10836 32676
rect 9772 32562 9828 32564
rect 9772 32510 9774 32562
rect 9774 32510 9826 32562
rect 9826 32510 9828 32562
rect 9772 32508 9828 32510
rect 9324 31612 9380 31668
rect 9884 31948 9940 32004
rect 9772 31890 9828 31892
rect 9772 31838 9774 31890
rect 9774 31838 9826 31890
rect 9826 31838 9828 31890
rect 9772 31836 9828 31838
rect 8316 31164 8372 31220
rect 8204 31106 8260 31108
rect 8204 31054 8206 31106
rect 8206 31054 8258 31106
rect 8258 31054 8260 31106
rect 8204 31052 8260 31054
rect 8652 31106 8708 31108
rect 8652 31054 8654 31106
rect 8654 31054 8706 31106
rect 8706 31054 8708 31106
rect 8652 31052 8708 31054
rect 9212 31052 9268 31108
rect 8316 30492 8372 30548
rect 7868 30380 7924 30436
rect 8316 30268 8372 30324
rect 6636 29372 6692 29428
rect 7308 29426 7364 29428
rect 7308 29374 7310 29426
rect 7310 29374 7362 29426
rect 7362 29374 7364 29426
rect 7308 29372 7364 29374
rect 6636 28588 6692 28644
rect 5852 27804 5908 27860
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4508 27298 4564 27300
rect 4508 27246 4510 27298
rect 4510 27246 4562 27298
rect 4562 27246 4564 27298
rect 4508 27244 4564 27246
rect 5068 27244 5124 27300
rect 4844 27074 4900 27076
rect 4844 27022 4846 27074
rect 4846 27022 4898 27074
rect 4898 27022 4900 27074
rect 4844 27020 4900 27022
rect 3948 26796 4004 26852
rect 5292 27020 5348 27076
rect 5068 26796 5124 26852
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4844 25788 4900 25844
rect 4172 25730 4228 25732
rect 4172 25678 4174 25730
rect 4174 25678 4226 25730
rect 4226 25678 4228 25730
rect 4172 25676 4228 25678
rect 5292 25676 5348 25732
rect 3724 25564 3780 25620
rect 2492 24610 2548 24612
rect 2492 24558 2494 24610
rect 2494 24558 2546 24610
rect 2546 24558 2548 24610
rect 2492 24556 2548 24558
rect 6524 27692 6580 27748
rect 5964 27244 6020 27300
rect 6076 27580 6132 27636
rect 6412 27298 6468 27300
rect 6412 27246 6414 27298
rect 6414 27246 6466 27298
rect 6466 27246 6468 27298
rect 6412 27244 6468 27246
rect 7084 28364 7140 28420
rect 7420 27804 7476 27860
rect 7084 27244 7140 27300
rect 6188 26290 6244 26292
rect 6188 26238 6190 26290
rect 6190 26238 6242 26290
rect 6242 26238 6244 26290
rect 6188 26236 6244 26238
rect 6076 25788 6132 25844
rect 7980 29426 8036 29428
rect 7980 29374 7982 29426
rect 7982 29374 8034 29426
rect 8034 29374 8036 29426
rect 7980 29372 8036 29374
rect 7756 28476 7812 28532
rect 7868 27746 7924 27748
rect 7868 27694 7870 27746
rect 7870 27694 7922 27746
rect 7922 27694 7924 27746
rect 7868 27692 7924 27694
rect 7196 25730 7252 25732
rect 7196 25678 7198 25730
rect 7198 25678 7250 25730
rect 7250 25678 7252 25730
rect 7196 25676 7252 25678
rect 3948 25116 4004 25172
rect 4620 24444 4676 24500
rect 5068 25116 5124 25172
rect 6300 25564 6356 25620
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 2492 23324 2548 23380
rect 4284 23324 4340 23380
rect 3388 23266 3444 23268
rect 3388 23214 3390 23266
rect 3390 23214 3442 23266
rect 3442 23214 3444 23266
rect 3388 23212 3444 23214
rect 2828 22988 2884 23044
rect 3500 23042 3556 23044
rect 3500 22990 3502 23042
rect 3502 22990 3554 23042
rect 3554 22990 3556 23042
rect 3500 22988 3556 22990
rect 4060 23154 4116 23156
rect 4060 23102 4062 23154
rect 4062 23102 4114 23154
rect 4114 23102 4116 23154
rect 4060 23100 4116 23102
rect 4620 24108 4676 24164
rect 5180 24444 5236 24500
rect 5180 23884 5236 23940
rect 4844 23772 4900 23828
rect 6860 25618 6916 25620
rect 6860 25566 6862 25618
rect 6862 25566 6914 25618
rect 6914 25566 6916 25618
rect 6860 25564 6916 25566
rect 7644 25564 7700 25620
rect 7084 25506 7140 25508
rect 7084 25454 7086 25506
rect 7086 25454 7138 25506
rect 7138 25454 7140 25506
rect 7084 25452 7140 25454
rect 6412 25394 6468 25396
rect 6412 25342 6414 25394
rect 6414 25342 6466 25394
rect 6466 25342 6468 25394
rect 6412 25340 6468 25342
rect 8764 28588 8820 28644
rect 9548 31218 9604 31220
rect 9548 31166 9550 31218
rect 9550 31166 9602 31218
rect 9602 31166 9604 31218
rect 9548 31164 9604 31166
rect 9996 31612 10052 31668
rect 9996 30268 10052 30324
rect 10780 31836 10836 31892
rect 12124 34018 12180 34020
rect 12124 33966 12126 34018
rect 12126 33966 12178 34018
rect 12178 33966 12180 34018
rect 12124 33964 12180 33966
rect 12684 33964 12740 34020
rect 11564 33068 11620 33124
rect 11228 32620 11284 32676
rect 11116 32562 11172 32564
rect 11116 32510 11118 32562
rect 11118 32510 11170 32562
rect 11170 32510 11172 32562
rect 11116 32508 11172 32510
rect 11676 32508 11732 32564
rect 12572 33292 12628 33348
rect 12572 31724 12628 31780
rect 10668 31164 10724 31220
rect 10444 31052 10500 31108
rect 12124 30940 12180 30996
rect 10220 30492 10276 30548
rect 8988 28364 9044 28420
rect 8988 27692 9044 27748
rect 8540 27634 8596 27636
rect 8540 27582 8542 27634
rect 8542 27582 8594 27634
rect 8594 27582 8596 27634
rect 8540 27580 8596 27582
rect 8428 26236 8484 26292
rect 12124 29314 12180 29316
rect 12124 29262 12126 29314
rect 12126 29262 12178 29314
rect 12178 29262 12180 29314
rect 12124 29260 12180 29262
rect 12348 28028 12404 28084
rect 11452 27746 11508 27748
rect 11452 27694 11454 27746
rect 11454 27694 11506 27746
rect 11506 27694 11508 27746
rect 11452 27692 11508 27694
rect 12012 27746 12068 27748
rect 12012 27694 12014 27746
rect 12014 27694 12066 27746
rect 12066 27694 12068 27746
rect 12012 27692 12068 27694
rect 12572 27356 12628 27412
rect 12796 27746 12852 27748
rect 12796 27694 12798 27746
rect 12798 27694 12850 27746
rect 12850 27694 12852 27746
rect 12796 27692 12852 27694
rect 13692 36204 13748 36260
rect 15484 39340 15540 39396
rect 15484 38556 15540 38612
rect 15148 38050 15204 38052
rect 15148 37998 15150 38050
rect 15150 37998 15202 38050
rect 15202 37998 15204 38050
rect 15148 37996 15204 37998
rect 15036 37826 15092 37828
rect 15036 37774 15038 37826
rect 15038 37774 15090 37826
rect 15090 37774 15092 37826
rect 15036 37772 15092 37774
rect 15372 37660 15428 37716
rect 15708 38722 15764 38724
rect 15708 38670 15710 38722
rect 15710 38670 15762 38722
rect 15762 38670 15764 38722
rect 15708 38668 15764 38670
rect 19852 47346 19908 47348
rect 19852 47294 19854 47346
rect 19854 47294 19906 47346
rect 19906 47294 19908 47346
rect 19852 47292 19908 47294
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 18396 45164 18452 45220
rect 16492 44322 16548 44324
rect 16492 44270 16494 44322
rect 16494 44270 16546 44322
rect 16546 44270 16548 44322
rect 16492 44268 16548 44270
rect 18396 44268 18452 44324
rect 16492 42642 16548 42644
rect 16492 42590 16494 42642
rect 16494 42590 16546 42642
rect 16546 42590 16548 42642
rect 16492 42588 16548 42590
rect 16380 41804 16436 41860
rect 16380 41298 16436 41300
rect 16380 41246 16382 41298
rect 16382 41246 16434 41298
rect 16434 41246 16436 41298
rect 16380 41244 16436 41246
rect 16156 40236 16212 40292
rect 16940 41804 16996 41860
rect 18508 44380 18564 44436
rect 18284 42530 18340 42532
rect 18284 42478 18286 42530
rect 18286 42478 18338 42530
rect 18338 42478 18340 42530
rect 18284 42476 18340 42478
rect 18620 42476 18676 42532
rect 21644 45218 21700 45220
rect 21644 45166 21646 45218
rect 21646 45166 21698 45218
rect 21698 45166 21700 45218
rect 21644 45164 21700 45166
rect 23884 46620 23940 46676
rect 21980 44380 22036 44436
rect 20300 44210 20356 44212
rect 20300 44158 20302 44210
rect 20302 44158 20354 44210
rect 20354 44158 20356 44210
rect 20300 44156 20356 44158
rect 22316 44210 22372 44212
rect 22316 44158 22318 44210
rect 22318 44158 22370 44210
rect 22370 44158 22372 44210
rect 22316 44156 22372 44158
rect 21644 44098 21700 44100
rect 21644 44046 21646 44098
rect 21646 44046 21698 44098
rect 21698 44046 21700 44098
rect 21644 44044 21700 44046
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20188 42924 20244 42980
rect 19180 42866 19236 42868
rect 19180 42814 19182 42866
rect 19182 42814 19234 42866
rect 19234 42814 19236 42866
rect 19180 42812 19236 42814
rect 20076 42642 20132 42644
rect 20076 42590 20078 42642
rect 20078 42590 20130 42642
rect 20130 42590 20132 42642
rect 20076 42588 20132 42590
rect 19068 42530 19124 42532
rect 19068 42478 19070 42530
rect 19070 42478 19122 42530
rect 19122 42478 19124 42530
rect 19068 42476 19124 42478
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 18732 42140 18788 42196
rect 18284 41916 18340 41972
rect 16716 41132 16772 41188
rect 17052 41020 17108 41076
rect 16604 40684 16660 40740
rect 16156 39452 16212 39508
rect 15932 38556 15988 38612
rect 15596 37996 15652 38052
rect 15596 37324 15652 37380
rect 14924 37100 14980 37156
rect 15932 38050 15988 38052
rect 15932 37998 15934 38050
rect 15934 37998 15986 38050
rect 15986 37998 15988 38050
rect 15932 37996 15988 37998
rect 17500 41804 17556 41860
rect 17500 40908 17556 40964
rect 17500 40684 17556 40740
rect 18172 41186 18228 41188
rect 18172 41134 18174 41186
rect 18174 41134 18226 41186
rect 18226 41134 18228 41186
rect 18172 41132 18228 41134
rect 18284 40796 18340 40852
rect 17948 40684 18004 40740
rect 18620 41746 18676 41748
rect 18620 41694 18622 41746
rect 18622 41694 18674 41746
rect 18674 41694 18676 41746
rect 18620 41692 18676 41694
rect 18732 41074 18788 41076
rect 18732 41022 18734 41074
rect 18734 41022 18786 41074
rect 18786 41022 18788 41074
rect 18732 41020 18788 41022
rect 18844 41244 18900 41300
rect 18508 40908 18564 40964
rect 18620 40572 18676 40628
rect 16716 39394 16772 39396
rect 16716 39342 16718 39394
rect 16718 39342 16770 39394
rect 16770 39342 16772 39394
rect 16716 39340 16772 39342
rect 16380 37996 16436 38052
rect 15820 37660 15876 37716
rect 16156 37772 16212 37828
rect 16268 37154 16324 37156
rect 16268 37102 16270 37154
rect 16270 37102 16322 37154
rect 16322 37102 16324 37154
rect 16268 37100 16324 37102
rect 14140 35756 14196 35812
rect 13020 34972 13076 35028
rect 14252 35026 14308 35028
rect 14252 34974 14254 35026
rect 14254 34974 14306 35026
rect 14306 34974 14308 35026
rect 14252 34972 14308 34974
rect 13132 33292 13188 33348
rect 15596 36258 15652 36260
rect 15596 36206 15598 36258
rect 15598 36206 15650 36258
rect 15650 36206 15652 36258
rect 15596 36204 15652 36206
rect 14812 35868 14868 35924
rect 15260 35810 15316 35812
rect 15260 35758 15262 35810
rect 15262 35758 15314 35810
rect 15314 35758 15316 35810
rect 15260 35756 15316 35758
rect 13468 33292 13524 33348
rect 13804 33234 13860 33236
rect 13804 33182 13806 33234
rect 13806 33182 13858 33234
rect 13858 33182 13860 33234
rect 13804 33180 13860 33182
rect 14588 32956 14644 33012
rect 15708 33234 15764 33236
rect 15708 33182 15710 33234
rect 15710 33182 15762 33234
rect 15762 33182 15764 33234
rect 15708 33180 15764 33182
rect 15372 33122 15428 33124
rect 15372 33070 15374 33122
rect 15374 33070 15426 33122
rect 15426 33070 15428 33122
rect 15372 33068 15428 33070
rect 15708 32786 15764 32788
rect 15708 32734 15710 32786
rect 15710 32734 15762 32786
rect 15762 32734 15764 32786
rect 15708 32732 15764 32734
rect 15932 34130 15988 34132
rect 15932 34078 15934 34130
rect 15934 34078 15986 34130
rect 15986 34078 15988 34130
rect 15932 34076 15988 34078
rect 18172 40124 18228 40180
rect 17948 40012 18004 40068
rect 17724 39900 17780 39956
rect 17052 39452 17108 39508
rect 16940 38050 16996 38052
rect 16940 37998 16942 38050
rect 16942 37998 16994 38050
rect 16994 37998 16996 38050
rect 16940 37996 16996 37998
rect 16828 36652 16884 36708
rect 16716 35868 16772 35924
rect 17724 39506 17780 39508
rect 17724 39454 17726 39506
rect 17726 39454 17778 39506
rect 17778 39454 17780 39506
rect 17724 39452 17780 39454
rect 17500 39394 17556 39396
rect 17500 39342 17502 39394
rect 17502 39342 17554 39394
rect 17554 39342 17556 39394
rect 17500 39340 17556 39342
rect 17612 39228 17668 39284
rect 19292 41692 19348 41748
rect 21532 42924 21588 42980
rect 21196 42812 21252 42868
rect 21868 42812 21924 42868
rect 21644 42364 21700 42420
rect 22428 44098 22484 44100
rect 22428 44046 22430 44098
rect 22430 44046 22482 44098
rect 22482 44046 22484 44098
rect 22428 44044 22484 44046
rect 22316 42700 22372 42756
rect 22204 42642 22260 42644
rect 22204 42590 22206 42642
rect 22206 42590 22258 42642
rect 22258 42590 22260 42642
rect 22204 42588 22260 42590
rect 22092 42530 22148 42532
rect 22092 42478 22094 42530
rect 22094 42478 22146 42530
rect 22146 42478 22148 42530
rect 22092 42476 22148 42478
rect 19740 41074 19796 41076
rect 19740 41022 19742 41074
rect 19742 41022 19794 41074
rect 19794 41022 19796 41074
rect 19740 41020 19796 41022
rect 19964 40962 20020 40964
rect 19964 40910 19966 40962
rect 19966 40910 20018 40962
rect 20018 40910 20020 40962
rect 19964 40908 20020 40910
rect 20636 41298 20692 41300
rect 20636 41246 20638 41298
rect 20638 41246 20690 41298
rect 20690 41246 20692 41298
rect 20636 41244 20692 41246
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 18844 40348 18900 40404
rect 20076 40626 20132 40628
rect 20076 40574 20078 40626
rect 20078 40574 20130 40626
rect 20130 40574 20132 40626
rect 20076 40572 20132 40574
rect 20412 40908 20468 40964
rect 19740 40348 19796 40404
rect 18620 39506 18676 39508
rect 18620 39454 18622 39506
rect 18622 39454 18674 39506
rect 18674 39454 18676 39506
rect 18620 39452 18676 39454
rect 19068 39340 19124 39396
rect 17164 38050 17220 38052
rect 17164 37998 17166 38050
rect 17166 37998 17218 38050
rect 17218 37998 17220 38050
rect 17164 37996 17220 37998
rect 17276 37826 17332 37828
rect 17276 37774 17278 37826
rect 17278 37774 17330 37826
rect 17330 37774 17332 37826
rect 17276 37772 17332 37774
rect 18172 38108 18228 38164
rect 17724 37996 17780 38052
rect 17388 37660 17444 37716
rect 17388 37378 17444 37380
rect 17388 37326 17390 37378
rect 17390 37326 17442 37378
rect 17442 37326 17444 37378
rect 17388 37324 17444 37326
rect 17948 37772 18004 37828
rect 18732 38108 18788 38164
rect 18284 37212 18340 37268
rect 18508 37772 18564 37828
rect 18956 37490 19012 37492
rect 18956 37438 18958 37490
rect 18958 37438 19010 37490
rect 19010 37438 19012 37490
rect 18956 37436 19012 37438
rect 19292 37212 19348 37268
rect 17612 36652 17668 36708
rect 17612 35420 17668 35476
rect 17052 35084 17108 35140
rect 16940 34860 16996 34916
rect 18172 35196 18228 35252
rect 18060 35084 18116 35140
rect 17836 34972 17892 35028
rect 20300 40402 20356 40404
rect 20300 40350 20302 40402
rect 20302 40350 20354 40402
rect 20354 40350 20356 40402
rect 20300 40348 20356 40350
rect 19964 40290 20020 40292
rect 19964 40238 19966 40290
rect 19966 40238 20018 40290
rect 20018 40238 20020 40290
rect 19964 40236 20020 40238
rect 20076 39564 20132 39620
rect 20300 39788 20356 39844
rect 20188 39340 20244 39396
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20300 38610 20356 38612
rect 20300 38558 20302 38610
rect 20302 38558 20354 38610
rect 20354 38558 20356 38610
rect 20300 38556 20356 38558
rect 20524 40236 20580 40292
rect 20636 39564 20692 39620
rect 21308 41020 21364 41076
rect 22876 42924 22932 42980
rect 23100 43596 23156 43652
rect 22540 42588 22596 42644
rect 22988 42588 23044 42644
rect 23436 42642 23492 42644
rect 23436 42590 23438 42642
rect 23438 42590 23490 42642
rect 23490 42590 23492 42642
rect 23436 42588 23492 42590
rect 23100 42530 23156 42532
rect 23100 42478 23102 42530
rect 23102 42478 23154 42530
rect 23154 42478 23156 42530
rect 23100 42476 23156 42478
rect 23324 42530 23380 42532
rect 23324 42478 23326 42530
rect 23326 42478 23378 42530
rect 23378 42478 23380 42530
rect 23324 42476 23380 42478
rect 25228 46674 25284 46676
rect 25228 46622 25230 46674
rect 25230 46622 25282 46674
rect 25282 46622 25284 46674
rect 25228 46620 25284 46622
rect 25004 46396 25060 46452
rect 24556 44434 24612 44436
rect 24556 44382 24558 44434
rect 24558 44382 24610 44434
rect 24610 44382 24612 44434
rect 24556 44380 24612 44382
rect 23660 43650 23716 43652
rect 23660 43598 23662 43650
rect 23662 43598 23714 43650
rect 23714 43598 23716 43650
rect 23660 43596 23716 43598
rect 23436 41916 23492 41972
rect 23100 41468 23156 41524
rect 21308 40796 21364 40852
rect 21196 39900 21252 39956
rect 21084 39788 21140 39844
rect 22092 40514 22148 40516
rect 22092 40462 22094 40514
rect 22094 40462 22146 40514
rect 22146 40462 22148 40514
rect 22092 40460 22148 40462
rect 21980 40402 22036 40404
rect 21980 40350 21982 40402
rect 21982 40350 22034 40402
rect 22034 40350 22036 40402
rect 21980 40348 22036 40350
rect 21420 40124 21476 40180
rect 20972 39340 21028 39396
rect 20524 38556 20580 38612
rect 20076 37938 20132 37940
rect 20076 37886 20078 37938
rect 20078 37886 20130 37938
rect 20130 37886 20132 37938
rect 20076 37884 20132 37886
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19628 37436 19684 37492
rect 22428 40460 22484 40516
rect 22204 39900 22260 39956
rect 21756 39506 21812 39508
rect 21756 39454 21758 39506
rect 21758 39454 21810 39506
rect 21810 39454 21812 39506
rect 21756 39452 21812 39454
rect 21532 39394 21588 39396
rect 21532 39342 21534 39394
rect 21534 39342 21586 39394
rect 21586 39342 21588 39394
rect 21532 39340 21588 39342
rect 22652 40796 22708 40852
rect 23548 41692 23604 41748
rect 24556 43372 24612 43428
rect 24108 41804 24164 41860
rect 24108 41186 24164 41188
rect 24108 41134 24110 41186
rect 24110 41134 24162 41186
rect 24162 41134 24164 41186
rect 24108 41132 24164 41134
rect 24780 41186 24836 41188
rect 24780 41134 24782 41186
rect 24782 41134 24834 41186
rect 24834 41134 24836 41186
rect 24780 41132 24836 41134
rect 22652 39340 22708 39396
rect 20972 38108 21028 38164
rect 20524 37212 20580 37268
rect 20076 36988 20132 37044
rect 19516 36204 19572 36260
rect 20524 36540 20580 36596
rect 18844 35196 18900 35252
rect 18172 34860 18228 34916
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20412 35026 20468 35028
rect 20412 34974 20414 35026
rect 20414 34974 20466 35026
rect 20466 34974 20468 35026
rect 20412 34972 20468 34974
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 17724 34188 17780 34244
rect 16380 34076 16436 34132
rect 17388 34130 17444 34132
rect 17388 34078 17390 34130
rect 17390 34078 17442 34130
rect 17442 34078 17444 34130
rect 17388 34076 17444 34078
rect 18620 34018 18676 34020
rect 18620 33966 18622 34018
rect 18622 33966 18674 34018
rect 18674 33966 18676 34018
rect 18620 33964 18676 33966
rect 17164 33570 17220 33572
rect 17164 33518 17166 33570
rect 17166 33518 17218 33570
rect 17218 33518 17220 33570
rect 17164 33516 17220 33518
rect 17500 33292 17556 33348
rect 17836 33516 17892 33572
rect 16156 33234 16212 33236
rect 16156 33182 16158 33234
rect 16158 33182 16210 33234
rect 16210 33182 16212 33234
rect 16156 33180 16212 33182
rect 16380 32956 16436 33012
rect 13580 31778 13636 31780
rect 13580 31726 13582 31778
rect 13582 31726 13634 31778
rect 13634 31726 13636 31778
rect 13580 31724 13636 31726
rect 13020 30994 13076 30996
rect 13020 30942 13022 30994
rect 13022 30942 13074 30994
rect 13074 30942 13076 30994
rect 13020 30940 13076 30942
rect 13804 30716 13860 30772
rect 13916 30268 13972 30324
rect 14476 30492 14532 30548
rect 14476 29260 14532 29316
rect 14028 28700 14084 28756
rect 13468 28028 13524 28084
rect 13132 27692 13188 27748
rect 9212 26236 9268 26292
rect 9548 26290 9604 26292
rect 9548 26238 9550 26290
rect 9550 26238 9602 26290
rect 9602 26238 9604 26290
rect 9548 26236 9604 26238
rect 12460 26236 12516 26292
rect 8428 25506 8484 25508
rect 8428 25454 8430 25506
rect 8430 25454 8482 25506
rect 8482 25454 8484 25506
rect 8428 25452 8484 25454
rect 9772 25506 9828 25508
rect 9772 25454 9774 25506
rect 9774 25454 9826 25506
rect 9826 25454 9828 25506
rect 9772 25452 9828 25454
rect 8316 25394 8372 25396
rect 8316 25342 8318 25394
rect 8318 25342 8370 25394
rect 8370 25342 8372 25394
rect 8316 25340 8372 25342
rect 10444 25506 10500 25508
rect 10444 25454 10446 25506
rect 10446 25454 10498 25506
rect 10498 25454 10500 25506
rect 10444 25452 10500 25454
rect 10780 25506 10836 25508
rect 10780 25454 10782 25506
rect 10782 25454 10834 25506
rect 10834 25454 10836 25506
rect 10780 25452 10836 25454
rect 6188 24610 6244 24612
rect 6188 24558 6190 24610
rect 6190 24558 6242 24610
rect 6242 24558 6244 24610
rect 6188 24556 6244 24558
rect 5404 24108 5460 24164
rect 5964 23996 6020 24052
rect 5628 23938 5684 23940
rect 5628 23886 5630 23938
rect 5630 23886 5682 23938
rect 5682 23886 5684 23938
rect 5628 23884 5684 23886
rect 4844 23212 4900 23268
rect 5292 23154 5348 23156
rect 5292 23102 5294 23154
rect 5294 23102 5346 23154
rect 5346 23102 5348 23154
rect 5292 23100 5348 23102
rect 6636 24050 6692 24052
rect 6636 23998 6638 24050
rect 6638 23998 6690 24050
rect 6690 23998 6692 24050
rect 6636 23996 6692 23998
rect 6300 23884 6356 23940
rect 6188 23826 6244 23828
rect 6188 23774 6190 23826
rect 6190 23774 6242 23826
rect 6242 23774 6244 23826
rect 6188 23772 6244 23774
rect 7868 24050 7924 24052
rect 7868 23998 7870 24050
rect 7870 23998 7922 24050
rect 7922 23998 7924 24050
rect 7868 23996 7924 23998
rect 7756 23772 7812 23828
rect 9100 23938 9156 23940
rect 9100 23886 9102 23938
rect 9102 23886 9154 23938
rect 9154 23886 9156 23938
rect 9100 23884 9156 23886
rect 8764 23714 8820 23716
rect 8764 23662 8766 23714
rect 8766 23662 8818 23714
rect 8818 23662 8820 23714
rect 8764 23660 8820 23662
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 3612 22540 3668 22596
rect 4620 22540 4676 22596
rect 5404 22540 5460 22596
rect 3948 21756 4004 21812
rect 1820 20802 1876 20804
rect 1820 20750 1822 20802
rect 1822 20750 1874 20802
rect 1874 20750 1876 20802
rect 1820 20748 1876 20750
rect 5516 21756 5572 21812
rect 8988 22652 9044 22708
rect 10780 24556 10836 24612
rect 12236 25506 12292 25508
rect 12236 25454 12238 25506
rect 12238 25454 12290 25506
rect 12290 25454 12292 25506
rect 12236 25452 12292 25454
rect 12460 25506 12516 25508
rect 12460 25454 12462 25506
rect 12462 25454 12514 25506
rect 12514 25454 12516 25506
rect 12460 25452 12516 25454
rect 11900 24610 11956 24612
rect 11900 24558 11902 24610
rect 11902 24558 11954 24610
rect 11954 24558 11956 24610
rect 11900 24556 11956 24558
rect 11004 23996 11060 24052
rect 11676 24444 11732 24500
rect 12012 24444 12068 24500
rect 12124 24220 12180 24276
rect 12012 23884 12068 23940
rect 12012 23266 12068 23268
rect 12012 23214 12014 23266
rect 12014 23214 12066 23266
rect 12066 23214 12068 23266
rect 12012 23212 12068 23214
rect 11004 22652 11060 22708
rect 6636 22370 6692 22372
rect 6636 22318 6638 22370
rect 6638 22318 6690 22370
rect 6690 22318 6692 22370
rect 6636 22316 6692 22318
rect 10332 22316 10388 22372
rect 6188 21756 6244 21812
rect 6748 21756 6804 21812
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3948 20748 4004 20804
rect 2492 20130 2548 20132
rect 2492 20078 2494 20130
rect 2494 20078 2546 20130
rect 2546 20078 2548 20130
rect 2492 20076 2548 20078
rect 1708 18060 1764 18116
rect 2604 18620 2660 18676
rect 2268 18450 2324 18452
rect 2268 18398 2270 18450
rect 2270 18398 2322 18450
rect 2322 18398 2324 18450
rect 2268 18396 2324 18398
rect 2492 17724 2548 17780
rect 2716 18284 2772 18340
rect 3052 18562 3108 18564
rect 3052 18510 3054 18562
rect 3054 18510 3106 18562
rect 3106 18510 3108 18562
rect 3052 18508 3108 18510
rect 3164 18172 3220 18228
rect 4620 20076 4676 20132
rect 5068 20076 5124 20132
rect 4620 19906 4676 19908
rect 4620 19854 4622 19906
rect 4622 19854 4674 19906
rect 4674 19854 4676 19906
rect 4620 19852 4676 19854
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4284 18508 4340 18564
rect 3724 18450 3780 18452
rect 3724 18398 3726 18450
rect 3726 18398 3778 18450
rect 3778 18398 3780 18450
rect 3724 18396 3780 18398
rect 3948 18450 4004 18452
rect 3948 18398 3950 18450
rect 3950 18398 4002 18450
rect 4002 18398 4004 18450
rect 3948 18396 4004 18398
rect 3612 18338 3668 18340
rect 3612 18286 3614 18338
rect 3614 18286 3666 18338
rect 3666 18286 3668 18338
rect 3612 18284 3668 18286
rect 3500 18060 3556 18116
rect 3948 18060 4004 18116
rect 4620 18620 4676 18676
rect 5852 19292 5908 19348
rect 5964 19852 6020 19908
rect 6524 21308 6580 21364
rect 8764 21810 8820 21812
rect 8764 21758 8766 21810
rect 8766 21758 8818 21810
rect 8818 21758 8820 21810
rect 8764 21756 8820 21758
rect 9660 21810 9716 21812
rect 9660 21758 9662 21810
rect 9662 21758 9714 21810
rect 9714 21758 9716 21810
rect 9660 21756 9716 21758
rect 10220 21698 10276 21700
rect 10220 21646 10222 21698
rect 10222 21646 10274 21698
rect 10274 21646 10276 21698
rect 10220 21644 10276 21646
rect 7420 20130 7476 20132
rect 7420 20078 7422 20130
rect 7422 20078 7474 20130
rect 7474 20078 7476 20130
rect 7420 20076 7476 20078
rect 6076 19180 6132 19236
rect 8316 20242 8372 20244
rect 8316 20190 8318 20242
rect 8318 20190 8370 20242
rect 8370 20190 8372 20242
rect 8316 20188 8372 20190
rect 7532 19740 7588 19796
rect 7420 19234 7476 19236
rect 7420 19182 7422 19234
rect 7422 19182 7474 19234
rect 7474 19182 7476 19234
rect 7420 19180 7476 19182
rect 6748 19122 6804 19124
rect 6748 19070 6750 19122
rect 6750 19070 6802 19122
rect 6802 19070 6804 19122
rect 6748 19068 6804 19070
rect 8316 19292 8372 19348
rect 5516 18396 5572 18452
rect 1820 16940 1876 16996
rect 2828 16994 2884 16996
rect 2828 16942 2830 16994
rect 2830 16942 2882 16994
rect 2882 16942 2884 16994
rect 2828 16940 2884 16942
rect 2604 16716 2660 16772
rect 2268 15538 2324 15540
rect 2268 15486 2270 15538
rect 2270 15486 2322 15538
rect 2322 15486 2324 15538
rect 2268 15484 2324 15486
rect 2492 15986 2548 15988
rect 2492 15934 2494 15986
rect 2494 15934 2546 15986
rect 2546 15934 2548 15986
rect 2492 15932 2548 15934
rect 2828 15426 2884 15428
rect 2828 15374 2830 15426
rect 2830 15374 2882 15426
rect 2882 15374 2884 15426
rect 2828 15372 2884 15374
rect 3052 16716 3108 16772
rect 4172 17724 4228 17780
rect 3388 15932 3444 15988
rect 4172 15484 4228 15540
rect 3276 15314 3332 15316
rect 3276 15262 3278 15314
rect 3278 15262 3330 15314
rect 3330 15262 3332 15314
rect 3276 15260 3332 15262
rect 4508 18226 4564 18228
rect 4508 18174 4510 18226
rect 4510 18174 4562 18226
rect 4562 18174 4564 18226
rect 4508 18172 4564 18174
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4620 17778 4676 17780
rect 4620 17726 4622 17778
rect 4622 17726 4674 17778
rect 4674 17726 4676 17778
rect 4620 17724 4676 17726
rect 6300 17666 6356 17668
rect 6300 17614 6302 17666
rect 6302 17614 6354 17666
rect 6354 17614 6356 17666
rect 6300 17612 6356 17614
rect 5852 16828 5908 16884
rect 6524 17442 6580 17444
rect 6524 17390 6526 17442
rect 6526 17390 6578 17442
rect 6578 17390 6580 17442
rect 6524 17388 6580 17390
rect 5964 16716 6020 16772
rect 6524 16828 6580 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4620 15372 4676 15428
rect 3836 15148 3892 15204
rect 4844 15148 4900 15204
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 3612 14700 3668 14756
rect 4844 14812 4900 14868
rect 2940 14252 2996 14308
rect 2492 13804 2548 13860
rect 3164 13916 3220 13972
rect 3836 13692 3892 13748
rect 4396 13858 4452 13860
rect 4396 13806 4398 13858
rect 4398 13806 4450 13858
rect 4450 13806 4452 13858
rect 4396 13804 4452 13806
rect 5964 15484 6020 15540
rect 6412 16044 6468 16100
rect 5852 15372 5908 15428
rect 6188 15148 6244 15204
rect 5740 14812 5796 14868
rect 5628 14306 5684 14308
rect 5628 14254 5630 14306
rect 5630 14254 5682 14306
rect 5682 14254 5684 14306
rect 5628 14252 5684 14254
rect 4620 13692 4676 13748
rect 3276 13132 3332 13188
rect 3724 13580 3780 13636
rect 2492 13074 2548 13076
rect 2492 13022 2494 13074
rect 2494 13022 2546 13074
rect 2546 13022 2548 13074
rect 2492 13020 2548 13022
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4620 13132 4676 13188
rect 4508 12908 4564 12964
rect 3500 12402 3556 12404
rect 3500 12350 3502 12402
rect 3502 12350 3554 12402
rect 3554 12350 3556 12402
rect 3500 12348 3556 12350
rect 5516 13916 5572 13972
rect 5964 13916 6020 13972
rect 6300 14028 6356 14084
rect 4956 12908 5012 12964
rect 4844 12684 4900 12740
rect 1820 11452 1876 11508
rect 2492 12012 2548 12068
rect 4060 12066 4116 12068
rect 4060 12014 4062 12066
rect 4062 12014 4114 12066
rect 4114 12014 4116 12066
rect 4060 12012 4116 12014
rect 5628 12962 5684 12964
rect 5628 12910 5630 12962
rect 5630 12910 5682 12962
rect 5682 12910 5684 12962
rect 5628 12908 5684 12910
rect 5964 13020 6020 13076
rect 5180 12572 5236 12628
rect 5068 12348 5124 12404
rect 6748 15484 6804 15540
rect 6748 15314 6804 15316
rect 6748 15262 6750 15314
rect 6750 15262 6802 15314
rect 6802 15262 6804 15314
rect 6748 15260 6804 15262
rect 6524 15148 6580 15204
rect 7196 16828 7252 16884
rect 7084 16716 7140 16772
rect 6972 15426 7028 15428
rect 6972 15374 6974 15426
rect 6974 15374 7026 15426
rect 7026 15374 7028 15426
rect 6972 15372 7028 15374
rect 7756 18396 7812 18452
rect 9660 21362 9716 21364
rect 9660 21310 9662 21362
rect 9662 21310 9714 21362
rect 9714 21310 9716 21362
rect 9660 21308 9716 21310
rect 8652 19740 8708 19796
rect 8876 19180 8932 19236
rect 10108 20802 10164 20804
rect 10108 20750 10110 20802
rect 10110 20750 10162 20802
rect 10162 20750 10164 20802
rect 10108 20748 10164 20750
rect 10892 21698 10948 21700
rect 10892 21646 10894 21698
rect 10894 21646 10946 21698
rect 10946 21646 10948 21698
rect 10892 21644 10948 21646
rect 9436 19180 9492 19236
rect 7868 18284 7924 18340
rect 7532 18172 7588 18228
rect 7756 17612 7812 17668
rect 9772 19068 9828 19124
rect 9548 18396 9604 18452
rect 8316 18172 8372 18228
rect 8092 17388 8148 17444
rect 9436 17388 9492 17444
rect 8540 16882 8596 16884
rect 8540 16830 8542 16882
rect 8542 16830 8594 16882
rect 8594 16830 8596 16882
rect 8540 16828 8596 16830
rect 7980 16156 8036 16212
rect 8876 16098 8932 16100
rect 8876 16046 8878 16098
rect 8878 16046 8930 16098
rect 8930 16046 8932 16098
rect 8876 16044 8932 16046
rect 6860 15036 6916 15092
rect 6860 14700 6916 14756
rect 7084 14812 7140 14868
rect 6748 13916 6804 13972
rect 6636 13580 6692 13636
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 5516 11954 5572 11956
rect 5516 11902 5518 11954
rect 5518 11902 5570 11954
rect 5570 11902 5572 11954
rect 5516 11900 5572 11902
rect 5292 11452 5348 11508
rect 4284 10780 4340 10836
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4732 9826 4788 9828
rect 4732 9774 4734 9826
rect 4734 9774 4786 9826
rect 4786 9774 4788 9826
rect 4732 9772 4788 9774
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4620 8428 4676 8484
rect 5180 9714 5236 9716
rect 5180 9662 5182 9714
rect 5182 9662 5234 9714
rect 5234 9662 5236 9714
rect 5180 9660 5236 9662
rect 5516 10834 5572 10836
rect 5516 10782 5518 10834
rect 5518 10782 5570 10834
rect 5570 10782 5572 10834
rect 5516 10780 5572 10782
rect 6972 13356 7028 13412
rect 7196 14028 7252 14084
rect 8092 15036 8148 15092
rect 8092 14476 8148 14532
rect 8204 15372 8260 15428
rect 8092 14140 8148 14196
rect 8428 15484 8484 15540
rect 8764 15426 8820 15428
rect 8764 15374 8766 15426
rect 8766 15374 8818 15426
rect 8818 15374 8820 15426
rect 8764 15372 8820 15374
rect 9324 16098 9380 16100
rect 9324 16046 9326 16098
rect 9326 16046 9378 16098
rect 9378 16046 9380 16098
rect 9324 16044 9380 16046
rect 10556 20188 10612 20244
rect 10220 18338 10276 18340
rect 10220 18286 10222 18338
rect 10222 18286 10274 18338
rect 10274 18286 10276 18338
rect 10220 18284 10276 18286
rect 9660 17724 9716 17780
rect 9884 16882 9940 16884
rect 9884 16830 9886 16882
rect 9886 16830 9938 16882
rect 9938 16830 9940 16882
rect 9884 16828 9940 16830
rect 9548 16492 9604 16548
rect 9884 16268 9940 16324
rect 8988 15820 9044 15876
rect 8876 15148 8932 15204
rect 10108 16492 10164 16548
rect 10780 17778 10836 17780
rect 10780 17726 10782 17778
rect 10782 17726 10834 17778
rect 10834 17726 10836 17778
rect 10780 17724 10836 17726
rect 10668 16268 10724 16324
rect 10556 15874 10612 15876
rect 10556 15822 10558 15874
rect 10558 15822 10610 15874
rect 10610 15822 10612 15874
rect 10556 15820 10612 15822
rect 9884 15484 9940 15540
rect 9212 14924 9268 14980
rect 9548 14588 9604 14644
rect 9436 14530 9492 14532
rect 9436 14478 9438 14530
rect 9438 14478 9490 14530
rect 9490 14478 9492 14530
rect 9436 14476 9492 14478
rect 8316 14028 8372 14084
rect 7980 13746 8036 13748
rect 7980 13694 7982 13746
rect 7982 13694 8034 13746
rect 8034 13694 8036 13746
rect 7980 13692 8036 13694
rect 9772 14306 9828 14308
rect 9772 14254 9774 14306
rect 9774 14254 9826 14306
rect 9826 14254 9828 14306
rect 9772 14252 9828 14254
rect 8876 14028 8932 14084
rect 7644 13356 7700 13412
rect 10892 15372 10948 15428
rect 10108 15202 10164 15204
rect 10108 15150 10110 15202
rect 10110 15150 10162 15202
rect 10162 15150 10164 15202
rect 10108 15148 10164 15150
rect 9996 13970 10052 13972
rect 9996 13918 9998 13970
rect 9998 13918 10050 13970
rect 10050 13918 10052 13970
rect 9996 13916 10052 13918
rect 6636 12738 6692 12740
rect 6636 12686 6638 12738
rect 6638 12686 6690 12738
rect 6690 12686 6692 12738
rect 6636 12684 6692 12686
rect 5740 10834 5796 10836
rect 5740 10782 5742 10834
rect 5742 10782 5794 10834
rect 5794 10782 5796 10834
rect 5740 10780 5796 10782
rect 6412 10780 6468 10836
rect 7196 11900 7252 11956
rect 7644 12348 7700 12404
rect 10556 14252 10612 14308
rect 10332 13858 10388 13860
rect 10332 13806 10334 13858
rect 10334 13806 10386 13858
rect 10386 13806 10388 13858
rect 10332 13804 10388 13806
rect 10892 13746 10948 13748
rect 10892 13694 10894 13746
rect 10894 13694 10946 13746
rect 10946 13694 10948 13746
rect 10892 13692 10948 13694
rect 9772 12402 9828 12404
rect 9772 12350 9774 12402
rect 9774 12350 9826 12402
rect 9826 12350 9828 12402
rect 9772 12348 9828 12350
rect 8764 11506 8820 11508
rect 8764 11454 8766 11506
rect 8766 11454 8818 11506
rect 8818 11454 8820 11506
rect 8764 11452 8820 11454
rect 9100 11676 9156 11732
rect 9996 11676 10052 11732
rect 5852 9996 5908 10052
rect 7644 9996 7700 10052
rect 9772 10444 9828 10500
rect 5964 9548 6020 9604
rect 5180 8540 5236 8596
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 5068 6748 5124 6804
rect 5292 8428 5348 8484
rect 6636 8652 6692 8708
rect 5292 7980 5348 8036
rect 6076 7532 6132 7588
rect 6524 7420 6580 7476
rect 6188 6860 6244 6916
rect 6300 6690 6356 6692
rect 6300 6638 6302 6690
rect 6302 6638 6354 6690
rect 6354 6638 6356 6690
rect 6300 6636 6356 6638
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 5180 5794 5236 5796
rect 5180 5742 5182 5794
rect 5182 5742 5234 5794
rect 5234 5742 5236 5794
rect 5180 5740 5236 5742
rect 5180 5404 5236 5460
rect 4844 5292 4900 5348
rect 5068 4956 5124 5012
rect 6076 5740 6132 5796
rect 5516 4956 5572 5012
rect 5852 4226 5908 4228
rect 5852 4174 5854 4226
rect 5854 4174 5906 4226
rect 5906 4174 5908 4226
rect 5852 4172 5908 4174
rect 5068 4060 5124 4116
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 6636 6972 6692 7028
rect 6636 6748 6692 6804
rect 7196 9602 7252 9604
rect 7196 9550 7198 9602
rect 7198 9550 7250 9602
rect 7250 9550 7252 9602
rect 7196 9548 7252 9550
rect 7644 9602 7700 9604
rect 7644 9550 7646 9602
rect 7646 9550 7698 9602
rect 7698 9550 7700 9602
rect 7644 9548 7700 9550
rect 8204 10108 8260 10164
rect 8092 9548 8148 9604
rect 8204 9884 8260 9940
rect 7084 8316 7140 8372
rect 8316 9548 8372 9604
rect 7756 8258 7812 8260
rect 7756 8206 7758 8258
rect 7758 8206 7810 8258
rect 7810 8206 7812 8258
rect 7756 8204 7812 8206
rect 6972 8146 7028 8148
rect 6972 8094 6974 8146
rect 6974 8094 7026 8146
rect 7026 8094 7028 8146
rect 6972 8092 7028 8094
rect 7084 8034 7140 8036
rect 7084 7982 7086 8034
rect 7086 7982 7138 8034
rect 7138 7982 7140 8034
rect 7084 7980 7140 7982
rect 7532 8034 7588 8036
rect 7532 7982 7534 8034
rect 7534 7982 7586 8034
rect 7586 7982 7588 8034
rect 7532 7980 7588 7982
rect 7868 7980 7924 8036
rect 8540 9324 8596 9380
rect 8428 8258 8484 8260
rect 8428 8206 8430 8258
rect 8430 8206 8482 8258
rect 8482 8206 8484 8258
rect 8428 8204 8484 8206
rect 7756 7196 7812 7252
rect 8092 7196 8148 7252
rect 7084 6914 7140 6916
rect 7084 6862 7086 6914
rect 7086 6862 7138 6914
rect 7138 6862 7140 6914
rect 7084 6860 7140 6862
rect 8428 7420 8484 7476
rect 6524 5292 6580 5348
rect 6860 4898 6916 4900
rect 6860 4846 6862 4898
rect 6862 4846 6914 4898
rect 6914 4846 6916 4898
rect 6860 4844 6916 4846
rect 4732 3276 4788 3332
rect 5516 3330 5572 3332
rect 5516 3278 5518 3330
rect 5518 3278 5570 3330
rect 5570 3278 5572 3330
rect 5516 3276 5572 3278
rect 9436 10332 9492 10388
rect 8652 8370 8708 8372
rect 8652 8318 8654 8370
rect 8654 8318 8706 8370
rect 8706 8318 8708 8370
rect 8652 8316 8708 8318
rect 8652 7868 8708 7924
rect 8988 9266 9044 9268
rect 8988 9214 8990 9266
rect 8990 9214 9042 9266
rect 9042 9214 9044 9266
rect 8988 9212 9044 9214
rect 8540 6748 8596 6804
rect 8988 8034 9044 8036
rect 8988 7982 8990 8034
rect 8990 7982 9042 8034
rect 9042 7982 9044 8034
rect 8988 7980 9044 7982
rect 8988 7474 9044 7476
rect 8988 7422 8990 7474
rect 8990 7422 9042 7474
rect 9042 7422 9044 7474
rect 8988 7420 9044 7422
rect 9660 7644 9716 7700
rect 9884 8764 9940 8820
rect 9884 8146 9940 8148
rect 9884 8094 9886 8146
rect 9886 8094 9938 8146
rect 9938 8094 9940 8146
rect 9884 8092 9940 8094
rect 8764 6636 8820 6692
rect 8428 6524 8484 6580
rect 8428 5122 8484 5124
rect 8428 5070 8430 5122
rect 8430 5070 8482 5122
rect 8482 5070 8484 5122
rect 8428 5068 8484 5070
rect 8540 4844 8596 4900
rect 8428 4226 8484 4228
rect 8428 4174 8430 4226
rect 8430 4174 8482 4226
rect 8482 4174 8484 4226
rect 8428 4172 8484 4174
rect 10556 10610 10612 10612
rect 10556 10558 10558 10610
rect 10558 10558 10610 10610
rect 10610 10558 10612 10610
rect 10556 10556 10612 10558
rect 11340 22370 11396 22372
rect 11340 22318 11342 22370
rect 11342 22318 11394 22370
rect 11394 22318 11396 22370
rect 11340 22316 11396 22318
rect 11452 21756 11508 21812
rect 11228 21474 11284 21476
rect 11228 21422 11230 21474
rect 11230 21422 11282 21474
rect 11282 21422 11284 21474
rect 11228 21420 11284 21422
rect 11788 21474 11844 21476
rect 11788 21422 11790 21474
rect 11790 21422 11842 21474
rect 11842 21422 11844 21474
rect 11788 21420 11844 21422
rect 13244 27244 13300 27300
rect 13804 27970 13860 27972
rect 13804 27918 13806 27970
rect 13806 27918 13858 27970
rect 13858 27918 13860 27970
rect 13804 27916 13860 27918
rect 13692 27746 13748 27748
rect 13692 27694 13694 27746
rect 13694 27694 13746 27746
rect 13746 27694 13748 27746
rect 13692 27692 13748 27694
rect 14700 29314 14756 29316
rect 14700 29262 14702 29314
rect 14702 29262 14754 29314
rect 14754 29262 14756 29314
rect 14700 29260 14756 29262
rect 15036 29986 15092 29988
rect 15036 29934 15038 29986
rect 15038 29934 15090 29986
rect 15090 29934 15092 29986
rect 15036 29932 15092 29934
rect 15484 29260 15540 29316
rect 14924 28700 14980 28756
rect 14700 27916 14756 27972
rect 15260 27916 15316 27972
rect 15036 27858 15092 27860
rect 15036 27806 15038 27858
rect 15038 27806 15090 27858
rect 15090 27806 15092 27858
rect 15036 27804 15092 27806
rect 15260 27244 15316 27300
rect 13580 26402 13636 26404
rect 13580 26350 13582 26402
rect 13582 26350 13634 26402
rect 13634 26350 13636 26402
rect 13580 26348 13636 26350
rect 13916 26796 13972 26852
rect 13692 26290 13748 26292
rect 13692 26238 13694 26290
rect 13694 26238 13746 26290
rect 13746 26238 13748 26290
rect 13692 26236 13748 26238
rect 14140 26348 14196 26404
rect 14588 26290 14644 26292
rect 14588 26238 14590 26290
rect 14590 26238 14642 26290
rect 14642 26238 14644 26290
rect 14588 26236 14644 26238
rect 14476 25730 14532 25732
rect 14476 25678 14478 25730
rect 14478 25678 14530 25730
rect 14530 25678 14532 25730
rect 14476 25676 14532 25678
rect 15484 26908 15540 26964
rect 15260 25900 15316 25956
rect 16044 30940 16100 30996
rect 16604 32562 16660 32564
rect 16604 32510 16606 32562
rect 16606 32510 16658 32562
rect 16658 32510 16660 32562
rect 16604 32508 16660 32510
rect 17388 33068 17444 33124
rect 17612 33180 17668 33236
rect 17276 32562 17332 32564
rect 17276 32510 17278 32562
rect 17278 32510 17330 32562
rect 17330 32510 17332 32562
rect 17276 32508 17332 32510
rect 16828 32396 16884 32452
rect 17276 32060 17332 32116
rect 16828 31836 16884 31892
rect 16716 31164 16772 31220
rect 16268 30716 16324 30772
rect 15708 29932 15764 29988
rect 16268 28588 16324 28644
rect 17052 28642 17108 28644
rect 17052 28590 17054 28642
rect 17054 28590 17106 28642
rect 17106 28590 17108 28642
rect 17052 28588 17108 28590
rect 16380 28082 16436 28084
rect 16380 28030 16382 28082
rect 16382 28030 16434 28082
rect 16434 28030 16436 28082
rect 16380 28028 16436 28030
rect 16716 28252 16772 28308
rect 16604 27970 16660 27972
rect 16604 27918 16606 27970
rect 16606 27918 16658 27970
rect 16658 27918 16660 27970
rect 16604 27916 16660 27918
rect 15932 27804 15988 27860
rect 15820 27244 15876 27300
rect 15708 26402 15764 26404
rect 15708 26350 15710 26402
rect 15710 26350 15762 26402
rect 15762 26350 15764 26402
rect 15708 26348 15764 26350
rect 15820 26290 15876 26292
rect 15820 26238 15822 26290
rect 15822 26238 15874 26290
rect 15874 26238 15876 26290
rect 15820 26236 15876 26238
rect 16156 27858 16212 27860
rect 16156 27806 16158 27858
rect 16158 27806 16210 27858
rect 16210 27806 16212 27858
rect 16156 27804 16212 27806
rect 16492 27804 16548 27860
rect 16828 27356 16884 27412
rect 16604 27074 16660 27076
rect 16604 27022 16606 27074
rect 16606 27022 16658 27074
rect 16658 27022 16660 27074
rect 16604 27020 16660 27022
rect 16380 26962 16436 26964
rect 16380 26910 16382 26962
rect 16382 26910 16434 26962
rect 16434 26910 16436 26962
rect 16380 26908 16436 26910
rect 17164 27020 17220 27076
rect 16716 26850 16772 26852
rect 16716 26798 16718 26850
rect 16718 26798 16770 26850
rect 16770 26798 16772 26850
rect 16716 26796 16772 26798
rect 16492 26514 16548 26516
rect 16492 26462 16494 26514
rect 16494 26462 16546 26514
rect 16546 26462 16548 26514
rect 16492 26460 16548 26462
rect 16044 25900 16100 25956
rect 14140 25452 14196 25508
rect 14812 25228 14868 25284
rect 16156 25676 16212 25732
rect 16044 25394 16100 25396
rect 16044 25342 16046 25394
rect 16046 25342 16098 25394
rect 16098 25342 16100 25394
rect 16044 25340 16100 25342
rect 13020 24668 13076 24724
rect 12572 24444 12628 24500
rect 12908 24162 12964 24164
rect 12908 24110 12910 24162
rect 12910 24110 12962 24162
rect 12962 24110 12964 24162
rect 12908 24108 12964 24110
rect 12348 24050 12404 24052
rect 12348 23998 12350 24050
rect 12350 23998 12402 24050
rect 12402 23998 12404 24050
rect 12348 23996 12404 23998
rect 12236 23884 12292 23940
rect 13132 23772 13188 23828
rect 13132 23212 13188 23268
rect 13916 24444 13972 24500
rect 13468 24220 13524 24276
rect 11116 20748 11172 20804
rect 14028 24108 14084 24164
rect 14028 23826 14084 23828
rect 14028 23774 14030 23826
rect 14030 23774 14082 23826
rect 14082 23774 14084 23826
rect 14028 23772 14084 23774
rect 14028 21810 14084 21812
rect 14028 21758 14030 21810
rect 14030 21758 14082 21810
rect 14082 21758 14084 21810
rect 14028 21756 14084 21758
rect 14588 24834 14644 24836
rect 14588 24782 14590 24834
rect 14590 24782 14642 24834
rect 14642 24782 14644 24834
rect 14588 24780 14644 24782
rect 14700 24610 14756 24612
rect 14700 24558 14702 24610
rect 14702 24558 14754 24610
rect 14754 24558 14756 24610
rect 14700 24556 14756 24558
rect 14252 23938 14308 23940
rect 14252 23886 14254 23938
rect 14254 23886 14306 23938
rect 14306 23886 14308 23938
rect 14252 23884 14308 23886
rect 15260 24556 15316 24612
rect 15036 23772 15092 23828
rect 15260 23772 15316 23828
rect 15036 23436 15092 23492
rect 14588 22988 14644 23044
rect 12684 20748 12740 20804
rect 14140 20802 14196 20804
rect 14140 20750 14142 20802
rect 14142 20750 14194 20802
rect 14194 20750 14196 20802
rect 14140 20748 14196 20750
rect 14924 20524 14980 20580
rect 15596 24610 15652 24612
rect 15596 24558 15598 24610
rect 15598 24558 15650 24610
rect 15650 24558 15652 24610
rect 15596 24556 15652 24558
rect 16604 26290 16660 26292
rect 16604 26238 16606 26290
rect 16606 26238 16658 26290
rect 16658 26238 16660 26290
rect 16604 26236 16660 26238
rect 16828 25564 16884 25620
rect 16716 25506 16772 25508
rect 16716 25454 16718 25506
rect 16718 25454 16770 25506
rect 16770 25454 16772 25506
rect 16716 25452 16772 25454
rect 16380 25228 16436 25284
rect 17052 25228 17108 25284
rect 16156 24556 16212 24612
rect 15484 23884 15540 23940
rect 16492 24108 16548 24164
rect 15820 23436 15876 23492
rect 16604 23772 16660 23828
rect 17612 32172 17668 32228
rect 17724 33068 17780 33124
rect 17500 31836 17556 31892
rect 17388 31218 17444 31220
rect 17388 31166 17390 31218
rect 17390 31166 17442 31218
rect 17442 31166 17444 31218
rect 17388 31164 17444 31166
rect 17724 31052 17780 31108
rect 18172 33346 18228 33348
rect 18172 33294 18174 33346
rect 18174 33294 18226 33346
rect 18226 33294 18228 33346
rect 18172 33292 18228 33294
rect 18060 33068 18116 33124
rect 18284 33122 18340 33124
rect 18284 33070 18286 33122
rect 18286 33070 18338 33122
rect 18338 33070 18340 33122
rect 18284 33068 18340 33070
rect 17836 31948 17892 32004
rect 18060 32172 18116 32228
rect 18508 32732 18564 32788
rect 18732 32732 18788 32788
rect 18620 32620 18676 32676
rect 18172 32060 18228 32116
rect 18172 31724 18228 31780
rect 17724 30770 17780 30772
rect 17724 30718 17726 30770
rect 17726 30718 17778 30770
rect 17778 30718 17780 30770
rect 17724 30716 17780 30718
rect 17500 30268 17556 30324
rect 18284 31388 18340 31444
rect 18396 31948 18452 32004
rect 18284 31106 18340 31108
rect 18284 31054 18286 31106
rect 18286 31054 18338 31106
rect 18338 31054 18340 31106
rect 18284 31052 18340 31054
rect 18508 31164 18564 31220
rect 19068 33122 19124 33124
rect 19068 33070 19070 33122
rect 19070 33070 19122 33122
rect 19122 33070 19124 33122
rect 19068 33068 19124 33070
rect 18956 32620 19012 32676
rect 19068 32732 19124 32788
rect 20412 34018 20468 34020
rect 20412 33966 20414 34018
rect 20414 33966 20466 34018
rect 20466 33966 20468 34018
rect 20412 33964 20468 33966
rect 19404 33404 19460 33460
rect 19292 33234 19348 33236
rect 19292 33182 19294 33234
rect 19294 33182 19346 33234
rect 19346 33182 19348 33234
rect 19292 33180 19348 33182
rect 19404 32956 19460 33012
rect 18844 32508 18900 32564
rect 18956 31500 19012 31556
rect 18844 30882 18900 30884
rect 18844 30830 18846 30882
rect 18846 30830 18898 30882
rect 18898 30830 18900 30882
rect 18844 30828 18900 30830
rect 18620 30716 18676 30772
rect 18396 30098 18452 30100
rect 18396 30046 18398 30098
rect 18398 30046 18450 30098
rect 18450 30046 18452 30098
rect 18396 30044 18452 30046
rect 17836 28530 17892 28532
rect 17836 28478 17838 28530
rect 17838 28478 17890 28530
rect 17890 28478 17892 28530
rect 17836 28476 17892 28478
rect 17724 28364 17780 28420
rect 17388 27858 17444 27860
rect 17388 27806 17390 27858
rect 17390 27806 17442 27858
rect 17442 27806 17444 27858
rect 17388 27804 17444 27806
rect 17388 27298 17444 27300
rect 17388 27246 17390 27298
rect 17390 27246 17442 27298
rect 17442 27246 17444 27298
rect 17388 27244 17444 27246
rect 17388 26796 17444 26852
rect 17836 26796 17892 26852
rect 17948 27580 18004 27636
rect 17612 26514 17668 26516
rect 17612 26462 17614 26514
rect 17614 26462 17666 26514
rect 17666 26462 17668 26514
rect 17612 26460 17668 26462
rect 17836 26402 17892 26404
rect 17836 26350 17838 26402
rect 17838 26350 17890 26402
rect 17890 26350 17892 26402
rect 17836 26348 17892 26350
rect 17500 26236 17556 26292
rect 18172 27858 18228 27860
rect 18172 27806 18174 27858
rect 18174 27806 18226 27858
rect 18226 27806 18228 27858
rect 18172 27804 18228 27806
rect 18396 27634 18452 27636
rect 18396 27582 18398 27634
rect 18398 27582 18450 27634
rect 18450 27582 18452 27634
rect 18396 27580 18452 27582
rect 18284 27468 18340 27524
rect 18060 27020 18116 27076
rect 18732 28252 18788 28308
rect 18284 27244 18340 27300
rect 18620 27356 18676 27412
rect 18508 27020 18564 27076
rect 20188 33404 20244 33460
rect 19516 32732 19572 32788
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19516 32562 19572 32564
rect 19516 32510 19518 32562
rect 19518 32510 19570 32562
rect 19570 32510 19572 32562
rect 19516 32508 19572 32510
rect 19180 31836 19236 31892
rect 20076 32786 20132 32788
rect 20076 32734 20078 32786
rect 20078 32734 20130 32786
rect 20130 32734 20132 32786
rect 20076 32732 20132 32734
rect 20412 33068 20468 33124
rect 20412 32674 20468 32676
rect 20412 32622 20414 32674
rect 20414 32622 20466 32674
rect 20466 32622 20468 32674
rect 20412 32620 20468 32622
rect 20300 32508 20356 32564
rect 19404 31724 19460 31780
rect 20412 31724 20468 31780
rect 19852 31612 19908 31668
rect 20524 31612 20580 31668
rect 19180 31388 19236 31444
rect 19628 31554 19684 31556
rect 19628 31502 19630 31554
rect 19630 31502 19682 31554
rect 19682 31502 19684 31554
rect 19628 31500 19684 31502
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20188 31388 20244 31444
rect 19404 29596 19460 29652
rect 19180 28476 19236 28532
rect 19404 28364 19460 28420
rect 19292 27916 19348 27972
rect 19180 27468 19236 27524
rect 17948 25618 18004 25620
rect 17948 25566 17950 25618
rect 17950 25566 18002 25618
rect 18002 25566 18004 25618
rect 17948 25564 18004 25566
rect 17724 25452 17780 25508
rect 17836 25116 17892 25172
rect 17164 24108 17220 24164
rect 17052 24050 17108 24052
rect 17052 23998 17054 24050
rect 17054 23998 17106 24050
rect 17106 23998 17108 24050
rect 17052 23996 17108 23998
rect 15484 23042 15540 23044
rect 15484 22990 15486 23042
rect 15486 22990 15538 23042
rect 15538 22990 15540 23042
rect 15484 22988 15540 22990
rect 16044 22988 16100 23044
rect 17276 22876 17332 22932
rect 17052 22540 17108 22596
rect 16044 21586 16100 21588
rect 16044 21534 16046 21586
rect 16046 21534 16098 21586
rect 16098 21534 16100 21586
rect 16044 21532 16100 21534
rect 16492 21474 16548 21476
rect 16492 21422 16494 21474
rect 16494 21422 16546 21474
rect 16546 21422 16548 21474
rect 16492 21420 16548 21422
rect 17836 24780 17892 24836
rect 18508 25564 18564 25620
rect 18396 25452 18452 25508
rect 18284 25228 18340 25284
rect 17388 21308 17444 21364
rect 17500 23938 17556 23940
rect 17500 23886 17502 23938
rect 17502 23886 17554 23938
rect 17554 23886 17556 23938
rect 17500 23884 17556 23886
rect 16828 21196 16884 21252
rect 17052 20748 17108 20804
rect 16604 20636 16660 20692
rect 15372 20300 15428 20356
rect 13804 20076 13860 20132
rect 14140 20076 14196 20132
rect 13692 19964 13748 20020
rect 12796 19740 12852 19796
rect 12124 18956 12180 19012
rect 11116 17724 11172 17780
rect 11228 17442 11284 17444
rect 11228 17390 11230 17442
rect 11230 17390 11282 17442
rect 11282 17390 11284 17442
rect 11228 17388 11284 17390
rect 11228 16268 11284 16324
rect 11116 15932 11172 15988
rect 12348 16492 12404 16548
rect 12124 15708 12180 15764
rect 11788 15036 11844 15092
rect 11116 14140 11172 14196
rect 11564 13858 11620 13860
rect 11564 13806 11566 13858
rect 11566 13806 11618 13858
rect 11618 13806 11620 13858
rect 11564 13804 11620 13806
rect 11116 13244 11172 13300
rect 11676 12962 11732 12964
rect 11676 12910 11678 12962
rect 11678 12910 11730 12962
rect 11730 12910 11732 12962
rect 11676 12908 11732 12910
rect 12124 14140 12180 14196
rect 13916 19794 13972 19796
rect 13916 19742 13918 19794
rect 13918 19742 13970 19794
rect 13970 19742 13972 19794
rect 13916 19740 13972 19742
rect 14028 19234 14084 19236
rect 14028 19182 14030 19234
rect 14030 19182 14082 19234
rect 14082 19182 14084 19234
rect 14028 19180 14084 19182
rect 13804 19122 13860 19124
rect 13804 19070 13806 19122
rect 13806 19070 13858 19122
rect 13858 19070 13860 19122
rect 13804 19068 13860 19070
rect 13580 18620 13636 18676
rect 13916 18508 13972 18564
rect 14364 20018 14420 20020
rect 14364 19966 14366 20018
rect 14366 19966 14418 20018
rect 14418 19966 14420 20018
rect 14364 19964 14420 19966
rect 14252 19010 14308 19012
rect 14252 18958 14254 19010
rect 14254 18958 14306 19010
rect 14306 18958 14308 19010
rect 14252 18956 14308 18958
rect 14700 19628 14756 19684
rect 14812 19234 14868 19236
rect 14812 19182 14814 19234
rect 14814 19182 14866 19234
rect 14866 19182 14868 19234
rect 14812 19180 14868 19182
rect 15932 20076 15988 20132
rect 15148 19852 15204 19908
rect 15372 19628 15428 19684
rect 16044 20018 16100 20020
rect 16044 19966 16046 20018
rect 16046 19966 16098 20018
rect 16098 19966 16100 20018
rect 16044 19964 16100 19966
rect 15484 19740 15540 19796
rect 16044 19740 16100 19796
rect 16268 19740 16324 19796
rect 15148 18508 15204 18564
rect 14812 18450 14868 18452
rect 14812 18398 14814 18450
rect 14814 18398 14866 18450
rect 14866 18398 14868 18450
rect 14812 18396 14868 18398
rect 16268 19068 16324 19124
rect 15708 18508 15764 18564
rect 15260 18450 15316 18452
rect 15260 18398 15262 18450
rect 15262 18398 15314 18450
rect 15314 18398 15316 18450
rect 15260 18396 15316 18398
rect 15036 18284 15092 18340
rect 12908 17724 12964 17780
rect 12908 17442 12964 17444
rect 12908 17390 12910 17442
rect 12910 17390 12962 17442
rect 12962 17390 12964 17442
rect 12908 17388 12964 17390
rect 13692 17778 13748 17780
rect 13692 17726 13694 17778
rect 13694 17726 13746 17778
rect 13746 17726 13748 17778
rect 13692 17724 13748 17726
rect 12796 16492 12852 16548
rect 12460 14476 12516 14532
rect 11900 13970 11956 13972
rect 11900 13918 11902 13970
rect 11902 13918 11954 13970
rect 11954 13918 11956 13970
rect 11900 13916 11956 13918
rect 12572 16268 12628 16324
rect 12684 15986 12740 15988
rect 12684 15934 12686 15986
rect 12686 15934 12738 15986
rect 12738 15934 12740 15986
rect 12684 15932 12740 15934
rect 13020 15986 13076 15988
rect 13020 15934 13022 15986
rect 13022 15934 13074 15986
rect 13074 15934 13076 15986
rect 13020 15932 13076 15934
rect 12796 15708 12852 15764
rect 13692 15932 13748 15988
rect 13580 15260 13636 15316
rect 13804 15708 13860 15764
rect 12684 13916 12740 13972
rect 12908 14642 12964 14644
rect 12908 14590 12910 14642
rect 12910 14590 12962 14642
rect 12962 14590 12964 14642
rect 12908 14588 12964 14590
rect 14140 17388 14196 17444
rect 14028 15708 14084 15764
rect 14476 15874 14532 15876
rect 14476 15822 14478 15874
rect 14478 15822 14530 15874
rect 14530 15822 14532 15874
rect 14476 15820 14532 15822
rect 14812 15708 14868 15764
rect 14252 15372 14308 15428
rect 17388 20636 17444 20692
rect 16828 19906 16884 19908
rect 16828 19854 16830 19906
rect 16830 19854 16882 19906
rect 16882 19854 16884 19906
rect 16828 19852 16884 19854
rect 17948 21196 18004 21252
rect 16716 19794 16772 19796
rect 16716 19742 16718 19794
rect 16718 19742 16770 19794
rect 16770 19742 16772 19794
rect 16716 19740 16772 19742
rect 17836 20578 17892 20580
rect 17836 20526 17838 20578
rect 17838 20526 17890 20578
rect 17890 20526 17892 20578
rect 17836 20524 17892 20526
rect 18172 20914 18228 20916
rect 18172 20862 18174 20914
rect 18174 20862 18226 20914
rect 18226 20862 18228 20914
rect 18172 20860 18228 20862
rect 17724 19628 17780 19684
rect 15820 18172 15876 18228
rect 15708 17948 15764 18004
rect 16492 18450 16548 18452
rect 16492 18398 16494 18450
rect 16494 18398 16546 18450
rect 16546 18398 16548 18450
rect 16492 18396 16548 18398
rect 16380 17836 16436 17892
rect 16828 17724 16884 17780
rect 15372 17612 15428 17668
rect 16492 17612 16548 17668
rect 15484 15986 15540 15988
rect 15484 15934 15486 15986
rect 15486 15934 15538 15986
rect 15538 15934 15540 15986
rect 15484 15932 15540 15934
rect 16828 16882 16884 16884
rect 16828 16830 16830 16882
rect 16830 16830 16882 16882
rect 16882 16830 16884 16882
rect 16828 16828 16884 16830
rect 17276 18620 17332 18676
rect 17612 18674 17668 18676
rect 17612 18622 17614 18674
rect 17614 18622 17666 18674
rect 17666 18622 17668 18674
rect 17612 18620 17668 18622
rect 17500 18508 17556 18564
rect 17388 17948 17444 18004
rect 17836 18284 17892 18340
rect 17836 18060 17892 18116
rect 17164 16210 17220 16212
rect 17164 16158 17166 16210
rect 17166 16158 17218 16210
rect 17218 16158 17220 16210
rect 17164 16156 17220 16158
rect 17276 16098 17332 16100
rect 17276 16046 17278 16098
rect 17278 16046 17330 16098
rect 17330 16046 17332 16098
rect 17276 16044 17332 16046
rect 17836 16044 17892 16100
rect 17612 15932 17668 15988
rect 15148 15874 15204 15876
rect 15148 15822 15150 15874
rect 15150 15822 15202 15874
rect 15202 15822 15204 15874
rect 15148 15820 15204 15822
rect 15036 15484 15092 15540
rect 14476 15260 14532 15316
rect 14140 15148 14196 15204
rect 14140 14588 14196 14644
rect 12124 13356 12180 13412
rect 11900 13074 11956 13076
rect 11900 13022 11902 13074
rect 11902 13022 11954 13074
rect 11954 13022 11956 13074
rect 11900 13020 11956 13022
rect 12348 13356 12404 13412
rect 12348 13020 12404 13076
rect 12460 12962 12516 12964
rect 12460 12910 12462 12962
rect 12462 12910 12514 12962
rect 12514 12910 12516 12962
rect 12460 12908 12516 12910
rect 14028 13356 14084 13412
rect 13244 12908 13300 12964
rect 12908 12850 12964 12852
rect 12908 12798 12910 12850
rect 12910 12798 12962 12850
rect 12962 12798 12964 12850
rect 12908 12796 12964 12798
rect 13692 12796 13748 12852
rect 11564 11228 11620 11284
rect 11004 10892 11060 10948
rect 10780 9266 10836 9268
rect 10780 9214 10782 9266
rect 10782 9214 10834 9266
rect 10834 9214 10836 9266
rect 10780 9212 10836 9214
rect 11228 10610 11284 10612
rect 11228 10558 11230 10610
rect 11230 10558 11282 10610
rect 11282 10558 11284 10610
rect 11228 10556 11284 10558
rect 11004 9548 11060 9604
rect 10444 8930 10500 8932
rect 10444 8878 10446 8930
rect 10446 8878 10498 8930
rect 10498 8878 10500 8930
rect 10444 8876 10500 8878
rect 10108 6524 10164 6580
rect 8876 5740 8932 5796
rect 8988 5122 9044 5124
rect 8988 5070 8990 5122
rect 8990 5070 9042 5122
rect 9042 5070 9044 5122
rect 8988 5068 9044 5070
rect 8876 4956 8932 5012
rect 8764 4060 8820 4116
rect 11340 9884 11396 9940
rect 11900 10386 11956 10388
rect 11900 10334 11902 10386
rect 11902 10334 11954 10386
rect 11954 10334 11956 10386
rect 11900 10332 11956 10334
rect 11564 9938 11620 9940
rect 11564 9886 11566 9938
rect 11566 9886 11618 9938
rect 11618 9886 11620 9938
rect 11564 9884 11620 9886
rect 11676 9548 11732 9604
rect 12236 9548 12292 9604
rect 12012 9324 12068 9380
rect 12796 11452 12852 11508
rect 12572 11282 12628 11284
rect 12572 11230 12574 11282
rect 12574 11230 12626 11282
rect 12626 11230 12628 11282
rect 12572 11228 12628 11230
rect 17276 15484 17332 15540
rect 14140 12572 14196 12628
rect 14364 12962 14420 12964
rect 14364 12910 14366 12962
rect 14366 12910 14418 12962
rect 14418 12910 14420 12962
rect 14364 12908 14420 12910
rect 14140 12066 14196 12068
rect 14140 12014 14142 12066
rect 14142 12014 14194 12066
rect 14194 12014 14196 12066
rect 14140 12012 14196 12014
rect 13804 11452 13860 11508
rect 14476 12178 14532 12180
rect 14476 12126 14478 12178
rect 14478 12126 14530 12178
rect 14530 12126 14532 12178
rect 14476 12124 14532 12126
rect 12460 9938 12516 9940
rect 12460 9886 12462 9938
rect 12462 9886 12514 9938
rect 12514 9886 12516 9938
rect 12460 9884 12516 9886
rect 13020 10444 13076 10500
rect 13580 10556 13636 10612
rect 12908 9826 12964 9828
rect 12908 9774 12910 9826
rect 12910 9774 12962 9826
rect 12962 9774 12964 9826
rect 12908 9772 12964 9774
rect 14700 12012 14756 12068
rect 14476 10892 14532 10948
rect 13692 10444 13748 10500
rect 13916 10556 13972 10612
rect 13692 9436 13748 9492
rect 11900 8818 11956 8820
rect 11900 8766 11902 8818
rect 11902 8766 11954 8818
rect 11954 8766 11956 8818
rect 11900 8764 11956 8766
rect 11676 8370 11732 8372
rect 11676 8318 11678 8370
rect 11678 8318 11730 8370
rect 11730 8318 11732 8370
rect 11676 8316 11732 8318
rect 10668 8146 10724 8148
rect 10668 8094 10670 8146
rect 10670 8094 10722 8146
rect 10722 8094 10724 8146
rect 10668 8092 10724 8094
rect 10556 6748 10612 6804
rect 10892 6972 10948 7028
rect 10444 5852 10500 5908
rect 9996 5794 10052 5796
rect 9996 5742 9998 5794
rect 9998 5742 10050 5794
rect 10050 5742 10052 5794
rect 9996 5740 10052 5742
rect 9436 3948 9492 4004
rect 9100 3836 9156 3892
rect 8652 3724 8708 3780
rect 9660 4898 9716 4900
rect 9660 4846 9662 4898
rect 9662 4846 9714 4898
rect 9714 4846 9716 4898
rect 9660 4844 9716 4846
rect 10780 5010 10836 5012
rect 10780 4958 10782 5010
rect 10782 4958 10834 5010
rect 10834 4958 10836 5010
rect 10780 4956 10836 4958
rect 10444 4844 10500 4900
rect 9772 3836 9828 3892
rect 8764 3500 8820 3556
rect 8204 3388 8260 3444
rect 6972 2716 7028 2772
rect 7868 3330 7924 3332
rect 7868 3278 7870 3330
rect 7870 3278 7922 3330
rect 7922 3278 7924 3330
rect 7868 3276 7924 3278
rect 10220 3948 10276 4004
rect 11788 4956 11844 5012
rect 10892 4620 10948 4676
rect 11228 4844 11284 4900
rect 10780 3778 10836 3780
rect 10780 3726 10782 3778
rect 10782 3726 10834 3778
rect 10834 3726 10836 3778
rect 10780 3724 10836 3726
rect 11676 4508 11732 4564
rect 11340 4396 11396 4452
rect 11676 3836 11732 3892
rect 12012 7532 12068 7588
rect 12684 8258 12740 8260
rect 12684 8206 12686 8258
rect 12686 8206 12738 8258
rect 12738 8206 12740 8258
rect 12684 8204 12740 8206
rect 13132 8316 13188 8372
rect 13020 8146 13076 8148
rect 13020 8094 13022 8146
rect 13022 8094 13074 8146
rect 13074 8094 13076 8146
rect 13020 8092 13076 8094
rect 12796 7756 12852 7812
rect 13020 7868 13076 7924
rect 12236 7308 12292 7364
rect 12684 7362 12740 7364
rect 12684 7310 12686 7362
rect 12686 7310 12738 7362
rect 12738 7310 12740 7362
rect 12684 7308 12740 7310
rect 12348 7196 12404 7252
rect 12684 7084 12740 7140
rect 12124 5740 12180 5796
rect 13020 7698 13076 7700
rect 13020 7646 13022 7698
rect 13022 7646 13074 7698
rect 13074 7646 13076 7698
rect 13020 7644 13076 7646
rect 13020 7084 13076 7140
rect 13244 7308 13300 7364
rect 14364 9212 14420 9268
rect 13132 6636 13188 6692
rect 13356 7084 13412 7140
rect 12908 4562 12964 4564
rect 12908 4510 12910 4562
rect 12910 4510 12962 4562
rect 12962 4510 12964 4562
rect 12908 4508 12964 4510
rect 11900 4060 11956 4116
rect 12124 4060 12180 4116
rect 12012 3724 12068 3780
rect 11900 3388 11956 3444
rect 10108 3276 10164 3332
rect 12460 4060 12516 4116
rect 13132 3724 13188 3780
rect 13020 3612 13076 3668
rect 13356 5068 13412 5124
rect 13692 7308 13748 7364
rect 13580 6748 13636 6804
rect 13916 7196 13972 7252
rect 13916 6690 13972 6692
rect 13916 6638 13918 6690
rect 13918 6638 13970 6690
rect 13970 6638 13972 6690
rect 13916 6636 13972 6638
rect 14476 9100 14532 9156
rect 15036 10780 15092 10836
rect 15260 11116 15316 11172
rect 14812 10444 14868 10500
rect 15820 15202 15876 15204
rect 15820 15150 15822 15202
rect 15822 15150 15874 15202
rect 15874 15150 15876 15202
rect 15820 15148 15876 15150
rect 16044 13692 16100 13748
rect 15932 13468 15988 13524
rect 16828 15260 16884 15316
rect 18060 18450 18116 18452
rect 18060 18398 18062 18450
rect 18062 18398 18114 18450
rect 18114 18398 18116 18450
rect 18060 18396 18116 18398
rect 18172 17388 18228 17444
rect 18172 16828 18228 16884
rect 19292 26572 19348 26628
rect 19292 25452 19348 25508
rect 19404 23884 19460 23940
rect 19628 30828 19684 30884
rect 20076 29932 20132 29988
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19852 29036 19908 29092
rect 19628 28588 19684 28644
rect 21644 38108 21700 38164
rect 21868 38050 21924 38052
rect 21868 37998 21870 38050
rect 21870 37998 21922 38050
rect 21922 37998 21924 38050
rect 21868 37996 21924 37998
rect 21756 37826 21812 37828
rect 21756 37774 21758 37826
rect 21758 37774 21810 37826
rect 21810 37774 21812 37826
rect 21756 37772 21812 37774
rect 21868 36988 21924 37044
rect 24444 40236 24500 40292
rect 24668 39900 24724 39956
rect 23772 38946 23828 38948
rect 23772 38894 23774 38946
rect 23774 38894 23826 38946
rect 23826 38894 23828 38946
rect 23772 38892 23828 38894
rect 23324 38834 23380 38836
rect 23324 38782 23326 38834
rect 23326 38782 23378 38834
rect 23378 38782 23380 38834
rect 23324 38780 23380 38782
rect 23884 38834 23940 38836
rect 23884 38782 23886 38834
rect 23886 38782 23938 38834
rect 23938 38782 23940 38834
rect 23884 38780 23940 38782
rect 24444 38780 24500 38836
rect 23996 38610 24052 38612
rect 23996 38558 23998 38610
rect 23998 38558 24050 38610
rect 24050 38558 24052 38610
rect 23996 38556 24052 38558
rect 21980 36540 22036 36596
rect 22764 38162 22820 38164
rect 22764 38110 22766 38162
rect 22766 38110 22818 38162
rect 22818 38110 22820 38162
rect 22764 38108 22820 38110
rect 22204 37772 22260 37828
rect 22428 38050 22484 38052
rect 22428 37998 22430 38050
rect 22430 37998 22482 38050
rect 22482 37998 22484 38050
rect 22428 37996 22484 37998
rect 22540 37884 22596 37940
rect 22540 36876 22596 36932
rect 22204 36652 22260 36708
rect 22316 36540 22372 36596
rect 21644 36258 21700 36260
rect 21644 36206 21646 36258
rect 21646 36206 21698 36258
rect 21698 36206 21700 36258
rect 21644 36204 21700 36206
rect 23100 37266 23156 37268
rect 23100 37214 23102 37266
rect 23102 37214 23154 37266
rect 23154 37214 23156 37266
rect 23100 37212 23156 37214
rect 24668 37884 24724 37940
rect 23324 37212 23380 37268
rect 23884 37212 23940 37268
rect 23324 36876 23380 36932
rect 22652 36204 22708 36260
rect 22428 35980 22484 36036
rect 22092 35810 22148 35812
rect 22092 35758 22094 35810
rect 22094 35758 22146 35810
rect 22146 35758 22148 35810
rect 22092 35756 22148 35758
rect 21308 34972 21364 35028
rect 20972 34860 21028 34916
rect 20860 34188 20916 34244
rect 21644 35698 21700 35700
rect 21644 35646 21646 35698
rect 21646 35646 21698 35698
rect 21698 35646 21700 35698
rect 21644 35644 21700 35646
rect 21532 35196 21588 35252
rect 21644 35308 21700 35364
rect 21532 34188 21588 34244
rect 20860 32396 20916 32452
rect 22876 36652 22932 36708
rect 24556 37154 24612 37156
rect 24556 37102 24558 37154
rect 24558 37102 24610 37154
rect 24610 37102 24612 37154
rect 24556 37100 24612 37102
rect 24668 36876 24724 36932
rect 24108 36258 24164 36260
rect 24108 36206 24110 36258
rect 24110 36206 24162 36258
rect 24162 36206 24164 36258
rect 24108 36204 24164 36206
rect 22876 35922 22932 35924
rect 22876 35870 22878 35922
rect 22878 35870 22930 35922
rect 22930 35870 22932 35922
rect 22876 35868 22932 35870
rect 23996 35922 24052 35924
rect 23996 35870 23998 35922
rect 23998 35870 24050 35922
rect 24050 35870 24052 35922
rect 23996 35868 24052 35870
rect 22540 35698 22596 35700
rect 22540 35646 22542 35698
rect 22542 35646 22594 35698
rect 22594 35646 22596 35698
rect 22540 35644 22596 35646
rect 22316 35420 22372 35476
rect 21196 31948 21252 32004
rect 21868 31778 21924 31780
rect 21868 31726 21870 31778
rect 21870 31726 21922 31778
rect 21922 31726 21924 31778
rect 21868 31724 21924 31726
rect 20636 31388 20692 31444
rect 20748 31500 20804 31556
rect 20524 31276 20580 31332
rect 21532 31388 21588 31444
rect 21532 31164 21588 31220
rect 20300 31106 20356 31108
rect 20300 31054 20302 31106
rect 20302 31054 20354 31106
rect 20354 31054 20356 31106
rect 20300 31052 20356 31054
rect 21308 31052 21364 31108
rect 21196 29932 21252 29988
rect 19852 28364 19908 28420
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19628 27804 19684 27860
rect 19740 27244 19796 27300
rect 19852 27580 19908 27636
rect 20636 28642 20692 28644
rect 20636 28590 20638 28642
rect 20638 28590 20690 28642
rect 20690 28590 20692 28642
rect 20636 28588 20692 28590
rect 20748 28082 20804 28084
rect 20748 28030 20750 28082
rect 20750 28030 20802 28082
rect 20802 28030 20804 28082
rect 20748 28028 20804 28030
rect 20300 27804 20356 27860
rect 20076 27580 20132 27636
rect 20412 27132 20468 27188
rect 20748 27132 20804 27188
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20524 26460 20580 26516
rect 19628 25506 19684 25508
rect 19628 25454 19630 25506
rect 19630 25454 19682 25506
rect 19682 25454 19684 25506
rect 19628 25452 19684 25454
rect 20412 25506 20468 25508
rect 20412 25454 20414 25506
rect 20414 25454 20466 25506
rect 20466 25454 20468 25506
rect 20412 25452 20468 25454
rect 20748 25506 20804 25508
rect 20748 25454 20750 25506
rect 20750 25454 20802 25506
rect 20802 25454 20804 25506
rect 20748 25452 20804 25454
rect 20076 25228 20132 25284
rect 20300 25282 20356 25284
rect 20300 25230 20302 25282
rect 20302 25230 20354 25282
rect 20354 25230 20356 25282
rect 20300 25228 20356 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20748 24108 20804 24164
rect 21084 28924 21140 28980
rect 21420 30994 21476 30996
rect 21420 30942 21422 30994
rect 21422 30942 21474 30994
rect 21474 30942 21476 30994
rect 21420 30940 21476 30942
rect 21420 29708 21476 29764
rect 21084 28476 21140 28532
rect 21420 27132 21476 27188
rect 21420 26908 21476 26964
rect 20972 26514 21028 26516
rect 20972 26462 20974 26514
rect 20974 26462 21026 26514
rect 21026 26462 21028 26514
rect 20972 26460 21028 26462
rect 21308 26178 21364 26180
rect 21308 26126 21310 26178
rect 21310 26126 21362 26178
rect 21362 26126 21364 26178
rect 21308 26124 21364 26126
rect 21196 25340 21252 25396
rect 23548 35756 23604 35812
rect 23324 35308 23380 35364
rect 23660 35196 23716 35252
rect 22988 34914 23044 34916
rect 22988 34862 22990 34914
rect 22990 34862 23042 34914
rect 23042 34862 23044 34914
rect 22988 34860 23044 34862
rect 23548 34188 23604 34244
rect 23436 33516 23492 33572
rect 21644 29820 21700 29876
rect 21644 28588 21700 28644
rect 22428 29986 22484 29988
rect 22428 29934 22430 29986
rect 22430 29934 22482 29986
rect 22482 29934 22484 29986
rect 22428 29932 22484 29934
rect 22764 30828 22820 30884
rect 22652 29820 22708 29876
rect 21868 28700 21924 28756
rect 21756 27916 21812 27972
rect 22540 28588 22596 28644
rect 22428 28530 22484 28532
rect 22428 28478 22430 28530
rect 22430 28478 22482 28530
rect 22482 28478 22484 28530
rect 22428 28476 22484 28478
rect 23436 30380 23492 30436
rect 23212 30156 23268 30212
rect 22764 28252 22820 28308
rect 22988 28812 23044 28868
rect 21980 27244 22036 27300
rect 23100 28754 23156 28756
rect 23100 28702 23102 28754
rect 23102 28702 23154 28754
rect 23154 28702 23156 28754
rect 23100 28700 23156 28702
rect 23324 28588 23380 28644
rect 24556 36204 24612 36260
rect 24556 35980 24612 36036
rect 24332 33516 24388 33572
rect 23884 32060 23940 32116
rect 23884 31388 23940 31444
rect 24556 30940 24612 30996
rect 23548 30044 23604 30100
rect 24220 30156 24276 30212
rect 24220 29932 24276 29988
rect 23772 29820 23828 29876
rect 23884 29708 23940 29764
rect 30268 46172 30324 46228
rect 26572 45890 26628 45892
rect 26572 45838 26574 45890
rect 26574 45838 26626 45890
rect 26626 45838 26628 45890
rect 26572 45836 26628 45838
rect 27356 45890 27412 45892
rect 27356 45838 27358 45890
rect 27358 45838 27410 45890
rect 27410 45838 27412 45890
rect 27356 45836 27412 45838
rect 27580 45890 27636 45892
rect 27580 45838 27582 45890
rect 27582 45838 27634 45890
rect 27634 45838 27636 45890
rect 27580 45836 27636 45838
rect 26684 45778 26740 45780
rect 26684 45726 26686 45778
rect 26686 45726 26738 45778
rect 26738 45726 26740 45778
rect 26684 45724 26740 45726
rect 26460 45276 26516 45332
rect 26796 45276 26852 45332
rect 25564 45106 25620 45108
rect 25564 45054 25566 45106
rect 25566 45054 25618 45106
rect 25618 45054 25620 45106
rect 25564 45052 25620 45054
rect 25228 44380 25284 44436
rect 26684 44434 26740 44436
rect 26684 44382 26686 44434
rect 26686 44382 26738 44434
rect 26738 44382 26740 44434
rect 26684 44380 26740 44382
rect 25900 44044 25956 44100
rect 26908 45164 26964 45220
rect 27020 45052 27076 45108
rect 28028 45778 28084 45780
rect 28028 45726 28030 45778
rect 28030 45726 28082 45778
rect 28082 45726 28084 45778
rect 28028 45724 28084 45726
rect 28140 45330 28196 45332
rect 28140 45278 28142 45330
rect 28142 45278 28194 45330
rect 28194 45278 28196 45330
rect 28140 45276 28196 45278
rect 27916 45164 27972 45220
rect 27132 44044 27188 44100
rect 27916 44380 27972 44436
rect 25900 43148 25956 43204
rect 25452 42476 25508 42532
rect 25228 41970 25284 41972
rect 25228 41918 25230 41970
rect 25230 41918 25282 41970
rect 25282 41918 25284 41970
rect 25228 41916 25284 41918
rect 25228 41132 25284 41188
rect 25452 40514 25508 40516
rect 25452 40462 25454 40514
rect 25454 40462 25506 40514
rect 25506 40462 25508 40514
rect 25452 40460 25508 40462
rect 25340 38834 25396 38836
rect 25340 38782 25342 38834
rect 25342 38782 25394 38834
rect 25394 38782 25396 38834
rect 25340 38780 25396 38782
rect 25900 40796 25956 40852
rect 26908 42866 26964 42868
rect 26908 42814 26910 42866
rect 26910 42814 26962 42866
rect 26962 42814 26964 42866
rect 26908 42812 26964 42814
rect 26796 42700 26852 42756
rect 26908 42476 26964 42532
rect 26908 40684 26964 40740
rect 26348 40572 26404 40628
rect 25788 40290 25844 40292
rect 25788 40238 25790 40290
rect 25790 40238 25842 40290
rect 25842 40238 25844 40290
rect 25788 40236 25844 40238
rect 25676 39900 25732 39956
rect 25676 39340 25732 39396
rect 26572 39900 26628 39956
rect 26124 39004 26180 39060
rect 26236 39564 26292 39620
rect 25788 38946 25844 38948
rect 25788 38894 25790 38946
rect 25790 38894 25842 38946
rect 25842 38894 25844 38946
rect 25788 38892 25844 38894
rect 25564 38444 25620 38500
rect 26348 39340 26404 39396
rect 26796 40178 26852 40180
rect 26796 40126 26798 40178
rect 26798 40126 26850 40178
rect 26850 40126 26852 40178
rect 26796 40124 26852 40126
rect 26908 39058 26964 39060
rect 26908 39006 26910 39058
rect 26910 39006 26962 39058
rect 26962 39006 26964 39058
rect 26908 39004 26964 39006
rect 26796 38834 26852 38836
rect 26796 38782 26798 38834
rect 26798 38782 26850 38834
rect 26850 38782 26852 38834
rect 26796 38780 26852 38782
rect 25452 37938 25508 37940
rect 25452 37886 25454 37938
rect 25454 37886 25506 37938
rect 25506 37886 25508 37938
rect 25452 37884 25508 37886
rect 26348 37436 26404 37492
rect 25676 37378 25732 37380
rect 25676 37326 25678 37378
rect 25678 37326 25730 37378
rect 25730 37326 25732 37378
rect 25676 37324 25732 37326
rect 25228 37266 25284 37268
rect 25228 37214 25230 37266
rect 25230 37214 25282 37266
rect 25282 37214 25284 37266
rect 25228 37212 25284 37214
rect 25900 37266 25956 37268
rect 25900 37214 25902 37266
rect 25902 37214 25954 37266
rect 25954 37214 25956 37266
rect 25900 37212 25956 37214
rect 25564 37154 25620 37156
rect 25564 37102 25566 37154
rect 25566 37102 25618 37154
rect 25618 37102 25620 37154
rect 25564 37100 25620 37102
rect 26236 36876 26292 36932
rect 26796 37266 26852 37268
rect 26796 37214 26798 37266
rect 26798 37214 26850 37266
rect 26850 37214 26852 37266
rect 26796 37212 26852 37214
rect 27916 44044 27972 44100
rect 27356 43260 27412 43316
rect 27244 42812 27300 42868
rect 27580 43426 27636 43428
rect 27580 43374 27582 43426
rect 27582 43374 27634 43426
rect 27634 43374 27636 43426
rect 27580 43372 27636 43374
rect 27804 43538 27860 43540
rect 27804 43486 27806 43538
rect 27806 43486 27858 43538
rect 27858 43486 27860 43538
rect 27804 43484 27860 43486
rect 28924 45948 28980 46004
rect 28588 45106 28644 45108
rect 28588 45054 28590 45106
rect 28590 45054 28642 45106
rect 28642 45054 28644 45106
rect 28588 45052 28644 45054
rect 29148 45890 29204 45892
rect 29148 45838 29150 45890
rect 29150 45838 29202 45890
rect 29202 45838 29204 45890
rect 29148 45836 29204 45838
rect 30604 45890 30660 45892
rect 30604 45838 30606 45890
rect 30606 45838 30658 45890
rect 30658 45838 30660 45890
rect 30604 45836 30660 45838
rect 29932 45218 29988 45220
rect 29932 45166 29934 45218
rect 29934 45166 29986 45218
rect 29986 45166 29988 45218
rect 29932 45164 29988 45166
rect 30604 44940 30660 44996
rect 30940 45106 30996 45108
rect 30940 45054 30942 45106
rect 30942 45054 30994 45106
rect 30994 45054 30996 45106
rect 30940 45052 30996 45054
rect 30828 44492 30884 44548
rect 28252 44098 28308 44100
rect 28252 44046 28254 44098
rect 28254 44046 28306 44098
rect 28306 44046 28308 44098
rect 28252 44044 28308 44046
rect 27692 43148 27748 43204
rect 28028 43484 28084 43540
rect 27916 42924 27972 42980
rect 27916 42252 27972 42308
rect 27244 41858 27300 41860
rect 27244 41806 27246 41858
rect 27246 41806 27298 41858
rect 27298 41806 27300 41858
rect 27244 41804 27300 41806
rect 27916 42028 27972 42084
rect 27692 40684 27748 40740
rect 27580 40626 27636 40628
rect 27580 40574 27582 40626
rect 27582 40574 27634 40626
rect 27634 40574 27636 40626
rect 27580 40572 27636 40574
rect 28140 43372 28196 43428
rect 29932 43484 29988 43540
rect 29148 43426 29204 43428
rect 29148 43374 29150 43426
rect 29150 43374 29202 43426
rect 29202 43374 29204 43426
rect 29148 43372 29204 43374
rect 28364 43260 28420 43316
rect 28252 43036 28308 43092
rect 28476 42924 28532 42980
rect 29372 43314 29428 43316
rect 29372 43262 29374 43314
rect 29374 43262 29426 43314
rect 29426 43262 29428 43314
rect 29372 43260 29428 43262
rect 28924 43148 28980 43204
rect 28588 41244 28644 41300
rect 29036 43036 29092 43092
rect 29148 42978 29204 42980
rect 29148 42926 29150 42978
rect 29150 42926 29202 42978
rect 29202 42926 29204 42978
rect 29148 42924 29204 42926
rect 29260 42866 29316 42868
rect 29260 42814 29262 42866
rect 29262 42814 29314 42866
rect 29314 42814 29316 42866
rect 29260 42812 29316 42814
rect 30380 43260 30436 43316
rect 29484 41916 29540 41972
rect 29372 41244 29428 41300
rect 30604 42754 30660 42756
rect 30604 42702 30606 42754
rect 30606 42702 30658 42754
rect 30658 42702 30660 42754
rect 30604 42700 30660 42702
rect 30156 41692 30212 41748
rect 30492 42028 30548 42084
rect 28140 40684 28196 40740
rect 30156 40460 30212 40516
rect 27804 40124 27860 40180
rect 27356 39058 27412 39060
rect 27356 39006 27358 39058
rect 27358 39006 27410 39058
rect 27410 39006 27412 39058
rect 27356 39004 27412 39006
rect 27132 38556 27188 38612
rect 27132 37436 27188 37492
rect 27692 38668 27748 38724
rect 27692 37772 27748 37828
rect 28588 39452 28644 39508
rect 29372 39506 29428 39508
rect 29372 39454 29374 39506
rect 29374 39454 29426 39506
rect 29426 39454 29428 39506
rect 29372 39452 29428 39454
rect 28476 39340 28532 39396
rect 28140 38834 28196 38836
rect 28140 38782 28142 38834
rect 28142 38782 28194 38834
rect 28194 38782 28196 38834
rect 28140 38780 28196 38782
rect 29484 39340 29540 39396
rect 28588 38162 28644 38164
rect 28588 38110 28590 38162
rect 28590 38110 28642 38162
rect 28642 38110 28644 38162
rect 28588 38108 28644 38110
rect 28812 38220 28868 38276
rect 28476 37996 28532 38052
rect 28252 37884 28308 37940
rect 27916 37826 27972 37828
rect 27916 37774 27918 37826
rect 27918 37774 27970 37826
rect 27970 37774 27972 37826
rect 27916 37772 27972 37774
rect 27356 37212 27412 37268
rect 25228 34188 25284 34244
rect 25676 33068 25732 33124
rect 27356 35756 27412 35812
rect 27580 36988 27636 37044
rect 28252 37490 28308 37492
rect 28252 37438 28254 37490
rect 28254 37438 28306 37490
rect 28306 37438 28308 37490
rect 28252 37436 28308 37438
rect 29820 38892 29876 38948
rect 29596 38220 29652 38276
rect 29372 38050 29428 38052
rect 29372 37998 29374 38050
rect 29374 37998 29426 38050
rect 29426 37998 29428 38050
rect 29372 37996 29428 37998
rect 30044 39004 30100 39060
rect 29372 37772 29428 37828
rect 28028 35756 28084 35812
rect 27580 35698 27636 35700
rect 27580 35646 27582 35698
rect 27582 35646 27634 35698
rect 27634 35646 27636 35698
rect 27580 35644 27636 35646
rect 28588 35698 28644 35700
rect 28588 35646 28590 35698
rect 28590 35646 28642 35698
rect 28642 35646 28644 35698
rect 28588 35644 28644 35646
rect 29820 37436 29876 37492
rect 30156 37996 30212 38052
rect 29932 37100 29988 37156
rect 30828 43260 30884 43316
rect 31276 45836 31332 45892
rect 31276 44828 31332 44884
rect 31164 43036 31220 43092
rect 30716 42028 30772 42084
rect 30828 41020 30884 41076
rect 30828 39452 30884 39508
rect 32060 46172 32116 46228
rect 32172 46620 32228 46676
rect 31948 46002 32004 46004
rect 31948 45950 31950 46002
rect 31950 45950 32002 46002
rect 32002 45950 32004 46002
rect 31948 45948 32004 45950
rect 32956 45218 33012 45220
rect 32956 45166 32958 45218
rect 32958 45166 33010 45218
rect 33010 45166 33012 45218
rect 32956 45164 33012 45166
rect 33404 45164 33460 45220
rect 31724 44828 31780 44884
rect 32172 45106 32228 45108
rect 32172 45054 32174 45106
rect 32174 45054 32226 45106
rect 32226 45054 32228 45106
rect 32172 45052 32228 45054
rect 33628 45106 33684 45108
rect 33628 45054 33630 45106
rect 33630 45054 33682 45106
rect 33682 45054 33684 45106
rect 33628 45052 33684 45054
rect 32396 44994 32452 44996
rect 32396 44942 32398 44994
rect 32398 44942 32450 44994
rect 32450 44942 32452 44994
rect 32396 44940 32452 44942
rect 32508 44434 32564 44436
rect 32508 44382 32510 44434
rect 32510 44382 32562 44434
rect 32562 44382 32564 44434
rect 32508 44380 32564 44382
rect 31612 43538 31668 43540
rect 31612 43486 31614 43538
rect 31614 43486 31666 43538
rect 31666 43486 31668 43538
rect 31612 43484 31668 43486
rect 31836 43148 31892 43204
rect 31948 43372 32004 43428
rect 31052 42642 31108 42644
rect 31052 42590 31054 42642
rect 31054 42590 31106 42642
rect 31106 42590 31108 42642
rect 31052 42588 31108 42590
rect 31948 42754 32004 42756
rect 31948 42702 31950 42754
rect 31950 42702 32002 42754
rect 32002 42702 32004 42754
rect 31948 42700 32004 42702
rect 31164 42140 31220 42196
rect 31276 42028 31332 42084
rect 32620 43484 32676 43540
rect 31612 42530 31668 42532
rect 31612 42478 31614 42530
rect 31614 42478 31666 42530
rect 31666 42478 31668 42530
rect 31612 42476 31668 42478
rect 31612 42140 31668 42196
rect 31836 42140 31892 42196
rect 32284 43148 32340 43204
rect 32620 42754 32676 42756
rect 32620 42702 32622 42754
rect 32622 42702 32674 42754
rect 32674 42702 32676 42754
rect 32620 42700 32676 42702
rect 32172 42476 32228 42532
rect 31388 41970 31444 41972
rect 31388 41918 31390 41970
rect 31390 41918 31442 41970
rect 31442 41918 31444 41970
rect 31388 41916 31444 41918
rect 31836 41132 31892 41188
rect 32732 42530 32788 42532
rect 32732 42478 32734 42530
rect 32734 42478 32786 42530
rect 32786 42478 32788 42530
rect 32732 42476 32788 42478
rect 32396 42194 32452 42196
rect 32396 42142 32398 42194
rect 32398 42142 32450 42194
rect 32450 42142 32452 42194
rect 32396 42140 32452 42142
rect 33852 44828 33908 44884
rect 33740 44380 33796 44436
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 42364 47682 42420 47684
rect 42364 47630 42366 47682
rect 42366 47630 42418 47682
rect 42418 47630 42420 47682
rect 42364 47628 42420 47630
rect 40572 47570 40628 47572
rect 40572 47518 40574 47570
rect 40574 47518 40626 47570
rect 40626 47518 40628 47570
rect 40572 47516 40628 47518
rect 37772 47404 37828 47460
rect 35196 47180 35252 47236
rect 34188 46898 34244 46900
rect 34188 46846 34190 46898
rect 34190 46846 34242 46898
rect 34242 46846 34244 46898
rect 34188 46844 34244 46846
rect 35980 47234 36036 47236
rect 35980 47182 35982 47234
rect 35982 47182 36034 47234
rect 36034 47182 36036 47234
rect 35980 47180 36036 47182
rect 34412 46674 34468 46676
rect 34412 46622 34414 46674
rect 34414 46622 34466 46674
rect 34466 46622 34468 46674
rect 34412 46620 34468 46622
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 36876 47234 36932 47236
rect 36876 47182 36878 47234
rect 36878 47182 36930 47234
rect 36930 47182 36932 47234
rect 36876 47180 36932 47182
rect 35196 45164 35252 45220
rect 35084 45106 35140 45108
rect 35084 45054 35086 45106
rect 35086 45054 35138 45106
rect 35138 45054 35140 45106
rect 35084 45052 35140 45054
rect 32956 43708 33012 43764
rect 33180 44044 33236 44100
rect 33740 44098 33796 44100
rect 33740 44046 33742 44098
rect 33742 44046 33794 44098
rect 33794 44046 33796 44098
rect 33740 44044 33796 44046
rect 33740 43708 33796 43764
rect 33068 43426 33124 43428
rect 33068 43374 33070 43426
rect 33070 43374 33122 43426
rect 33122 43374 33124 43426
rect 33068 43372 33124 43374
rect 33516 43426 33572 43428
rect 33516 43374 33518 43426
rect 33518 43374 33570 43426
rect 33570 43374 33572 43426
rect 33516 43372 33572 43374
rect 34188 44940 34244 44996
rect 36204 45052 36260 45108
rect 35084 44828 35140 44884
rect 34748 44434 34804 44436
rect 34748 44382 34750 44434
rect 34750 44382 34802 44434
rect 34802 44382 34804 44434
rect 34748 44380 34804 44382
rect 33852 42754 33908 42756
rect 33852 42702 33854 42754
rect 33854 42702 33906 42754
rect 33906 42702 33908 42754
rect 33852 42700 33908 42702
rect 32956 42140 33012 42196
rect 33068 42476 33124 42532
rect 32396 41804 32452 41860
rect 32284 41020 32340 41076
rect 33068 40908 33124 40964
rect 32172 39058 32228 39060
rect 32172 39006 32174 39058
rect 32174 39006 32226 39058
rect 32226 39006 32228 39058
rect 32172 39004 32228 39006
rect 32284 39340 32340 39396
rect 30604 38556 30660 38612
rect 30604 38050 30660 38052
rect 30604 37998 30606 38050
rect 30606 37998 30658 38050
rect 30658 37998 30660 38050
rect 30604 37996 30660 37998
rect 30492 37772 30548 37828
rect 30380 37324 30436 37380
rect 30156 37212 30212 37268
rect 30492 37100 30548 37156
rect 29484 36540 29540 36596
rect 29372 35756 29428 35812
rect 30380 36428 30436 36484
rect 29148 35644 29204 35700
rect 30268 35698 30324 35700
rect 30268 35646 30270 35698
rect 30270 35646 30322 35698
rect 30322 35646 30324 35698
rect 30268 35644 30324 35646
rect 27468 35138 27524 35140
rect 27468 35086 27470 35138
rect 27470 35086 27522 35138
rect 27522 35086 27524 35138
rect 27468 35084 27524 35086
rect 25788 31836 25844 31892
rect 24668 30044 24724 30100
rect 24780 29932 24836 29988
rect 25004 29986 25060 29988
rect 25004 29934 25006 29986
rect 25006 29934 25058 29986
rect 25058 29934 25060 29986
rect 25004 29932 25060 29934
rect 24668 29372 24724 29428
rect 25564 29484 25620 29540
rect 22988 26796 23044 26852
rect 23212 28140 23268 28196
rect 23212 26460 23268 26516
rect 21756 25564 21812 25620
rect 22092 26124 22148 26180
rect 23100 26124 23156 26180
rect 22204 25788 22260 25844
rect 21980 25506 22036 25508
rect 21980 25454 21982 25506
rect 21982 25454 22034 25506
rect 22034 25454 22036 25506
rect 21980 25452 22036 25454
rect 21308 24892 21364 24948
rect 21420 25004 21476 25060
rect 20860 23996 20916 24052
rect 19180 23100 19236 23156
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18508 23042 18564 23044
rect 18508 22990 18510 23042
rect 18510 22990 18562 23042
rect 18562 22990 18564 23042
rect 18508 22988 18564 22990
rect 19404 22876 19460 22932
rect 18956 21756 19012 21812
rect 19068 22204 19124 22260
rect 18396 21420 18452 21476
rect 19404 21644 19460 21700
rect 19516 22092 19572 22148
rect 20188 22652 20244 22708
rect 20636 22652 20692 22708
rect 20076 22092 20132 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20972 23042 21028 23044
rect 20972 22990 20974 23042
rect 20974 22990 21026 23042
rect 21026 22990 21028 23042
rect 20972 22988 21028 22990
rect 21196 23100 21252 23156
rect 21532 24220 21588 24276
rect 21644 25116 21700 25172
rect 21532 24050 21588 24052
rect 21532 23998 21534 24050
rect 21534 23998 21586 24050
rect 21586 23998 21588 24050
rect 21532 23996 21588 23998
rect 21644 22652 21700 22708
rect 22540 25340 22596 25396
rect 24108 28252 24164 28308
rect 23884 27746 23940 27748
rect 23884 27694 23886 27746
rect 23886 27694 23938 27746
rect 23938 27694 23940 27746
rect 23884 27692 23940 27694
rect 23436 26962 23492 26964
rect 23436 26910 23438 26962
rect 23438 26910 23490 26962
rect 23490 26910 23492 26962
rect 23436 26908 23492 26910
rect 24780 27804 24836 27860
rect 24892 27580 24948 27636
rect 23884 26178 23940 26180
rect 23884 26126 23886 26178
rect 23886 26126 23938 26178
rect 23938 26126 23940 26178
rect 23884 26124 23940 26126
rect 23996 26012 24052 26068
rect 22876 25452 22932 25508
rect 22428 25282 22484 25284
rect 22428 25230 22430 25282
rect 22430 25230 22482 25282
rect 22482 25230 22484 25282
rect 22428 25228 22484 25230
rect 22652 25228 22708 25284
rect 22428 25004 22484 25060
rect 22764 24946 22820 24948
rect 22764 24894 22766 24946
rect 22766 24894 22818 24946
rect 22818 24894 22820 24946
rect 22764 24892 22820 24894
rect 23436 25564 23492 25620
rect 22988 25394 23044 25396
rect 22988 25342 22990 25394
rect 22990 25342 23042 25394
rect 23042 25342 23044 25394
rect 22988 25340 23044 25342
rect 22876 23884 22932 23940
rect 21084 22204 21140 22260
rect 20860 21810 20916 21812
rect 20860 21758 20862 21810
rect 20862 21758 20914 21810
rect 20914 21758 20916 21810
rect 20860 21756 20916 21758
rect 21196 21698 21252 21700
rect 21196 21646 21198 21698
rect 21198 21646 21250 21698
rect 21250 21646 21252 21698
rect 21196 21644 21252 21646
rect 19628 21420 19684 21476
rect 20412 21420 20468 21476
rect 19180 21084 19236 21140
rect 19740 20802 19796 20804
rect 19740 20750 19742 20802
rect 19742 20750 19794 20802
rect 19794 20750 19796 20802
rect 19740 20748 19796 20750
rect 19628 20636 19684 20692
rect 20748 20690 20804 20692
rect 20748 20638 20750 20690
rect 20750 20638 20802 20690
rect 20802 20638 20804 20690
rect 20748 20636 20804 20638
rect 19516 20300 19572 20356
rect 18396 19346 18452 19348
rect 18396 19294 18398 19346
rect 18398 19294 18450 19346
rect 18450 19294 18452 19346
rect 18396 19292 18452 19294
rect 18732 19180 18788 19236
rect 18732 18620 18788 18676
rect 18620 18284 18676 18340
rect 18508 17948 18564 18004
rect 18060 15314 18116 15316
rect 18060 15262 18062 15314
rect 18062 15262 18114 15314
rect 18114 15262 18116 15314
rect 18060 15260 18116 15262
rect 17948 15148 18004 15204
rect 19068 19404 19124 19460
rect 19180 18562 19236 18564
rect 19180 18510 19182 18562
rect 19182 18510 19234 18562
rect 19234 18510 19236 18562
rect 19180 18508 19236 18510
rect 19404 18674 19460 18676
rect 19404 18622 19406 18674
rect 19406 18622 19458 18674
rect 19458 18622 19460 18674
rect 19404 18620 19460 18622
rect 19068 18060 19124 18116
rect 19404 17778 19460 17780
rect 19404 17726 19406 17778
rect 19406 17726 19458 17778
rect 19458 17726 19460 17778
rect 19404 17724 19460 17726
rect 18956 17052 19012 17108
rect 18620 16156 18676 16212
rect 18844 16268 18900 16324
rect 18396 15484 18452 15540
rect 17948 14812 18004 14868
rect 18172 14306 18228 14308
rect 18172 14254 18174 14306
rect 18174 14254 18226 14306
rect 18226 14254 18228 14306
rect 18172 14252 18228 14254
rect 16268 13468 16324 13524
rect 16604 13580 16660 13636
rect 16380 12908 16436 12964
rect 16380 12348 16436 12404
rect 17612 13746 17668 13748
rect 17612 13694 17614 13746
rect 17614 13694 17666 13746
rect 17666 13694 17668 13746
rect 17612 13692 17668 13694
rect 17500 13634 17556 13636
rect 17500 13582 17502 13634
rect 17502 13582 17554 13634
rect 17554 13582 17556 13634
rect 17500 13580 17556 13582
rect 17276 13468 17332 13524
rect 16828 12908 16884 12964
rect 17724 12796 17780 12852
rect 16716 12178 16772 12180
rect 16716 12126 16718 12178
rect 16718 12126 16770 12178
rect 16770 12126 16772 12178
rect 16716 12124 16772 12126
rect 16380 11676 16436 11732
rect 16716 10834 16772 10836
rect 16716 10782 16718 10834
rect 16718 10782 16770 10834
rect 16770 10782 16772 10834
rect 16716 10780 16772 10782
rect 17388 12178 17444 12180
rect 17388 12126 17390 12178
rect 17390 12126 17442 12178
rect 17442 12126 17444 12178
rect 17388 12124 17444 12126
rect 15372 10556 15428 10612
rect 16156 10610 16212 10612
rect 16156 10558 16158 10610
rect 16158 10558 16210 10610
rect 16210 10558 16212 10610
rect 16156 10556 16212 10558
rect 15932 10498 15988 10500
rect 15932 10446 15934 10498
rect 15934 10446 15986 10498
rect 15986 10446 15988 10498
rect 15932 10444 15988 10446
rect 15596 9826 15652 9828
rect 15596 9774 15598 9826
rect 15598 9774 15650 9826
rect 15650 9774 15652 9826
rect 15596 9772 15652 9774
rect 16604 10444 16660 10500
rect 16940 11564 16996 11620
rect 16044 9996 16100 10052
rect 16044 9266 16100 9268
rect 16044 9214 16046 9266
rect 16046 9214 16098 9266
rect 16098 9214 16100 9266
rect 16044 9212 16100 9214
rect 14812 8428 14868 8484
rect 15036 8930 15092 8932
rect 15036 8878 15038 8930
rect 15038 8878 15090 8930
rect 15090 8878 15092 8930
rect 15036 8876 15092 8878
rect 15036 8316 15092 8372
rect 14700 7420 14756 7476
rect 14700 7084 14756 7140
rect 14588 6690 14644 6692
rect 14588 6638 14590 6690
rect 14590 6638 14642 6690
rect 14642 6638 14644 6690
rect 14588 6636 14644 6638
rect 15372 8316 15428 8372
rect 16492 8316 16548 8372
rect 16156 8258 16212 8260
rect 16156 8206 16158 8258
rect 16158 8206 16210 8258
rect 16210 8206 16212 8258
rect 16156 8204 16212 8206
rect 16716 8316 16772 8372
rect 16492 7980 16548 8036
rect 18060 13692 18116 13748
rect 17724 10610 17780 10612
rect 17724 10558 17726 10610
rect 17726 10558 17778 10610
rect 17778 10558 17780 10610
rect 17724 10556 17780 10558
rect 18732 15260 18788 15316
rect 18620 13468 18676 13524
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 21308 21420 21364 21476
rect 21532 21308 21588 21364
rect 21756 22482 21812 22484
rect 21756 22430 21758 22482
rect 21758 22430 21810 22482
rect 21810 22430 21812 22482
rect 21756 22428 21812 22430
rect 22876 22764 22932 22820
rect 22764 22204 22820 22260
rect 21756 21586 21812 21588
rect 21756 21534 21758 21586
rect 21758 21534 21810 21586
rect 21810 21534 21812 21586
rect 21756 21532 21812 21534
rect 21756 21084 21812 21140
rect 22316 20914 22372 20916
rect 22316 20862 22318 20914
rect 22318 20862 22370 20914
rect 22370 20862 22372 20914
rect 22316 20860 22372 20862
rect 20076 19234 20132 19236
rect 20076 19182 20078 19234
rect 20078 19182 20130 19234
rect 20130 19182 20132 19234
rect 20076 19180 20132 19182
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19740 18450 19796 18452
rect 19740 18398 19742 18450
rect 19742 18398 19794 18450
rect 19794 18398 19796 18450
rect 19740 18396 19796 18398
rect 20076 18226 20132 18228
rect 20076 18174 20078 18226
rect 20078 18174 20130 18226
rect 20130 18174 20132 18226
rect 20076 18172 20132 18174
rect 20188 17948 20244 18004
rect 20412 18284 20468 18340
rect 20188 17666 20244 17668
rect 20188 17614 20190 17666
rect 20190 17614 20242 17666
rect 20242 17614 20244 17666
rect 20188 17612 20244 17614
rect 21980 20018 22036 20020
rect 21980 19966 21982 20018
rect 21982 19966 22034 20018
rect 22034 19966 22036 20018
rect 21980 19964 22036 19966
rect 21308 19292 21364 19348
rect 21756 19292 21812 19348
rect 21532 19234 21588 19236
rect 21532 19182 21534 19234
rect 21534 19182 21586 19234
rect 21586 19182 21588 19234
rect 21532 19180 21588 19182
rect 21308 17948 21364 18004
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19964 16716 20020 16772
rect 22652 21420 22708 21476
rect 22876 20860 22932 20916
rect 23996 25506 24052 25508
rect 23996 25454 23998 25506
rect 23998 25454 24050 25506
rect 24050 25454 24052 25506
rect 23996 25452 24052 25454
rect 23772 25394 23828 25396
rect 23772 25342 23774 25394
rect 23774 25342 23826 25394
rect 23826 25342 23828 25394
rect 23772 25340 23828 25342
rect 23660 25282 23716 25284
rect 23660 25230 23662 25282
rect 23662 25230 23714 25282
rect 23714 25230 23716 25282
rect 23660 25228 23716 25230
rect 24444 25282 24500 25284
rect 24444 25230 24446 25282
rect 24446 25230 24498 25282
rect 24498 25230 24500 25282
rect 24444 25228 24500 25230
rect 23884 24722 23940 24724
rect 23884 24670 23886 24722
rect 23886 24670 23938 24722
rect 23938 24670 23940 24722
rect 23884 24668 23940 24670
rect 23436 24220 23492 24276
rect 23772 22428 23828 22484
rect 23548 21756 23604 21812
rect 23324 21308 23380 21364
rect 22988 21196 23044 21252
rect 23212 21196 23268 21252
rect 22316 19180 22372 19236
rect 22428 19404 22484 19460
rect 22764 19068 22820 19124
rect 23212 20636 23268 20692
rect 23100 20076 23156 20132
rect 22988 19516 23044 19572
rect 21756 17612 21812 17668
rect 21308 17554 21364 17556
rect 21308 17502 21310 17554
rect 21310 17502 21362 17554
rect 21362 17502 21364 17554
rect 21308 17500 21364 17502
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19404 15538 19460 15540
rect 19404 15486 19406 15538
rect 19406 15486 19458 15538
rect 19458 15486 19460 15538
rect 19404 15484 19460 15486
rect 18956 14924 19012 14980
rect 20524 15538 20580 15540
rect 20524 15486 20526 15538
rect 20526 15486 20578 15538
rect 20578 15486 20580 15538
rect 20524 15484 20580 15486
rect 20748 15036 20804 15092
rect 20412 14924 20468 14980
rect 19292 13692 19348 13748
rect 19516 14306 19572 14308
rect 19516 14254 19518 14306
rect 19518 14254 19570 14306
rect 19570 14254 19572 14306
rect 19516 14252 19572 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18956 13580 19012 13636
rect 18732 13132 18788 13188
rect 19628 13634 19684 13636
rect 19628 13582 19630 13634
rect 19630 13582 19682 13634
rect 19682 13582 19684 13634
rect 19628 13580 19684 13582
rect 19740 13020 19796 13076
rect 19516 12684 19572 12740
rect 20748 13580 20804 13636
rect 20636 13074 20692 13076
rect 20636 13022 20638 13074
rect 20638 13022 20690 13074
rect 20690 13022 20692 13074
rect 20636 13020 20692 13022
rect 20412 12796 20468 12852
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 18844 12066 18900 12068
rect 18844 12014 18846 12066
rect 18846 12014 18898 12066
rect 18898 12014 18900 12066
rect 18844 12012 18900 12014
rect 18284 11452 18340 11508
rect 18396 11900 18452 11956
rect 19068 11954 19124 11956
rect 19068 11902 19070 11954
rect 19070 11902 19122 11954
rect 19122 11902 19124 11954
rect 19068 11900 19124 11902
rect 19180 11506 19236 11508
rect 19180 11454 19182 11506
rect 19182 11454 19234 11506
rect 19234 11454 19236 11506
rect 19180 11452 19236 11454
rect 19964 11394 20020 11396
rect 19964 11342 19966 11394
rect 19966 11342 20018 11394
rect 20018 11342 20020 11394
rect 19964 11340 20020 11342
rect 18284 9996 18340 10052
rect 16940 9772 16996 9828
rect 17164 9100 17220 9156
rect 16940 8370 16996 8372
rect 16940 8318 16942 8370
rect 16942 8318 16994 8370
rect 16994 8318 16996 8370
rect 16940 8316 16996 8318
rect 16828 8204 16884 8260
rect 15596 7868 15652 7924
rect 16940 8092 16996 8148
rect 16828 7308 16884 7364
rect 15484 7196 15540 7252
rect 15596 7084 15652 7140
rect 13916 5740 13972 5796
rect 13692 5122 13748 5124
rect 13692 5070 13694 5122
rect 13694 5070 13746 5122
rect 13746 5070 13748 5122
rect 13692 5068 13748 5070
rect 15596 6076 15652 6132
rect 16268 7084 16324 7140
rect 16156 5964 16212 6020
rect 16828 6636 16884 6692
rect 15596 4844 15652 4900
rect 16716 4284 16772 4340
rect 16940 5906 16996 5908
rect 16940 5854 16942 5906
rect 16942 5854 16994 5906
rect 16994 5854 16996 5906
rect 16940 5852 16996 5854
rect 13692 3500 13748 3556
rect 12236 2940 12292 2996
rect 16380 3554 16436 3556
rect 16380 3502 16382 3554
rect 16382 3502 16434 3554
rect 16434 3502 16436 3554
rect 16380 3500 16436 3502
rect 17388 7084 17444 7140
rect 18284 9548 18340 9604
rect 18844 9996 18900 10052
rect 20300 11340 20356 11396
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 20412 11788 20468 11844
rect 21196 16156 21252 16212
rect 21532 17442 21588 17444
rect 21532 17390 21534 17442
rect 21534 17390 21586 17442
rect 21586 17390 21588 17442
rect 21532 17388 21588 17390
rect 22316 18060 22372 18116
rect 22204 17778 22260 17780
rect 22204 17726 22206 17778
rect 22206 17726 22258 17778
rect 22258 17726 22260 17778
rect 22204 17724 22260 17726
rect 22092 17666 22148 17668
rect 22092 17614 22094 17666
rect 22094 17614 22146 17666
rect 22146 17614 22148 17666
rect 22092 17612 22148 17614
rect 21644 16882 21700 16884
rect 21644 16830 21646 16882
rect 21646 16830 21698 16882
rect 21698 16830 21700 16882
rect 21644 16828 21700 16830
rect 21532 16770 21588 16772
rect 21532 16718 21534 16770
rect 21534 16718 21586 16770
rect 21586 16718 21588 16770
rect 21532 16716 21588 16718
rect 21532 16098 21588 16100
rect 21532 16046 21534 16098
rect 21534 16046 21586 16098
rect 21586 16046 21588 16098
rect 21532 16044 21588 16046
rect 22540 16156 22596 16212
rect 22540 15986 22596 15988
rect 22540 15934 22542 15986
rect 22542 15934 22594 15986
rect 22594 15934 22596 15986
rect 22540 15932 22596 15934
rect 22204 15874 22260 15876
rect 22204 15822 22206 15874
rect 22206 15822 22258 15874
rect 22258 15822 22260 15874
rect 22204 15820 22260 15822
rect 21084 15036 21140 15092
rect 22316 15314 22372 15316
rect 22316 15262 22318 15314
rect 22318 15262 22370 15314
rect 22370 15262 22372 15314
rect 22316 15260 22372 15262
rect 22204 15148 22260 15204
rect 21644 15036 21700 15092
rect 21644 14364 21700 14420
rect 23436 21084 23492 21140
rect 23436 19852 23492 19908
rect 23436 19516 23492 19572
rect 23660 20076 23716 20132
rect 24220 22428 24276 22484
rect 23884 22258 23940 22260
rect 23884 22206 23886 22258
rect 23886 22206 23938 22258
rect 23938 22206 23940 22258
rect 23884 22204 23940 22206
rect 23996 21532 24052 21588
rect 24780 25676 24836 25732
rect 24780 23884 24836 23940
rect 24668 22428 24724 22484
rect 24892 21868 24948 21924
rect 24556 21532 24612 21588
rect 24556 20914 24612 20916
rect 24556 20862 24558 20914
rect 24558 20862 24610 20914
rect 24610 20862 24612 20914
rect 24556 20860 24612 20862
rect 23996 20242 24052 20244
rect 23996 20190 23998 20242
rect 23998 20190 24050 20242
rect 24050 20190 24052 20242
rect 23996 20188 24052 20190
rect 25228 29426 25284 29428
rect 25228 29374 25230 29426
rect 25230 29374 25282 29426
rect 25282 29374 25284 29426
rect 25228 29372 25284 29374
rect 25452 28812 25508 28868
rect 25340 28588 25396 28644
rect 27244 34076 27300 34132
rect 28364 35308 28420 35364
rect 29260 35308 29316 35364
rect 29148 35196 29204 35252
rect 28028 34300 28084 34356
rect 27580 33516 27636 33572
rect 26796 33122 26852 33124
rect 26796 33070 26798 33122
rect 26798 33070 26850 33122
rect 26850 33070 26852 33122
rect 26796 33068 26852 33070
rect 26908 32674 26964 32676
rect 26908 32622 26910 32674
rect 26910 32622 26962 32674
rect 26962 32622 26964 32674
rect 26908 32620 26964 32622
rect 27132 32508 27188 32564
rect 26124 31164 26180 31220
rect 25228 27746 25284 27748
rect 25228 27694 25230 27746
rect 25230 27694 25282 27746
rect 25282 27694 25284 27746
rect 25228 27692 25284 27694
rect 25452 27692 25508 27748
rect 26236 30210 26292 30212
rect 26236 30158 26238 30210
rect 26238 30158 26290 30210
rect 26290 30158 26292 30210
rect 26236 30156 26292 30158
rect 27804 34076 27860 34132
rect 27468 31948 27524 32004
rect 28700 35084 28756 35140
rect 28588 34354 28644 34356
rect 28588 34302 28590 34354
rect 28590 34302 28642 34354
rect 28642 34302 28644 34354
rect 28588 34300 28644 34302
rect 28364 34130 28420 34132
rect 28364 34078 28366 34130
rect 28366 34078 28418 34130
rect 28418 34078 28420 34130
rect 28364 34076 28420 34078
rect 27916 32732 27972 32788
rect 28700 32786 28756 32788
rect 28700 32734 28702 32786
rect 28702 32734 28754 32786
rect 28754 32734 28756 32786
rect 28700 32732 28756 32734
rect 28364 32620 28420 32676
rect 28028 31948 28084 32004
rect 27916 31666 27972 31668
rect 27916 31614 27918 31666
rect 27918 31614 27970 31666
rect 27970 31614 27972 31666
rect 27916 31612 27972 31614
rect 27692 30380 27748 30436
rect 27468 30268 27524 30324
rect 27356 30210 27412 30212
rect 27356 30158 27358 30210
rect 27358 30158 27410 30210
rect 27410 30158 27412 30210
rect 27356 30156 27412 30158
rect 28140 30434 28196 30436
rect 28140 30382 28142 30434
rect 28142 30382 28194 30434
rect 28194 30382 28196 30434
rect 28140 30380 28196 30382
rect 26348 28700 26404 28756
rect 26348 27580 26404 27636
rect 25228 25900 25284 25956
rect 25116 25452 25172 25508
rect 25228 24722 25284 24724
rect 25228 24670 25230 24722
rect 25230 24670 25282 24722
rect 25282 24670 25284 24722
rect 25228 24668 25284 24670
rect 25452 26236 25508 26292
rect 25788 26124 25844 26180
rect 25340 22428 25396 22484
rect 25228 20524 25284 20580
rect 23884 19964 23940 20020
rect 23548 19068 23604 19124
rect 23212 17948 23268 18004
rect 23324 17724 23380 17780
rect 23660 18732 23716 18788
rect 23436 17554 23492 17556
rect 23436 17502 23438 17554
rect 23438 17502 23490 17554
rect 23490 17502 23492 17554
rect 23436 17500 23492 17502
rect 24220 20076 24276 20132
rect 24668 20130 24724 20132
rect 24668 20078 24670 20130
rect 24670 20078 24722 20130
rect 24722 20078 24724 20130
rect 24668 20076 24724 20078
rect 24332 19292 24388 19348
rect 25004 19404 25060 19460
rect 24444 19010 24500 19012
rect 24444 18958 24446 19010
rect 24446 18958 24498 19010
rect 24498 18958 24500 19010
rect 24444 18956 24500 18958
rect 24332 18844 24388 18900
rect 24220 18172 24276 18228
rect 23884 17836 23940 17892
rect 24556 17948 24612 18004
rect 24892 17724 24948 17780
rect 24780 17666 24836 17668
rect 24780 17614 24782 17666
rect 24782 17614 24834 17666
rect 24834 17614 24836 17666
rect 24780 17612 24836 17614
rect 24444 17052 24500 17108
rect 24668 17052 24724 17108
rect 24556 16044 24612 16100
rect 23548 15932 23604 15988
rect 23660 14418 23716 14420
rect 23660 14366 23662 14418
rect 23662 14366 23714 14418
rect 23714 14366 23716 14418
rect 23660 14364 23716 14366
rect 22652 13916 22708 13972
rect 21084 13244 21140 13300
rect 21756 13580 21812 13636
rect 21644 12684 21700 12740
rect 21084 12460 21140 12516
rect 20860 11676 20916 11732
rect 20860 11282 20916 11284
rect 20860 11230 20862 11282
rect 20862 11230 20914 11282
rect 20914 11230 20916 11282
rect 20860 11228 20916 11230
rect 20972 10834 21028 10836
rect 20972 10782 20974 10834
rect 20974 10782 21026 10834
rect 21026 10782 21028 10834
rect 20972 10780 21028 10782
rect 20300 10050 20356 10052
rect 20300 9998 20302 10050
rect 20302 9998 20354 10050
rect 20354 9998 20356 10050
rect 20300 9996 20356 9998
rect 19516 9660 19572 9716
rect 20636 9602 20692 9604
rect 20636 9550 20638 9602
rect 20638 9550 20690 9602
rect 20690 9550 20692 9602
rect 20636 9548 20692 9550
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20188 9436 20244 9492
rect 20636 9154 20692 9156
rect 20636 9102 20638 9154
rect 20638 9102 20690 9154
rect 20690 9102 20692 9154
rect 20636 9100 20692 9102
rect 20076 8930 20132 8932
rect 20076 8878 20078 8930
rect 20078 8878 20130 8930
rect 20130 8878 20132 8930
rect 20076 8876 20132 8878
rect 17948 8092 18004 8148
rect 17724 7362 17780 7364
rect 17724 7310 17726 7362
rect 17726 7310 17778 7362
rect 17778 7310 17780 7362
rect 17724 7308 17780 7310
rect 17724 6300 17780 6356
rect 17836 6524 17892 6580
rect 17724 6130 17780 6132
rect 17724 6078 17726 6130
rect 17726 6078 17778 6130
rect 17778 6078 17780 6130
rect 17724 6076 17780 6078
rect 18508 6578 18564 6580
rect 18508 6526 18510 6578
rect 18510 6526 18562 6578
rect 18562 6526 18564 6578
rect 18508 6524 18564 6526
rect 18508 6300 18564 6356
rect 17164 5740 17220 5796
rect 18620 5906 18676 5908
rect 18620 5854 18622 5906
rect 18622 5854 18674 5906
rect 18674 5854 18676 5906
rect 18620 5852 18676 5854
rect 20188 8316 20244 8372
rect 19180 7420 19236 7476
rect 18956 5964 19012 6020
rect 19852 7980 19908 8036
rect 20748 8876 20804 8932
rect 20524 8540 20580 8596
rect 20636 8204 20692 8260
rect 20412 7980 20468 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20636 6802 20692 6804
rect 20636 6750 20638 6802
rect 20638 6750 20690 6802
rect 20690 6750 20692 6802
rect 20636 6748 20692 6750
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19404 5964 19460 6020
rect 18620 5068 18676 5124
rect 17500 4338 17556 4340
rect 17500 4286 17502 4338
rect 17502 4286 17554 4338
rect 17554 4286 17556 4338
rect 17500 4284 17556 4286
rect 17500 4060 17556 4116
rect 18508 4114 18564 4116
rect 18508 4062 18510 4114
rect 18510 4062 18562 4114
rect 18562 4062 18564 4114
rect 18508 4060 18564 4062
rect 20188 5964 20244 6020
rect 20076 5906 20132 5908
rect 20076 5854 20078 5906
rect 20078 5854 20130 5906
rect 20130 5854 20132 5906
rect 20076 5852 20132 5854
rect 19740 5122 19796 5124
rect 19740 5070 19742 5122
rect 19742 5070 19794 5122
rect 19794 5070 19796 5122
rect 19740 5068 19796 5070
rect 21308 10610 21364 10612
rect 21308 10558 21310 10610
rect 21310 10558 21362 10610
rect 21362 10558 21364 10610
rect 21308 10556 21364 10558
rect 22764 13692 22820 13748
rect 21980 12850 22036 12852
rect 21980 12798 21982 12850
rect 21982 12798 22034 12850
rect 22034 12798 22036 12850
rect 21980 12796 22036 12798
rect 22764 12908 22820 12964
rect 22876 12850 22932 12852
rect 22876 12798 22878 12850
rect 22878 12798 22930 12850
rect 22930 12798 22932 12850
rect 22876 12796 22932 12798
rect 23212 12796 23268 12852
rect 22652 12684 22708 12740
rect 23100 12572 23156 12628
rect 22092 11788 22148 11844
rect 21644 11282 21700 11284
rect 21644 11230 21646 11282
rect 21646 11230 21698 11282
rect 21698 11230 21700 11282
rect 21644 11228 21700 11230
rect 21980 11004 22036 11060
rect 22428 12012 22484 12068
rect 21980 9826 22036 9828
rect 21980 9774 21982 9826
rect 21982 9774 22034 9826
rect 22034 9774 22036 9826
rect 21980 9772 22036 9774
rect 21644 9660 21700 9716
rect 22428 9436 22484 9492
rect 21308 9212 21364 9268
rect 22988 11228 23044 11284
rect 22652 9772 22708 9828
rect 22876 9826 22932 9828
rect 22876 9774 22878 9826
rect 22878 9774 22930 9826
rect 22930 9774 22932 9826
rect 22876 9772 22932 9774
rect 22652 9602 22708 9604
rect 22652 9550 22654 9602
rect 22654 9550 22706 9602
rect 22706 9550 22708 9602
rect 22652 9548 22708 9550
rect 22316 9266 22372 9268
rect 22316 9214 22318 9266
rect 22318 9214 22370 9266
rect 22370 9214 22372 9266
rect 22316 9212 22372 9214
rect 23324 11676 23380 11732
rect 23212 9714 23268 9716
rect 23212 9662 23214 9714
rect 23214 9662 23266 9714
rect 23266 9662 23268 9714
rect 23212 9660 23268 9662
rect 22876 9324 22932 9380
rect 21420 8540 21476 8596
rect 21420 8258 21476 8260
rect 21420 8206 21422 8258
rect 21422 8206 21474 8258
rect 21474 8206 21476 8258
rect 21420 8204 21476 8206
rect 21308 8146 21364 8148
rect 21308 8094 21310 8146
rect 21310 8094 21362 8146
rect 21362 8094 21364 8146
rect 21308 8092 21364 8094
rect 21980 8652 22036 8708
rect 21644 7980 21700 8036
rect 20972 7868 21028 7924
rect 21756 7532 21812 7588
rect 21756 6748 21812 6804
rect 20972 6524 21028 6580
rect 21420 5964 21476 6020
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 21532 5180 21588 5236
rect 21196 4284 21252 4340
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22540 8988 22596 9044
rect 22204 8092 22260 8148
rect 22204 7644 22260 7700
rect 21980 6300 22036 6356
rect 21980 5404 22036 5460
rect 22428 5628 22484 5684
rect 22316 5234 22372 5236
rect 22316 5182 22318 5234
rect 22318 5182 22370 5234
rect 22370 5182 22372 5234
rect 22316 5180 22372 5182
rect 22428 5068 22484 5124
rect 21868 4396 21924 4452
rect 21756 3500 21812 3556
rect 22652 8764 22708 8820
rect 22876 8428 22932 8484
rect 23212 9100 23268 9156
rect 23996 13970 24052 13972
rect 23996 13918 23998 13970
rect 23998 13918 24050 13970
rect 24050 13918 24052 13970
rect 23996 13916 24052 13918
rect 24444 13916 24500 13972
rect 23772 13746 23828 13748
rect 23772 13694 23774 13746
rect 23774 13694 23826 13746
rect 23826 13694 23828 13746
rect 23772 13692 23828 13694
rect 24668 12796 24724 12852
rect 24444 12572 24500 12628
rect 24668 12236 24724 12292
rect 23996 11676 24052 11732
rect 24668 12066 24724 12068
rect 24668 12014 24670 12066
rect 24670 12014 24722 12066
rect 24722 12014 24724 12066
rect 24668 12012 24724 12014
rect 25676 22428 25732 22484
rect 26908 29932 26964 29988
rect 27132 29484 27188 29540
rect 26572 28364 26628 28420
rect 26908 28082 26964 28084
rect 26908 28030 26910 28082
rect 26910 28030 26962 28082
rect 26962 28030 26964 28082
rect 26908 28028 26964 28030
rect 25900 25788 25956 25844
rect 29260 34300 29316 34356
rect 29260 33292 29316 33348
rect 29708 35196 29764 35252
rect 29932 35084 29988 35140
rect 29484 34914 29540 34916
rect 29484 34862 29486 34914
rect 29486 34862 29538 34914
rect 29538 34862 29540 34914
rect 29484 34860 29540 34862
rect 30044 34914 30100 34916
rect 30044 34862 30046 34914
rect 30046 34862 30098 34914
rect 30098 34862 30100 34914
rect 30044 34860 30100 34862
rect 29484 34354 29540 34356
rect 29484 34302 29486 34354
rect 29486 34302 29538 34354
rect 29538 34302 29540 34354
rect 29484 34300 29540 34302
rect 29484 34076 29540 34132
rect 29820 34300 29876 34356
rect 29708 33404 29764 33460
rect 29596 33346 29652 33348
rect 29596 33294 29598 33346
rect 29598 33294 29650 33346
rect 29650 33294 29652 33346
rect 29596 33292 29652 33294
rect 30156 34300 30212 34356
rect 30268 35084 30324 35140
rect 30716 37324 30772 37380
rect 30604 36876 30660 36932
rect 30492 34300 30548 34356
rect 30604 34242 30660 34244
rect 30604 34190 30606 34242
rect 30606 34190 30658 34242
rect 30658 34190 30660 34242
rect 30604 34188 30660 34190
rect 29932 34130 29988 34132
rect 29932 34078 29934 34130
rect 29934 34078 29986 34130
rect 29986 34078 29988 34130
rect 29932 34076 29988 34078
rect 28924 32620 28980 32676
rect 28476 32284 28532 32340
rect 28476 31836 28532 31892
rect 28476 30044 28532 30100
rect 27916 29820 27972 29876
rect 27692 29484 27748 29540
rect 27356 27916 27412 27972
rect 27692 28642 27748 28644
rect 27692 28590 27694 28642
rect 27694 28590 27746 28642
rect 27746 28590 27748 28642
rect 27692 28588 27748 28590
rect 27468 27858 27524 27860
rect 27468 27806 27470 27858
rect 27470 27806 27522 27858
rect 27522 27806 27524 27858
rect 27468 27804 27524 27806
rect 27580 28418 27636 28420
rect 27580 28366 27582 28418
rect 27582 28366 27634 28418
rect 27634 28366 27636 28418
rect 27580 28364 27636 28366
rect 27804 28418 27860 28420
rect 27804 28366 27806 28418
rect 27806 28366 27858 28418
rect 27858 28366 27860 28418
rect 27804 28364 27860 28366
rect 27580 26908 27636 26964
rect 26796 26796 26852 26852
rect 27356 25900 27412 25956
rect 26684 25394 26740 25396
rect 26684 25342 26686 25394
rect 26686 25342 26738 25394
rect 26738 25342 26740 25394
rect 26684 25340 26740 25342
rect 27916 28028 27972 28084
rect 28700 30716 28756 30772
rect 28588 29932 28644 29988
rect 28252 26850 28308 26852
rect 28252 26798 28254 26850
rect 28254 26798 28306 26850
rect 28306 26798 28308 26850
rect 28252 26796 28308 26798
rect 28252 26348 28308 26404
rect 28028 26012 28084 26068
rect 27804 25564 27860 25620
rect 28140 25452 28196 25508
rect 27692 25394 27748 25396
rect 27692 25342 27694 25394
rect 27694 25342 27746 25394
rect 27746 25342 27748 25394
rect 27692 25340 27748 25342
rect 27804 25228 27860 25284
rect 26460 23884 26516 23940
rect 27020 23884 27076 23940
rect 25788 21756 25844 21812
rect 26236 23548 26292 23604
rect 26012 22258 26068 22260
rect 26012 22206 26014 22258
rect 26014 22206 26066 22258
rect 26066 22206 26068 22258
rect 26012 22204 26068 22206
rect 25788 20972 25844 21028
rect 25900 20860 25956 20916
rect 26124 21420 26180 21476
rect 26124 20748 26180 20804
rect 25452 19292 25508 19348
rect 25452 19068 25508 19124
rect 25340 18450 25396 18452
rect 25340 18398 25342 18450
rect 25342 18398 25394 18450
rect 25394 18398 25396 18450
rect 25340 18396 25396 18398
rect 25228 17612 25284 17668
rect 26124 20524 26180 20580
rect 25900 19292 25956 19348
rect 25564 18956 25620 19012
rect 25788 18956 25844 19012
rect 25676 17052 25732 17108
rect 25788 16492 25844 16548
rect 26460 22204 26516 22260
rect 27356 22428 27412 22484
rect 27804 23212 27860 23268
rect 27468 21810 27524 21812
rect 27468 21758 27470 21810
rect 27470 21758 27522 21810
rect 27522 21758 27524 21810
rect 27468 21756 27524 21758
rect 26236 19404 26292 19460
rect 26012 19068 26068 19124
rect 26236 17164 26292 17220
rect 26852 21420 26908 21476
rect 27020 21420 27076 21476
rect 26908 21084 26964 21140
rect 26460 19234 26516 19236
rect 26460 19182 26462 19234
rect 26462 19182 26514 19234
rect 26514 19182 26516 19234
rect 26460 19180 26516 19182
rect 27468 21532 27524 21588
rect 27356 21362 27412 21364
rect 27356 21310 27358 21362
rect 27358 21310 27410 21362
rect 27410 21310 27412 21362
rect 27356 21308 27412 21310
rect 27356 20972 27412 21028
rect 27244 20802 27300 20804
rect 27244 20750 27246 20802
rect 27246 20750 27298 20802
rect 27298 20750 27300 20802
rect 27244 20748 27300 20750
rect 28028 23938 28084 23940
rect 28028 23886 28030 23938
rect 28030 23886 28082 23938
rect 28082 23886 28084 23938
rect 28028 23884 28084 23886
rect 28028 23660 28084 23716
rect 27132 19852 27188 19908
rect 27244 20300 27300 20356
rect 26796 19234 26852 19236
rect 26796 19182 26798 19234
rect 26798 19182 26850 19234
rect 26850 19182 26852 19234
rect 26796 19180 26852 19182
rect 27020 19180 27076 19236
rect 26572 18338 26628 18340
rect 26572 18286 26574 18338
rect 26574 18286 26626 18338
rect 26626 18286 26628 18338
rect 26572 18284 26628 18286
rect 26460 17948 26516 18004
rect 26124 16268 26180 16324
rect 26124 15538 26180 15540
rect 26124 15486 26126 15538
rect 26126 15486 26178 15538
rect 26178 15486 26180 15538
rect 26124 15484 26180 15486
rect 26684 16716 26740 16772
rect 26460 15932 26516 15988
rect 27020 18172 27076 18228
rect 26908 17500 26964 17556
rect 27244 19234 27300 19236
rect 27244 19182 27246 19234
rect 27246 19182 27298 19234
rect 27298 19182 27300 19234
rect 27244 19180 27300 19182
rect 27356 18172 27412 18228
rect 27580 20690 27636 20692
rect 27580 20638 27582 20690
rect 27582 20638 27634 20690
rect 27634 20638 27636 20690
rect 27580 20636 27636 20638
rect 28140 23436 28196 23492
rect 28588 28642 28644 28644
rect 28588 28590 28590 28642
rect 28590 28590 28642 28642
rect 28642 28590 28644 28642
rect 28588 28588 28644 28590
rect 28476 28530 28532 28532
rect 28476 28478 28478 28530
rect 28478 28478 28530 28530
rect 28530 28478 28532 28530
rect 28476 28476 28532 28478
rect 28700 28364 28756 28420
rect 28476 26908 28532 26964
rect 28364 23772 28420 23828
rect 28588 26236 28644 26292
rect 28588 25788 28644 25844
rect 28588 25564 28644 25620
rect 28588 24780 28644 24836
rect 28476 23660 28532 23716
rect 28588 24444 28644 24500
rect 28588 23884 28644 23940
rect 27692 20188 27748 20244
rect 28476 22428 28532 22484
rect 27580 18508 27636 18564
rect 27692 18396 27748 18452
rect 27916 20636 27972 20692
rect 28028 20860 28084 20916
rect 27916 20300 27972 20356
rect 28028 19404 28084 19460
rect 27804 17948 27860 18004
rect 27356 17554 27412 17556
rect 27356 17502 27358 17554
rect 27358 17502 27410 17554
rect 27410 17502 27412 17554
rect 27356 17500 27412 17502
rect 27804 17442 27860 17444
rect 27804 17390 27806 17442
rect 27806 17390 27858 17442
rect 27858 17390 27860 17442
rect 27804 17388 27860 17390
rect 27692 16994 27748 16996
rect 27692 16942 27694 16994
rect 27694 16942 27746 16994
rect 27746 16942 27748 16994
rect 27692 16940 27748 16942
rect 27244 16716 27300 16772
rect 26348 14812 26404 14868
rect 25116 10780 25172 10836
rect 25228 11676 25284 11732
rect 23548 10556 23604 10612
rect 23548 9660 23604 9716
rect 24668 10108 24724 10164
rect 23772 9548 23828 9604
rect 24108 9324 24164 9380
rect 23660 8930 23716 8932
rect 23660 8878 23662 8930
rect 23662 8878 23714 8930
rect 23714 8878 23716 8930
rect 23660 8876 23716 8878
rect 23548 8764 23604 8820
rect 23324 8652 23380 8708
rect 23212 8428 23268 8484
rect 23100 8258 23156 8260
rect 23100 8206 23102 8258
rect 23102 8206 23154 8258
rect 23154 8206 23156 8258
rect 23100 8204 23156 8206
rect 22988 8092 23044 8148
rect 22764 7868 22820 7924
rect 22876 7756 22932 7812
rect 22652 7474 22708 7476
rect 22652 7422 22654 7474
rect 22654 7422 22706 7474
rect 22706 7422 22708 7474
rect 22652 7420 22708 7422
rect 23100 7644 23156 7700
rect 22988 5964 23044 6020
rect 23772 8540 23828 8596
rect 23324 7586 23380 7588
rect 23324 7534 23326 7586
rect 23326 7534 23378 7586
rect 23378 7534 23380 7586
rect 23324 7532 23380 7534
rect 23436 6636 23492 6692
rect 24444 9212 24500 9268
rect 24444 8764 24500 8820
rect 24332 7756 24388 7812
rect 23660 6524 23716 6580
rect 23436 5852 23492 5908
rect 23548 5740 23604 5796
rect 23212 5628 23268 5684
rect 28588 21756 28644 21812
rect 29708 32674 29764 32676
rect 29708 32622 29710 32674
rect 29710 32622 29762 32674
rect 29762 32622 29764 32674
rect 29708 32620 29764 32622
rect 29260 32338 29316 32340
rect 29260 32286 29262 32338
rect 29262 32286 29314 32338
rect 29314 32286 29316 32338
rect 29260 32284 29316 32286
rect 30156 33404 30212 33460
rect 30716 32956 30772 33012
rect 29372 31666 29428 31668
rect 29372 31614 29374 31666
rect 29374 31614 29426 31666
rect 29426 31614 29428 31666
rect 29372 31612 29428 31614
rect 30044 31612 30100 31668
rect 29148 30882 29204 30884
rect 29148 30830 29150 30882
rect 29150 30830 29202 30882
rect 29202 30830 29204 30882
rect 29148 30828 29204 30830
rect 29820 31554 29876 31556
rect 29820 31502 29822 31554
rect 29822 31502 29874 31554
rect 29874 31502 29876 31554
rect 29820 31500 29876 31502
rect 30492 31106 30548 31108
rect 30492 31054 30494 31106
rect 30494 31054 30546 31106
rect 30546 31054 30548 31106
rect 30492 31052 30548 31054
rect 29932 30770 29988 30772
rect 29932 30718 29934 30770
rect 29934 30718 29986 30770
rect 29986 30718 29988 30770
rect 29932 30716 29988 30718
rect 29148 29036 29204 29092
rect 29708 29986 29764 29988
rect 29708 29934 29710 29986
rect 29710 29934 29762 29986
rect 29762 29934 29764 29986
rect 29708 29932 29764 29934
rect 29372 28364 29428 28420
rect 29484 28476 29540 28532
rect 29372 26962 29428 26964
rect 29372 26910 29374 26962
rect 29374 26910 29426 26962
rect 29426 26910 29428 26962
rect 29372 26908 29428 26910
rect 28812 26290 28868 26292
rect 28812 26238 28814 26290
rect 28814 26238 28866 26290
rect 28866 26238 28868 26290
rect 28812 26236 28868 26238
rect 28812 25676 28868 25732
rect 28812 24780 28868 24836
rect 29596 26962 29652 26964
rect 29596 26910 29598 26962
rect 29598 26910 29650 26962
rect 29650 26910 29652 26962
rect 29596 26908 29652 26910
rect 29148 26012 29204 26068
rect 29372 25788 29428 25844
rect 30268 30156 30324 30212
rect 30492 29932 30548 29988
rect 30268 29484 30324 29540
rect 29932 28700 29988 28756
rect 30716 31612 30772 31668
rect 31052 37490 31108 37492
rect 31052 37438 31054 37490
rect 31054 37438 31106 37490
rect 31106 37438 31108 37490
rect 31052 37436 31108 37438
rect 31052 36988 31108 37044
rect 31724 38556 31780 38612
rect 31724 37436 31780 37492
rect 31276 36876 31332 36932
rect 31276 36594 31332 36596
rect 31276 36542 31278 36594
rect 31278 36542 31330 36594
rect 31330 36542 31332 36594
rect 31276 36540 31332 36542
rect 31164 35644 31220 35700
rect 31612 35698 31668 35700
rect 31612 35646 31614 35698
rect 31614 35646 31666 35698
rect 31666 35646 31668 35698
rect 31612 35644 31668 35646
rect 31724 34972 31780 35028
rect 33292 41746 33348 41748
rect 33292 41694 33294 41746
rect 33294 41694 33346 41746
rect 33346 41694 33348 41746
rect 33292 41692 33348 41694
rect 33292 40572 33348 40628
rect 33740 42530 33796 42532
rect 33740 42478 33742 42530
rect 33742 42478 33794 42530
rect 33794 42478 33796 42530
rect 33740 42476 33796 42478
rect 33516 41858 33572 41860
rect 33516 41806 33518 41858
rect 33518 41806 33570 41858
rect 33570 41806 33572 41858
rect 33516 41804 33572 41806
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35868 44492 35924 44548
rect 34860 43596 34916 43652
rect 35420 43596 35476 43652
rect 35196 43538 35252 43540
rect 35196 43486 35198 43538
rect 35198 43486 35250 43538
rect 35250 43486 35252 43538
rect 35196 43484 35252 43486
rect 34748 42812 34804 42868
rect 35084 43372 35140 43428
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34188 41692 34244 41748
rect 34412 42140 34468 42196
rect 34300 41356 34356 41412
rect 34076 41244 34132 41300
rect 33628 41186 33684 41188
rect 33628 41134 33630 41186
rect 33630 41134 33682 41186
rect 33682 41134 33684 41186
rect 33628 41132 33684 41134
rect 34748 41858 34804 41860
rect 34748 41806 34750 41858
rect 34750 41806 34802 41858
rect 34802 41806 34804 41858
rect 34748 41804 34804 41806
rect 34860 41692 34916 41748
rect 34860 41132 34916 41188
rect 33852 40796 33908 40852
rect 32956 38780 33012 38836
rect 32284 37884 32340 37940
rect 32732 37884 32788 37940
rect 32508 37772 32564 37828
rect 32060 37660 32116 37716
rect 32396 37490 32452 37492
rect 32396 37438 32398 37490
rect 32398 37438 32450 37490
rect 32450 37438 32452 37490
rect 32396 37436 32452 37438
rect 32284 37100 32340 37156
rect 31948 36988 32004 37044
rect 32508 36316 32564 36372
rect 32620 36258 32676 36260
rect 32620 36206 32622 36258
rect 32622 36206 32674 36258
rect 32674 36206 32676 36258
rect 32620 36204 32676 36206
rect 32620 35420 32676 35476
rect 32284 35308 32340 35364
rect 32172 35084 32228 35140
rect 30940 34130 30996 34132
rect 30940 34078 30942 34130
rect 30942 34078 30994 34130
rect 30994 34078 30996 34130
rect 30940 34076 30996 34078
rect 31164 33122 31220 33124
rect 31164 33070 31166 33122
rect 31166 33070 31218 33122
rect 31218 33070 31220 33122
rect 31164 33068 31220 33070
rect 31500 32562 31556 32564
rect 31500 32510 31502 32562
rect 31502 32510 31554 32562
rect 31554 32510 31556 32562
rect 31500 32508 31556 32510
rect 31388 31778 31444 31780
rect 31388 31726 31390 31778
rect 31390 31726 31442 31778
rect 31442 31726 31444 31778
rect 31388 31724 31444 31726
rect 30940 31500 30996 31556
rect 30940 31276 30996 31332
rect 31164 31276 31220 31332
rect 31836 34076 31892 34132
rect 31612 31836 31668 31892
rect 31500 31612 31556 31668
rect 30716 30268 30772 30324
rect 30716 30044 30772 30100
rect 30716 29148 30772 29204
rect 30828 29932 30884 29988
rect 30828 28812 30884 28868
rect 30716 27746 30772 27748
rect 30716 27694 30718 27746
rect 30718 27694 30770 27746
rect 30770 27694 30772 27746
rect 30716 27692 30772 27694
rect 30156 27132 30212 27188
rect 30380 26962 30436 26964
rect 30380 26910 30382 26962
rect 30382 26910 30434 26962
rect 30434 26910 30436 26962
rect 30380 26908 30436 26910
rect 29820 25676 29876 25732
rect 30156 26460 30212 26516
rect 30604 26796 30660 26852
rect 29260 25506 29316 25508
rect 29260 25454 29262 25506
rect 29262 25454 29314 25506
rect 29314 25454 29316 25506
rect 29260 25452 29316 25454
rect 29260 25116 29316 25172
rect 30492 26402 30548 26404
rect 30492 26350 30494 26402
rect 30494 26350 30546 26402
rect 30546 26350 30548 26402
rect 30492 26348 30548 26350
rect 30716 26460 30772 26516
rect 31052 30210 31108 30212
rect 31052 30158 31054 30210
rect 31054 30158 31106 30210
rect 31106 30158 31108 30210
rect 31052 30156 31108 30158
rect 31388 29426 31444 29428
rect 31388 29374 31390 29426
rect 31390 29374 31442 29426
rect 31442 29374 31444 29426
rect 31388 29372 31444 29374
rect 31052 29202 31108 29204
rect 31052 29150 31054 29202
rect 31054 29150 31106 29202
rect 31106 29150 31108 29202
rect 31052 29148 31108 29150
rect 31276 28642 31332 28644
rect 31276 28590 31278 28642
rect 31278 28590 31330 28642
rect 31330 28590 31332 28642
rect 31276 28588 31332 28590
rect 31164 27858 31220 27860
rect 31164 27806 31166 27858
rect 31166 27806 31218 27858
rect 31218 27806 31220 27858
rect 31164 27804 31220 27806
rect 32060 33516 32116 33572
rect 31836 33068 31892 33124
rect 32844 35084 32900 35140
rect 32620 35026 32676 35028
rect 32620 34974 32622 35026
rect 32622 34974 32674 35026
rect 32674 34974 32676 35026
rect 32620 34972 32676 34974
rect 34860 40796 34916 40852
rect 34524 40626 34580 40628
rect 34524 40574 34526 40626
rect 34526 40574 34578 40626
rect 34578 40574 34580 40626
rect 34524 40572 34580 40574
rect 35308 42700 35364 42756
rect 35756 43484 35812 43540
rect 35644 43426 35700 43428
rect 35644 43374 35646 43426
rect 35646 43374 35698 43426
rect 35698 43374 35700 43426
rect 35644 43372 35700 43374
rect 35980 43932 36036 43988
rect 35980 43650 36036 43652
rect 35980 43598 35982 43650
rect 35982 43598 36034 43650
rect 36034 43598 36036 43650
rect 35980 43596 36036 43598
rect 37100 45164 37156 45220
rect 40012 47458 40068 47460
rect 40012 47406 40014 47458
rect 40014 47406 40066 47458
rect 40066 47406 40068 47458
rect 40012 47404 40068 47406
rect 41244 47404 41300 47460
rect 38780 47346 38836 47348
rect 38780 47294 38782 47346
rect 38782 47294 38834 47346
rect 38834 47294 38836 47346
rect 38780 47292 38836 47294
rect 37772 46844 37828 46900
rect 37212 45052 37268 45108
rect 37324 44828 37380 44884
rect 36988 44380 37044 44436
rect 37212 44434 37268 44436
rect 37212 44382 37214 44434
rect 37214 44382 37266 44434
rect 37266 44382 37268 44434
rect 37212 44380 37268 44382
rect 35868 42924 35924 42980
rect 35084 41804 35140 41860
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35532 41186 35588 41188
rect 35532 41134 35534 41186
rect 35534 41134 35586 41186
rect 35586 41134 35588 41186
rect 35532 41132 35588 41134
rect 35196 41020 35252 41076
rect 35868 42140 35924 42196
rect 36988 43932 37044 43988
rect 36540 43538 36596 43540
rect 36540 43486 36542 43538
rect 36542 43486 36594 43538
rect 36594 43486 36596 43538
rect 36540 43484 36596 43486
rect 36652 43260 36708 43316
rect 36428 42530 36484 42532
rect 36428 42478 36430 42530
rect 36430 42478 36482 42530
rect 36482 42478 36484 42530
rect 36428 42476 36484 42478
rect 37100 43820 37156 43876
rect 37212 43372 37268 43428
rect 37100 43260 37156 43316
rect 36876 42140 36932 42196
rect 36204 42028 36260 42084
rect 37772 43260 37828 43316
rect 37548 43148 37604 43204
rect 37548 42978 37604 42980
rect 37548 42926 37550 42978
rect 37550 42926 37602 42978
rect 37602 42926 37604 42978
rect 37548 42924 37604 42926
rect 37436 42028 37492 42084
rect 37100 41692 37156 41748
rect 36204 41410 36260 41412
rect 36204 41358 36206 41410
rect 36206 41358 36258 41410
rect 36258 41358 36260 41410
rect 36204 41356 36260 41358
rect 35756 41020 35812 41076
rect 35196 40796 35252 40852
rect 34412 40402 34468 40404
rect 34412 40350 34414 40402
rect 34414 40350 34466 40402
rect 34466 40350 34468 40402
rect 34412 40348 34468 40350
rect 33964 40290 34020 40292
rect 33964 40238 33966 40290
rect 33966 40238 34018 40290
rect 34018 40238 34020 40290
rect 33964 40236 34020 40238
rect 33852 38780 33908 38836
rect 33180 38610 33236 38612
rect 33180 38558 33182 38610
rect 33182 38558 33234 38610
rect 33234 38558 33236 38610
rect 33180 38556 33236 38558
rect 33068 36988 33124 37044
rect 33628 36876 33684 36932
rect 33292 36482 33348 36484
rect 33292 36430 33294 36482
rect 33294 36430 33346 36482
rect 33346 36430 33348 36482
rect 33292 36428 33348 36430
rect 33404 35644 33460 35700
rect 33068 34130 33124 34132
rect 33068 34078 33070 34130
rect 33070 34078 33122 34130
rect 33122 34078 33124 34130
rect 33068 34076 33124 34078
rect 32284 32956 32340 33012
rect 32396 33292 32452 33348
rect 32284 32732 32340 32788
rect 31948 31836 32004 31892
rect 31836 31666 31892 31668
rect 31836 31614 31838 31666
rect 31838 31614 31890 31666
rect 31890 31614 31892 31666
rect 31836 31612 31892 31614
rect 31948 31106 32004 31108
rect 31948 31054 31950 31106
rect 31950 31054 32002 31106
rect 32002 31054 32004 31106
rect 31948 31052 32004 31054
rect 31724 30994 31780 30996
rect 31724 30942 31726 30994
rect 31726 30942 31778 30994
rect 31778 30942 31780 30994
rect 31724 30940 31780 30942
rect 31836 30268 31892 30324
rect 31724 30044 31780 30100
rect 31724 28812 31780 28868
rect 31500 27356 31556 27412
rect 31724 26908 31780 26964
rect 30940 26572 30996 26628
rect 31612 26796 31668 26852
rect 30156 25340 30212 25396
rect 30156 25116 30212 25172
rect 29596 25004 29652 25060
rect 29484 24668 29540 24724
rect 29484 23772 29540 23828
rect 29260 23548 29316 23604
rect 28924 23436 28980 23492
rect 28924 23266 28980 23268
rect 28924 23214 28926 23266
rect 28926 23214 28978 23266
rect 28978 23214 28980 23266
rect 28924 23212 28980 23214
rect 30044 24610 30100 24612
rect 30044 24558 30046 24610
rect 30046 24558 30098 24610
rect 30098 24558 30100 24610
rect 30044 24556 30100 24558
rect 29820 24444 29876 24500
rect 30828 24892 30884 24948
rect 30716 24498 30772 24500
rect 30716 24446 30718 24498
rect 30718 24446 30770 24498
rect 30770 24446 30772 24498
rect 30716 24444 30772 24446
rect 30380 23772 30436 23828
rect 28252 21308 28308 21364
rect 28700 20972 28756 21028
rect 28364 20524 28420 20580
rect 28252 20188 28308 20244
rect 28252 19346 28308 19348
rect 28252 19294 28254 19346
rect 28254 19294 28306 19346
rect 28306 19294 28308 19346
rect 28252 19292 28308 19294
rect 28588 19292 28644 19348
rect 28140 18844 28196 18900
rect 28028 18172 28084 18228
rect 28140 17724 28196 17780
rect 28588 18956 28644 19012
rect 28700 18732 28756 18788
rect 29260 22482 29316 22484
rect 29260 22430 29262 22482
rect 29262 22430 29314 22482
rect 29314 22430 29316 22482
rect 29260 22428 29316 22430
rect 28924 18396 28980 18452
rect 29372 21868 29428 21924
rect 29932 23436 29988 23492
rect 30268 23378 30324 23380
rect 30268 23326 30270 23378
rect 30270 23326 30322 23378
rect 30322 23326 30324 23378
rect 30268 23324 30324 23326
rect 30492 23266 30548 23268
rect 30492 23214 30494 23266
rect 30494 23214 30546 23266
rect 30546 23214 30548 23266
rect 30492 23212 30548 23214
rect 30492 22764 30548 22820
rect 29484 21532 29540 21588
rect 29596 21308 29652 21364
rect 29708 21756 29764 21812
rect 30828 23826 30884 23828
rect 30828 23774 30830 23826
rect 30830 23774 30882 23826
rect 30882 23774 30884 23826
rect 30828 23772 30884 23774
rect 31052 26178 31108 26180
rect 31052 26126 31054 26178
rect 31054 26126 31106 26178
rect 31106 26126 31108 26178
rect 31052 26124 31108 26126
rect 31052 25676 31108 25732
rect 31612 25228 31668 25284
rect 31612 24946 31668 24948
rect 31612 24894 31614 24946
rect 31614 24894 31666 24946
rect 31666 24894 31668 24946
rect 31612 24892 31668 24894
rect 31836 24946 31892 24948
rect 31836 24894 31838 24946
rect 31838 24894 31890 24946
rect 31890 24894 31892 24946
rect 31836 24892 31892 24894
rect 31388 24722 31444 24724
rect 31388 24670 31390 24722
rect 31390 24670 31442 24722
rect 31442 24670 31444 24722
rect 31388 24668 31444 24670
rect 31164 23378 31220 23380
rect 31164 23326 31166 23378
rect 31166 23326 31218 23378
rect 31218 23326 31220 23378
rect 31164 23324 31220 23326
rect 31612 24444 31668 24500
rect 31500 23436 31556 23492
rect 31724 24332 31780 24388
rect 30940 22316 30996 22372
rect 29708 21084 29764 21140
rect 30268 21586 30324 21588
rect 30268 21534 30270 21586
rect 30270 21534 30322 21586
rect 30322 21534 30324 21586
rect 30268 21532 30324 21534
rect 29820 20972 29876 21028
rect 29932 21420 29988 21476
rect 29708 20578 29764 20580
rect 29708 20526 29710 20578
rect 29710 20526 29762 20578
rect 29762 20526 29764 20578
rect 29708 20524 29764 20526
rect 29596 19404 29652 19460
rect 29708 19346 29764 19348
rect 29708 19294 29710 19346
rect 29710 19294 29762 19346
rect 29762 19294 29764 19346
rect 29708 19292 29764 19294
rect 29148 19234 29204 19236
rect 29148 19182 29150 19234
rect 29150 19182 29202 19234
rect 29202 19182 29204 19234
rect 29148 19180 29204 19182
rect 29484 19068 29540 19124
rect 29372 18508 29428 18564
rect 29708 19010 29764 19012
rect 29708 18958 29710 19010
rect 29710 18958 29762 19010
rect 29762 18958 29764 19010
rect 29708 18956 29764 18958
rect 29036 18284 29092 18340
rect 29260 18396 29316 18452
rect 28364 17778 28420 17780
rect 28364 17726 28366 17778
rect 28366 17726 28418 17778
rect 28418 17726 28420 17778
rect 28364 17724 28420 17726
rect 28588 17724 28644 17780
rect 28252 17612 28308 17668
rect 30156 20972 30212 21028
rect 30044 20524 30100 20580
rect 30268 20860 30324 20916
rect 29932 19516 29988 19572
rect 30044 18956 30100 19012
rect 30940 21532 30996 21588
rect 30716 20914 30772 20916
rect 30716 20862 30718 20914
rect 30718 20862 30770 20914
rect 30770 20862 30772 20914
rect 30716 20860 30772 20862
rect 31500 21586 31556 21588
rect 31500 21534 31502 21586
rect 31502 21534 31554 21586
rect 31554 21534 31556 21586
rect 31500 21532 31556 21534
rect 31388 21420 31444 21476
rect 32060 30940 32116 30996
rect 32620 31612 32676 31668
rect 32172 29426 32228 29428
rect 32172 29374 32174 29426
rect 32174 29374 32226 29426
rect 32226 29374 32228 29426
rect 32172 29372 32228 29374
rect 32284 28028 32340 28084
rect 32060 27692 32116 27748
rect 32284 27692 32340 27748
rect 32508 27858 32564 27860
rect 32508 27806 32510 27858
rect 32510 27806 32562 27858
rect 32562 27806 32564 27858
rect 32508 27804 32564 27806
rect 32060 26796 32116 26852
rect 32060 25676 32116 25732
rect 32508 26796 32564 26852
rect 34636 39788 34692 39844
rect 34972 40348 35028 40404
rect 33852 38556 33908 38612
rect 33964 37996 34020 38052
rect 34076 37212 34132 37268
rect 34076 36540 34132 36596
rect 33740 35420 33796 35476
rect 33852 35756 33908 35812
rect 33516 33292 33572 33348
rect 33180 32732 33236 32788
rect 33292 33180 33348 33236
rect 33180 32450 33236 32452
rect 33180 32398 33182 32450
rect 33182 32398 33234 32450
rect 33234 32398 33236 32450
rect 33180 32396 33236 32398
rect 33628 32060 33684 32116
rect 33180 30940 33236 30996
rect 33068 29596 33124 29652
rect 33404 30156 33460 30212
rect 33292 29708 33348 29764
rect 33516 29596 33572 29652
rect 33068 29426 33124 29428
rect 33068 29374 33070 29426
rect 33070 29374 33122 29426
rect 33122 29374 33124 29426
rect 33068 29372 33124 29374
rect 33180 28028 33236 28084
rect 32732 26236 32788 26292
rect 33180 27634 33236 27636
rect 33180 27582 33182 27634
rect 33182 27582 33234 27634
rect 33234 27582 33236 27634
rect 33180 27580 33236 27582
rect 33292 26796 33348 26852
rect 33516 29372 33572 29428
rect 33740 31836 33796 31892
rect 33852 31276 33908 31332
rect 33964 34018 34020 34020
rect 33964 33966 33966 34018
rect 33966 33966 34018 34018
rect 34018 33966 34020 34018
rect 33964 33964 34020 33966
rect 33852 30380 33908 30436
rect 35196 40124 35252 40180
rect 35420 40962 35476 40964
rect 35420 40910 35422 40962
rect 35422 40910 35474 40962
rect 35474 40910 35476 40962
rect 35420 40908 35476 40910
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35308 39788 35364 39844
rect 36092 40460 36148 40516
rect 35532 39564 35588 39620
rect 35420 38946 35476 38948
rect 35420 38894 35422 38946
rect 35422 38894 35474 38946
rect 35474 38894 35476 38946
rect 35420 38892 35476 38894
rect 34300 38722 34356 38724
rect 34300 38670 34302 38722
rect 34302 38670 34354 38722
rect 34354 38670 34356 38722
rect 34300 38668 34356 38670
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34860 38108 34916 38164
rect 35196 38108 35252 38164
rect 34860 37938 34916 37940
rect 34860 37886 34862 37938
rect 34862 37886 34914 37938
rect 34914 37886 34916 37938
rect 34860 37884 34916 37886
rect 34412 37100 34468 37156
rect 34972 37548 35028 37604
rect 34972 36652 35028 36708
rect 34300 36370 34356 36372
rect 34300 36318 34302 36370
rect 34302 36318 34354 36370
rect 34354 36318 34356 36370
rect 34300 36316 34356 36318
rect 34188 35644 34244 35700
rect 35644 39394 35700 39396
rect 35644 39342 35646 39394
rect 35646 39342 35698 39394
rect 35698 39342 35700 39394
rect 35644 39340 35700 39342
rect 35980 39564 36036 39620
rect 35532 38108 35588 38164
rect 35868 39116 35924 39172
rect 35756 38444 35812 38500
rect 35756 37938 35812 37940
rect 35756 37886 35758 37938
rect 35758 37886 35810 37938
rect 35810 37886 35812 37938
rect 35756 37884 35812 37886
rect 35868 37826 35924 37828
rect 35868 37774 35870 37826
rect 35870 37774 35922 37826
rect 35922 37774 35924 37826
rect 35868 37772 35924 37774
rect 36204 40236 36260 40292
rect 36876 41020 36932 41076
rect 36428 40348 36484 40404
rect 36540 40236 36596 40292
rect 36316 39506 36372 39508
rect 36316 39454 36318 39506
rect 36318 39454 36370 39506
rect 36370 39454 36372 39506
rect 36316 39452 36372 39454
rect 35980 37660 36036 37716
rect 36092 38444 36148 38500
rect 36204 38050 36260 38052
rect 36204 37998 36206 38050
rect 36206 37998 36258 38050
rect 36258 37998 36260 38050
rect 36204 37996 36260 37998
rect 36428 38444 36484 38500
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34300 33234 34356 33236
rect 34300 33182 34302 33234
rect 34302 33182 34354 33234
rect 34354 33182 34356 33234
rect 34300 33180 34356 33182
rect 34300 32786 34356 32788
rect 34300 32734 34302 32786
rect 34302 32734 34354 32786
rect 34354 32734 34356 32786
rect 34300 32732 34356 32734
rect 34076 32060 34132 32116
rect 34412 32450 34468 32452
rect 34412 32398 34414 32450
rect 34414 32398 34466 32450
rect 34466 32398 34468 32450
rect 34412 32396 34468 32398
rect 34188 31388 34244 31444
rect 34076 31276 34132 31332
rect 34524 31276 34580 31332
rect 34412 31106 34468 31108
rect 34412 31054 34414 31106
rect 34414 31054 34466 31106
rect 34466 31054 34468 31106
rect 34412 31052 34468 31054
rect 33964 29932 34020 29988
rect 34188 30940 34244 30996
rect 33740 29426 33796 29428
rect 33740 29374 33742 29426
rect 33742 29374 33794 29426
rect 33794 29374 33796 29426
rect 33740 29372 33796 29374
rect 33852 29314 33908 29316
rect 33852 29262 33854 29314
rect 33854 29262 33906 29314
rect 33906 29262 33908 29314
rect 33852 29260 33908 29262
rect 33628 27970 33684 27972
rect 33628 27918 33630 27970
rect 33630 27918 33682 27970
rect 33682 27918 33684 27970
rect 33628 27916 33684 27918
rect 34076 28588 34132 28644
rect 33852 27580 33908 27636
rect 33404 26236 33460 26292
rect 34076 27468 34132 27524
rect 33068 26178 33124 26180
rect 33068 26126 33070 26178
rect 33070 26126 33122 26178
rect 33122 26126 33124 26178
rect 33068 26124 33124 26126
rect 33068 25788 33124 25844
rect 32844 25676 32900 25732
rect 32396 25116 32452 25172
rect 32060 24722 32116 24724
rect 32060 24670 32062 24722
rect 32062 24670 32114 24722
rect 32114 24670 32116 24722
rect 32060 24668 32116 24670
rect 31948 23266 32004 23268
rect 31948 23214 31950 23266
rect 31950 23214 32002 23266
rect 32002 23214 32004 23266
rect 31948 23212 32004 23214
rect 31836 22092 31892 22148
rect 32172 22258 32228 22260
rect 32172 22206 32174 22258
rect 32174 22206 32226 22258
rect 32226 22206 32228 22258
rect 32172 22204 32228 22206
rect 32172 21756 32228 21812
rect 31836 21532 31892 21588
rect 33180 25116 33236 25172
rect 32956 24892 33012 24948
rect 33516 25618 33572 25620
rect 33516 25566 33518 25618
rect 33518 25566 33570 25618
rect 33570 25566 33572 25618
rect 33516 25564 33572 25566
rect 33516 23436 33572 23492
rect 33852 26124 33908 26180
rect 33740 25506 33796 25508
rect 33740 25454 33742 25506
rect 33742 25454 33794 25506
rect 33794 25454 33796 25506
rect 33740 25452 33796 25454
rect 33964 25340 34020 25396
rect 33964 24108 34020 24164
rect 33628 23324 33684 23380
rect 33964 23436 34020 23492
rect 33852 23042 33908 23044
rect 33852 22990 33854 23042
rect 33854 22990 33906 23042
rect 33906 22990 33908 23042
rect 33852 22988 33908 22990
rect 33516 22876 33572 22932
rect 32620 22258 32676 22260
rect 32620 22206 32622 22258
rect 32622 22206 32674 22258
rect 32674 22206 32676 22258
rect 32620 22204 32676 22206
rect 33068 22258 33124 22260
rect 33068 22206 33070 22258
rect 33070 22206 33122 22258
rect 33122 22206 33124 22258
rect 33068 22204 33124 22206
rect 33068 21810 33124 21812
rect 33068 21758 33070 21810
rect 33070 21758 33122 21810
rect 33122 21758 33124 21810
rect 33068 21756 33124 21758
rect 32508 21532 32564 21588
rect 31612 21420 31668 21476
rect 32396 21474 32452 21476
rect 32396 21422 32398 21474
rect 32398 21422 32450 21474
rect 32450 21422 32452 21474
rect 32396 21420 32452 21422
rect 31276 20860 31332 20916
rect 31052 19964 31108 20020
rect 31612 20524 31668 20580
rect 30604 19628 30660 19684
rect 30604 19404 30660 19460
rect 30492 19346 30548 19348
rect 30492 19294 30494 19346
rect 30494 19294 30546 19346
rect 30546 19294 30548 19346
rect 30492 19292 30548 19294
rect 30268 19068 30324 19124
rect 29708 18172 29764 18228
rect 29820 18396 29876 18452
rect 29036 17612 29092 17668
rect 28140 17388 28196 17444
rect 28140 16716 28196 16772
rect 28028 16604 28084 16660
rect 27692 16156 27748 16212
rect 27244 15986 27300 15988
rect 27244 15934 27246 15986
rect 27246 15934 27298 15986
rect 27298 15934 27300 15986
rect 27244 15932 27300 15934
rect 27580 16044 27636 16100
rect 28028 15932 28084 15988
rect 27804 15260 27860 15316
rect 26572 13916 26628 13972
rect 25452 12572 25508 12628
rect 25340 11564 25396 11620
rect 26572 13580 26628 13636
rect 26460 13132 26516 13188
rect 26124 12178 26180 12180
rect 26124 12126 26126 12178
rect 26126 12126 26178 12178
rect 26178 12126 26180 12178
rect 26124 12124 26180 12126
rect 25564 12066 25620 12068
rect 25564 12014 25566 12066
rect 25566 12014 25618 12066
rect 25618 12014 25620 12066
rect 25564 12012 25620 12014
rect 27020 13746 27076 13748
rect 27020 13694 27022 13746
rect 27022 13694 27074 13746
rect 27074 13694 27076 13746
rect 27020 13692 27076 13694
rect 26796 12236 26852 12292
rect 26908 12124 26964 12180
rect 25788 11564 25844 11620
rect 25340 9100 25396 9156
rect 24780 8988 24836 9044
rect 24668 8540 24724 8596
rect 25228 8204 25284 8260
rect 24892 8092 24948 8148
rect 24556 7420 24612 7476
rect 24780 7868 24836 7924
rect 24780 7308 24836 7364
rect 24220 6636 24276 6692
rect 24220 6018 24276 6020
rect 24220 5966 24222 6018
rect 24222 5966 24274 6018
rect 24274 5966 24276 6018
rect 24220 5964 24276 5966
rect 23772 5180 23828 5236
rect 25228 7980 25284 8036
rect 25340 7756 25396 7812
rect 25788 10892 25844 10948
rect 26460 11116 26516 11172
rect 25788 10220 25844 10276
rect 26684 10444 26740 10500
rect 25564 9266 25620 9268
rect 25564 9214 25566 9266
rect 25566 9214 25618 9266
rect 25618 9214 25620 9266
rect 25564 9212 25620 9214
rect 28252 16098 28308 16100
rect 28252 16046 28254 16098
rect 28254 16046 28306 16098
rect 28306 16046 28308 16098
rect 28252 16044 28308 16046
rect 27356 13580 27412 13636
rect 27468 13356 27524 13412
rect 27692 13692 27748 13748
rect 28476 16156 28532 16212
rect 28588 16044 28644 16100
rect 28252 13692 28308 13748
rect 27804 13132 27860 13188
rect 28028 13244 28084 13300
rect 28364 13020 28420 13076
rect 29148 17500 29204 17556
rect 29260 17388 29316 17444
rect 29596 17836 29652 17892
rect 30380 19010 30436 19012
rect 30380 18958 30382 19010
rect 30382 18958 30434 19010
rect 30434 18958 30436 19010
rect 30380 18956 30436 18958
rect 30828 18956 30884 19012
rect 30828 18508 30884 18564
rect 30604 18338 30660 18340
rect 30604 18286 30606 18338
rect 30606 18286 30658 18338
rect 30658 18286 30660 18338
rect 30604 18284 30660 18286
rect 31276 19346 31332 19348
rect 31276 19294 31278 19346
rect 31278 19294 31330 19346
rect 31330 19294 31332 19346
rect 31276 19292 31332 19294
rect 31388 19122 31444 19124
rect 31388 19070 31390 19122
rect 31390 19070 31442 19122
rect 31442 19070 31444 19122
rect 31388 19068 31444 19070
rect 31164 18956 31220 19012
rect 31276 18844 31332 18900
rect 31612 19740 31668 19796
rect 32060 19292 32116 19348
rect 31612 18620 31668 18676
rect 31052 18396 31108 18452
rect 31052 18172 31108 18228
rect 29596 16492 29652 16548
rect 29932 15484 29988 15540
rect 29260 15260 29316 15316
rect 29372 14530 29428 14532
rect 29372 14478 29374 14530
rect 29374 14478 29426 14530
rect 29426 14478 29428 14530
rect 29372 14476 29428 14478
rect 28812 13746 28868 13748
rect 28812 13694 28814 13746
rect 28814 13694 28866 13746
rect 28866 13694 28868 13746
rect 28812 13692 28868 13694
rect 29484 13356 29540 13412
rect 28028 12796 28084 12852
rect 27916 12236 27972 12292
rect 27244 10444 27300 10500
rect 27468 11170 27524 11172
rect 27468 11118 27470 11170
rect 27470 11118 27522 11170
rect 27522 11118 27524 11170
rect 27468 11116 27524 11118
rect 28028 11170 28084 11172
rect 28028 11118 28030 11170
rect 28030 11118 28082 11170
rect 28082 11118 28084 11170
rect 28028 11116 28084 11118
rect 28364 10556 28420 10612
rect 28140 10498 28196 10500
rect 28140 10446 28142 10498
rect 28142 10446 28194 10498
rect 28194 10446 28196 10498
rect 28140 10444 28196 10446
rect 27356 10220 27412 10276
rect 27804 10108 27860 10164
rect 27468 9884 27524 9940
rect 28140 9660 28196 9716
rect 27132 9266 27188 9268
rect 27132 9214 27134 9266
rect 27134 9214 27186 9266
rect 27186 9214 27188 9266
rect 27132 9212 27188 9214
rect 25900 9154 25956 9156
rect 25900 9102 25902 9154
rect 25902 9102 25954 9154
rect 25954 9102 25956 9154
rect 25900 9100 25956 9102
rect 25564 8316 25620 8372
rect 25676 7362 25732 7364
rect 25676 7310 25678 7362
rect 25678 7310 25730 7362
rect 25730 7310 25732 7362
rect 25676 7308 25732 7310
rect 25788 7980 25844 8036
rect 25452 6636 25508 6692
rect 25228 5180 25284 5236
rect 24668 4450 24724 4452
rect 24668 4398 24670 4450
rect 24670 4398 24722 4450
rect 24722 4398 24724 4450
rect 24668 4396 24724 4398
rect 28588 11394 28644 11396
rect 28588 11342 28590 11394
rect 28590 11342 28642 11394
rect 28642 11342 28644 11394
rect 28588 11340 28644 11342
rect 28812 11116 28868 11172
rect 29260 11676 29316 11732
rect 29372 11452 29428 11508
rect 29484 11676 29540 11732
rect 28924 10780 28980 10836
rect 29148 10668 29204 10724
rect 29372 10610 29428 10612
rect 29372 10558 29374 10610
rect 29374 10558 29426 10610
rect 29426 10558 29428 10610
rect 29372 10556 29428 10558
rect 31276 17836 31332 17892
rect 32172 19010 32228 19012
rect 32172 18958 32174 19010
rect 32174 18958 32226 19010
rect 32226 18958 32228 19010
rect 32172 18956 32228 18958
rect 32060 18732 32116 18788
rect 31948 18620 32004 18676
rect 32620 20300 32676 20356
rect 33180 19906 33236 19908
rect 33180 19854 33182 19906
rect 33182 19854 33234 19906
rect 33234 19854 33236 19906
rect 33180 19852 33236 19854
rect 32620 19234 32676 19236
rect 32620 19182 32622 19234
rect 32622 19182 32674 19234
rect 32674 19182 32676 19234
rect 32620 19180 32676 19182
rect 33628 22764 33684 22820
rect 35532 35084 35588 35140
rect 35644 36652 35700 36708
rect 35980 36428 36036 36484
rect 37100 40908 37156 40964
rect 37660 42140 37716 42196
rect 40348 47180 40404 47236
rect 38332 44604 38388 44660
rect 38332 44434 38388 44436
rect 38332 44382 38334 44434
rect 38334 44382 38386 44434
rect 38386 44382 38388 44434
rect 38332 44380 38388 44382
rect 38332 43484 38388 43540
rect 37884 41692 37940 41748
rect 38108 43148 38164 43204
rect 38108 41970 38164 41972
rect 38108 41918 38110 41970
rect 38110 41918 38162 41970
rect 38162 41918 38164 41970
rect 38108 41916 38164 41918
rect 37548 40684 37604 40740
rect 36988 40124 37044 40180
rect 36764 38668 36820 38724
rect 37324 40402 37380 40404
rect 37324 40350 37326 40402
rect 37326 40350 37378 40402
rect 37378 40350 37380 40402
rect 37324 40348 37380 40350
rect 37212 39618 37268 39620
rect 37212 39566 37214 39618
rect 37214 39566 37266 39618
rect 37266 39566 37268 39618
rect 37212 39564 37268 39566
rect 37884 40348 37940 40404
rect 37548 39564 37604 39620
rect 37324 39506 37380 39508
rect 37324 39454 37326 39506
rect 37326 39454 37378 39506
rect 37378 39454 37380 39506
rect 37324 39452 37380 39454
rect 37660 39116 37716 39172
rect 37548 39004 37604 39060
rect 36652 36428 36708 36484
rect 36876 38220 36932 38276
rect 36988 38162 37044 38164
rect 36988 38110 36990 38162
rect 36990 38110 37042 38162
rect 37042 38110 37044 38162
rect 36988 38108 37044 38110
rect 36876 37324 36932 37380
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35084 33516 35140 33572
rect 34748 33404 34804 33460
rect 36428 33458 36484 33460
rect 36428 33406 36430 33458
rect 36430 33406 36482 33458
rect 36482 33406 36484 33458
rect 36428 33404 36484 33406
rect 36204 32450 36260 32452
rect 36204 32398 36206 32450
rect 36206 32398 36258 32450
rect 36258 32398 36260 32450
rect 36204 32396 36260 32398
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35868 31890 35924 31892
rect 35868 31838 35870 31890
rect 35870 31838 35922 31890
rect 35922 31838 35924 31890
rect 35868 31836 35924 31838
rect 35980 31778 36036 31780
rect 35980 31726 35982 31778
rect 35982 31726 36034 31778
rect 36034 31726 36036 31778
rect 35980 31724 36036 31726
rect 34524 30940 34580 30996
rect 34748 31388 34804 31444
rect 34412 30716 34468 30772
rect 35084 31276 35140 31332
rect 34860 29708 34916 29764
rect 36092 31388 36148 31444
rect 35756 31276 35812 31332
rect 35308 30994 35364 30996
rect 35308 30942 35310 30994
rect 35310 30942 35362 30994
rect 35362 30942 35364 30994
rect 35308 30940 35364 30942
rect 35196 30716 35252 30772
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 30210 35252 30212
rect 35196 30158 35198 30210
rect 35198 30158 35250 30210
rect 35250 30158 35252 30210
rect 35196 30156 35252 30158
rect 36316 31500 36372 31556
rect 36652 31052 36708 31108
rect 36540 30492 36596 30548
rect 36428 30098 36484 30100
rect 36428 30046 36430 30098
rect 36430 30046 36482 30098
rect 36482 30046 36484 30098
rect 36428 30044 36484 30046
rect 36428 29650 36484 29652
rect 36428 29598 36430 29650
rect 36430 29598 36482 29650
rect 36482 29598 36484 29650
rect 36428 29596 36484 29598
rect 34860 29538 34916 29540
rect 34860 29486 34862 29538
rect 34862 29486 34914 29538
rect 34914 29486 34916 29538
rect 34860 29484 34916 29486
rect 35196 29426 35252 29428
rect 35196 29374 35198 29426
rect 35198 29374 35250 29426
rect 35250 29374 35252 29426
rect 35196 29372 35252 29374
rect 35756 29260 35812 29316
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34636 28812 34692 28868
rect 34412 27858 34468 27860
rect 34412 27806 34414 27858
rect 34414 27806 34466 27858
rect 34466 27806 34468 27858
rect 34412 27804 34468 27806
rect 35308 28754 35364 28756
rect 35308 28702 35310 28754
rect 35310 28702 35362 28754
rect 35362 28702 35364 28754
rect 35308 28700 35364 28702
rect 35980 29202 36036 29204
rect 35980 29150 35982 29202
rect 35982 29150 36034 29202
rect 36034 29150 36036 29202
rect 35980 29148 36036 29150
rect 35980 28700 36036 28756
rect 35868 28642 35924 28644
rect 35868 28590 35870 28642
rect 35870 28590 35922 28642
rect 35922 28590 35924 28642
rect 35868 28588 35924 28590
rect 35644 27916 35700 27972
rect 35196 27466 35252 27468
rect 34860 27356 34916 27412
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34524 25506 34580 25508
rect 34524 25454 34526 25506
rect 34526 25454 34578 25506
rect 34578 25454 34580 25506
rect 34524 25452 34580 25454
rect 34636 26236 34692 26292
rect 34300 25340 34356 25396
rect 35756 28476 35812 28532
rect 36204 27916 36260 27972
rect 35756 27132 35812 27188
rect 36204 27692 36260 27748
rect 35644 27020 35700 27076
rect 36988 35698 37044 35700
rect 36988 35646 36990 35698
rect 36990 35646 37042 35698
rect 37042 35646 37044 35698
rect 36988 35644 37044 35646
rect 37884 38444 37940 38500
rect 38668 43148 38724 43204
rect 38780 42924 38836 42980
rect 38556 42530 38612 42532
rect 38556 42478 38558 42530
rect 38558 42478 38610 42530
rect 38610 42478 38612 42530
rect 38556 42476 38612 42478
rect 38444 42364 38500 42420
rect 38220 41804 38276 41860
rect 38444 41916 38500 41972
rect 38668 42140 38724 42196
rect 38556 41580 38612 41636
rect 38108 40402 38164 40404
rect 38108 40350 38110 40402
rect 38110 40350 38162 40402
rect 38162 40350 38164 40402
rect 38108 40348 38164 40350
rect 38220 40796 38276 40852
rect 37660 38332 37716 38388
rect 37324 36370 37380 36372
rect 37324 36318 37326 36370
rect 37326 36318 37378 36370
rect 37378 36318 37380 36370
rect 37324 36316 37380 36318
rect 37548 35756 37604 35812
rect 37212 35084 37268 35140
rect 37548 35532 37604 35588
rect 37324 35026 37380 35028
rect 37324 34974 37326 35026
rect 37326 34974 37378 35026
rect 37378 34974 37380 35026
rect 37324 34972 37380 34974
rect 37436 34242 37492 34244
rect 37436 34190 37438 34242
rect 37438 34190 37490 34242
rect 37490 34190 37492 34242
rect 37436 34188 37492 34190
rect 36988 33964 37044 34020
rect 37548 32508 37604 32564
rect 36988 32396 37044 32452
rect 37324 31666 37380 31668
rect 37324 31614 37326 31666
rect 37326 31614 37378 31666
rect 37378 31614 37380 31666
rect 37324 31612 37380 31614
rect 37436 31554 37492 31556
rect 37436 31502 37438 31554
rect 37438 31502 37490 31554
rect 37490 31502 37492 31554
rect 37436 31500 37492 31502
rect 37212 31052 37268 31108
rect 37548 30492 37604 30548
rect 37884 36258 37940 36260
rect 37884 36206 37886 36258
rect 37886 36206 37938 36258
rect 37938 36206 37940 36258
rect 37884 36204 37940 36206
rect 39116 42588 39172 42644
rect 39900 44156 39956 44212
rect 39228 41916 39284 41972
rect 39340 41580 39396 41636
rect 39676 42194 39732 42196
rect 39676 42142 39678 42194
rect 39678 42142 39730 42194
rect 39730 42142 39732 42194
rect 39676 42140 39732 42142
rect 41020 47234 41076 47236
rect 41020 47182 41022 47234
rect 41022 47182 41074 47234
rect 41074 47182 41076 47234
rect 41020 47180 41076 47182
rect 41020 46674 41076 46676
rect 41020 46622 41022 46674
rect 41022 46622 41074 46674
rect 41074 46622 41076 46674
rect 41020 46620 41076 46622
rect 41916 47458 41972 47460
rect 41916 47406 41918 47458
rect 41918 47406 41970 47458
rect 41970 47406 41972 47458
rect 41916 47404 41972 47406
rect 42140 47458 42196 47460
rect 42140 47406 42142 47458
rect 42142 47406 42194 47458
rect 42194 47406 42196 47458
rect 42140 47404 42196 47406
rect 41356 47234 41412 47236
rect 41356 47182 41358 47234
rect 41358 47182 41410 47234
rect 41410 47182 41412 47234
rect 41356 47180 41412 47182
rect 41356 46620 41412 46676
rect 41580 46060 41636 46116
rect 41692 46172 41748 46228
rect 41468 45388 41524 45444
rect 41132 44434 41188 44436
rect 41132 44382 41134 44434
rect 41134 44382 41186 44434
rect 41186 44382 41188 44434
rect 41132 44380 41188 44382
rect 41356 44994 41412 44996
rect 41356 44942 41358 44994
rect 41358 44942 41410 44994
rect 41410 44942 41412 44994
rect 41356 44940 41412 44942
rect 40460 44044 40516 44100
rect 40348 43148 40404 43204
rect 39676 41692 39732 41748
rect 39004 41132 39060 41188
rect 38668 40572 38724 40628
rect 38332 39394 38388 39396
rect 38332 39342 38334 39394
rect 38334 39342 38386 39394
rect 38386 39342 38388 39394
rect 38332 39340 38388 39342
rect 38332 39004 38388 39060
rect 38444 37212 38500 37268
rect 38780 40908 38836 40964
rect 38892 39452 38948 39508
rect 38892 38780 38948 38836
rect 39004 39228 39060 39284
rect 38892 38556 38948 38612
rect 38892 37884 38948 37940
rect 38892 37660 38948 37716
rect 39228 39676 39284 39732
rect 39228 39340 39284 39396
rect 39116 38668 39172 38724
rect 39228 38892 39284 38948
rect 39004 37436 39060 37492
rect 37996 35868 38052 35924
rect 38668 35810 38724 35812
rect 38668 35758 38670 35810
rect 38670 35758 38722 35810
rect 38722 35758 38724 35810
rect 38668 35756 38724 35758
rect 38556 35644 38612 35700
rect 38108 34748 38164 34804
rect 37772 33234 37828 33236
rect 37772 33182 37774 33234
rect 37774 33182 37826 33234
rect 37826 33182 37828 33234
rect 37772 33180 37828 33182
rect 37996 32956 38052 33012
rect 37660 29932 37716 29988
rect 36988 29708 37044 29764
rect 37660 29708 37716 29764
rect 37884 30156 37940 30212
rect 37996 32508 38052 32564
rect 36988 27916 37044 27972
rect 36988 27074 37044 27076
rect 36988 27022 36990 27074
rect 36990 27022 37042 27074
rect 37042 27022 37044 27074
rect 36988 27020 37044 27022
rect 37436 28476 37492 28532
rect 37548 27634 37604 27636
rect 37548 27582 37550 27634
rect 37550 27582 37602 27634
rect 37602 27582 37604 27634
rect 37548 27580 37604 27582
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34972 25452 35028 25508
rect 35532 25618 35588 25620
rect 35532 25566 35534 25618
rect 35534 25566 35586 25618
rect 35586 25566 35588 25618
rect 35532 25564 35588 25566
rect 35644 25506 35700 25508
rect 35644 25454 35646 25506
rect 35646 25454 35698 25506
rect 35698 25454 35700 25506
rect 35644 25452 35700 25454
rect 34188 24556 34244 24612
rect 34860 24162 34916 24164
rect 34860 24110 34862 24162
rect 34862 24110 34914 24162
rect 34914 24110 34916 24162
rect 34860 24108 34916 24110
rect 34412 23436 34468 23492
rect 33964 21868 34020 21924
rect 34188 22876 34244 22932
rect 34188 22370 34244 22372
rect 34188 22318 34190 22370
rect 34190 22318 34242 22370
rect 34242 22318 34244 22370
rect 34188 22316 34244 22318
rect 34188 21868 34244 21924
rect 33852 21420 33908 21476
rect 33516 19404 33572 19460
rect 33628 20636 33684 20692
rect 34076 21362 34132 21364
rect 34076 21310 34078 21362
rect 34078 21310 34130 21362
rect 34130 21310 34132 21362
rect 34076 21308 34132 21310
rect 34188 21084 34244 21140
rect 33852 20188 33908 20244
rect 32844 18844 32900 18900
rect 32508 18508 32564 18564
rect 31836 18172 31892 18228
rect 31724 17724 31780 17780
rect 30268 17276 30324 17332
rect 33180 18396 33236 18452
rect 33852 18956 33908 19012
rect 34524 23324 34580 23380
rect 34524 22930 34580 22932
rect 34524 22878 34526 22930
rect 34526 22878 34578 22930
rect 34578 22878 34580 22930
rect 34524 22876 34580 22878
rect 34300 20524 34356 20580
rect 34300 20188 34356 20244
rect 34188 20018 34244 20020
rect 34188 19966 34190 20018
rect 34190 19966 34242 20018
rect 34242 19966 34244 20018
rect 34188 19964 34244 19966
rect 34972 23938 35028 23940
rect 34972 23886 34974 23938
rect 34974 23886 35026 23938
rect 35026 23886 35028 23938
rect 34972 23884 35028 23886
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 23938 35252 23940
rect 35196 23886 35198 23938
rect 35198 23886 35250 23938
rect 35250 23886 35252 23938
rect 35196 23884 35252 23886
rect 36204 26012 36260 26068
rect 36428 25394 36484 25396
rect 36428 25342 36430 25394
rect 36430 25342 36482 25394
rect 36482 25342 36484 25394
rect 36428 25340 36484 25342
rect 35980 25116 36036 25172
rect 36316 25228 36372 25284
rect 36428 24556 36484 24612
rect 36092 24050 36148 24052
rect 36092 23998 36094 24050
rect 36094 23998 36146 24050
rect 36146 23998 36148 24050
rect 36092 23996 36148 23998
rect 35868 23772 35924 23828
rect 35084 23378 35140 23380
rect 35084 23326 35086 23378
rect 35086 23326 35138 23378
rect 35138 23326 35140 23378
rect 35084 23324 35140 23326
rect 34748 23042 34804 23044
rect 34748 22990 34750 23042
rect 34750 22990 34802 23042
rect 34802 22990 34804 23042
rect 34748 22988 34804 22990
rect 34636 22482 34692 22484
rect 34636 22430 34638 22482
rect 34638 22430 34690 22482
rect 34690 22430 34692 22482
rect 34636 22428 34692 22430
rect 34524 19964 34580 20020
rect 34636 21474 34692 21476
rect 34636 21422 34638 21474
rect 34638 21422 34690 21474
rect 34690 21422 34692 21474
rect 34636 21420 34692 21422
rect 36764 25788 36820 25844
rect 36652 25452 36708 25508
rect 35420 23100 35476 23156
rect 35980 23042 36036 23044
rect 35980 22990 35982 23042
rect 35982 22990 36034 23042
rect 36034 22990 36036 23042
rect 35980 22988 36036 22990
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35644 22764 35700 22820
rect 37212 25506 37268 25508
rect 37212 25454 37214 25506
rect 37214 25454 37266 25506
rect 37266 25454 37268 25506
rect 37212 25452 37268 25454
rect 36988 25228 37044 25284
rect 37100 24610 37156 24612
rect 37100 24558 37102 24610
rect 37102 24558 37154 24610
rect 37154 24558 37156 24610
rect 37100 24556 37156 24558
rect 36876 23884 36932 23940
rect 37660 26796 37716 26852
rect 37660 25788 37716 25844
rect 39452 40514 39508 40516
rect 39452 40462 39454 40514
rect 39454 40462 39506 40514
rect 39506 40462 39508 40514
rect 39452 40460 39508 40462
rect 38556 32508 38612 32564
rect 38668 35420 38724 35476
rect 38444 32396 38500 32452
rect 38108 31724 38164 31780
rect 38332 31554 38388 31556
rect 38332 31502 38334 31554
rect 38334 31502 38386 31554
rect 38386 31502 38388 31554
rect 38332 31500 38388 31502
rect 38220 31388 38276 31444
rect 38444 31276 38500 31332
rect 38892 35084 38948 35140
rect 38892 32562 38948 32564
rect 38892 32510 38894 32562
rect 38894 32510 38946 32562
rect 38946 32510 38948 32562
rect 38892 32508 38948 32510
rect 38668 31052 38724 31108
rect 38108 30268 38164 30324
rect 38892 31612 38948 31668
rect 40348 42476 40404 42532
rect 40236 41858 40292 41860
rect 40236 41806 40238 41858
rect 40238 41806 40290 41858
rect 40290 41806 40292 41858
rect 40236 41804 40292 41806
rect 41020 43820 41076 43876
rect 40796 42252 40852 42308
rect 41804 45890 41860 45892
rect 41804 45838 41806 45890
rect 41806 45838 41858 45890
rect 41858 45838 41860 45890
rect 41804 45836 41860 45838
rect 41468 43820 41524 43876
rect 41692 43426 41748 43428
rect 41692 43374 41694 43426
rect 41694 43374 41746 43426
rect 41746 43374 41748 43426
rect 41692 43372 41748 43374
rect 48188 47964 48244 48020
rect 45388 47682 45444 47684
rect 45388 47630 45390 47682
rect 45390 47630 45442 47682
rect 45442 47630 45444 47682
rect 45388 47628 45444 47630
rect 47516 47628 47572 47684
rect 42588 45836 42644 45892
rect 42700 44940 42756 44996
rect 42588 44882 42644 44884
rect 42588 44830 42590 44882
rect 42590 44830 42642 44882
rect 42642 44830 42644 44882
rect 42588 44828 42644 44830
rect 42476 44492 42532 44548
rect 42364 44380 42420 44436
rect 43036 45948 43092 46004
rect 44156 47404 44212 47460
rect 42924 44268 42980 44324
rect 43036 45500 43092 45556
rect 43260 44940 43316 44996
rect 42140 43260 42196 43316
rect 42588 43372 42644 43428
rect 41804 42700 41860 42756
rect 41244 42140 41300 42196
rect 41132 41580 41188 41636
rect 40460 41132 40516 41188
rect 41244 41132 41300 41188
rect 42476 42754 42532 42756
rect 42476 42702 42478 42754
rect 42478 42702 42530 42754
rect 42530 42702 42532 42754
rect 42476 42700 42532 42702
rect 42812 42754 42868 42756
rect 42812 42702 42814 42754
rect 42814 42702 42866 42754
rect 42866 42702 42868 42754
rect 42812 42700 42868 42702
rect 42700 42588 42756 42644
rect 41804 41858 41860 41860
rect 41804 41806 41806 41858
rect 41806 41806 41858 41858
rect 41858 41806 41860 41858
rect 41804 41804 41860 41806
rect 41020 40626 41076 40628
rect 41020 40574 41022 40626
rect 41022 40574 41074 40626
rect 41074 40574 41076 40626
rect 41020 40572 41076 40574
rect 39676 40348 39732 40404
rect 41468 40290 41524 40292
rect 41468 40238 41470 40290
rect 41470 40238 41522 40290
rect 41522 40238 41524 40290
rect 41468 40236 41524 40238
rect 39788 39788 39844 39844
rect 41244 39788 41300 39844
rect 41020 39228 41076 39284
rect 40684 39116 40740 39172
rect 40012 38892 40068 38948
rect 39900 37660 39956 37716
rect 40236 38722 40292 38724
rect 40236 38670 40238 38722
rect 40238 38670 40290 38722
rect 40290 38670 40292 38722
rect 40236 38668 40292 38670
rect 40348 38444 40404 38500
rect 39676 37490 39732 37492
rect 39676 37438 39678 37490
rect 39678 37438 39730 37490
rect 39730 37438 39732 37490
rect 39676 37436 39732 37438
rect 40236 37996 40292 38052
rect 39564 37324 39620 37380
rect 39452 35586 39508 35588
rect 39452 35534 39454 35586
rect 39454 35534 39506 35586
rect 39506 35534 39508 35586
rect 39452 35532 39508 35534
rect 39676 35756 39732 35812
rect 39340 34972 39396 35028
rect 39676 35196 39732 35252
rect 39564 33852 39620 33908
rect 39228 32956 39284 33012
rect 40012 37266 40068 37268
rect 40012 37214 40014 37266
rect 40014 37214 40066 37266
rect 40066 37214 40068 37266
rect 40012 37212 40068 37214
rect 39900 37154 39956 37156
rect 39900 37102 39902 37154
rect 39902 37102 39954 37154
rect 39954 37102 39956 37154
rect 39900 37100 39956 37102
rect 39900 35084 39956 35140
rect 39788 34748 39844 34804
rect 40124 35980 40180 36036
rect 40236 35922 40292 35924
rect 40236 35870 40238 35922
rect 40238 35870 40290 35922
rect 40290 35870 40292 35922
rect 40236 35868 40292 35870
rect 41132 39116 41188 39172
rect 41356 39676 41412 39732
rect 41020 37884 41076 37940
rect 41244 37772 41300 37828
rect 40908 37324 40964 37380
rect 40908 37154 40964 37156
rect 40908 37102 40910 37154
rect 40910 37102 40962 37154
rect 40962 37102 40964 37154
rect 40908 37100 40964 37102
rect 40908 36540 40964 36596
rect 41804 40514 41860 40516
rect 41804 40462 41806 40514
rect 41806 40462 41858 40514
rect 41858 40462 41860 40514
rect 41804 40460 41860 40462
rect 42364 41746 42420 41748
rect 42364 41694 42366 41746
rect 42366 41694 42418 41746
rect 42418 41694 42420 41746
rect 42364 41692 42420 41694
rect 42252 41580 42308 41636
rect 42140 41186 42196 41188
rect 42140 41134 42142 41186
rect 42142 41134 42194 41186
rect 42194 41134 42196 41186
rect 42140 41132 42196 41134
rect 42364 40908 42420 40964
rect 41916 40178 41972 40180
rect 41916 40126 41918 40178
rect 41918 40126 41970 40178
rect 41970 40126 41972 40178
rect 41916 40124 41972 40126
rect 41804 39116 41860 39172
rect 41580 37938 41636 37940
rect 41580 37886 41582 37938
rect 41582 37886 41634 37938
rect 41634 37886 41636 37938
rect 41580 37884 41636 37886
rect 41356 35756 41412 35812
rect 40348 35474 40404 35476
rect 40348 35422 40350 35474
rect 40350 35422 40402 35474
rect 40402 35422 40404 35474
rect 40348 35420 40404 35422
rect 40236 35196 40292 35252
rect 40236 34914 40292 34916
rect 40236 34862 40238 34914
rect 40238 34862 40290 34914
rect 40290 34862 40292 34914
rect 40236 34860 40292 34862
rect 41020 34914 41076 34916
rect 41020 34862 41022 34914
rect 41022 34862 41074 34914
rect 41074 34862 41076 34914
rect 41020 34860 41076 34862
rect 39900 33404 39956 33460
rect 39116 31388 39172 31444
rect 39340 31612 39396 31668
rect 38220 30156 38276 30212
rect 37996 29372 38052 29428
rect 37996 27692 38052 27748
rect 38108 29932 38164 29988
rect 38108 28140 38164 28196
rect 38892 31276 38948 31332
rect 38444 28700 38500 28756
rect 38332 28476 38388 28532
rect 38668 29148 38724 29204
rect 37996 26962 38052 26964
rect 37996 26910 37998 26962
rect 37998 26910 38050 26962
rect 38050 26910 38052 26962
rect 37996 26908 38052 26910
rect 38668 27692 38724 27748
rect 37884 25900 37940 25956
rect 37324 23996 37380 24052
rect 37436 25452 37492 25508
rect 37548 23884 37604 23940
rect 37324 22876 37380 22932
rect 36876 22764 36932 22820
rect 36764 22428 36820 22484
rect 36204 22316 36260 22372
rect 35980 21810 36036 21812
rect 35980 21758 35982 21810
rect 35982 21758 36034 21810
rect 36034 21758 36036 21810
rect 35980 21756 36036 21758
rect 35084 21586 35140 21588
rect 35084 21534 35086 21586
rect 35086 21534 35138 21586
rect 35138 21534 35140 21586
rect 35084 21532 35140 21534
rect 35756 21420 35812 21476
rect 36428 22146 36484 22148
rect 36428 22094 36430 22146
rect 36430 22094 36482 22146
rect 36482 22094 36484 22146
rect 36428 22092 36484 22094
rect 36092 21420 36148 21476
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35868 21362 35924 21364
rect 35868 21310 35870 21362
rect 35870 21310 35922 21362
rect 35922 21310 35924 21362
rect 35868 21308 35924 21310
rect 35532 20972 35588 21028
rect 35980 20972 36036 21028
rect 35196 20748 35252 20804
rect 36428 21420 36484 21476
rect 34748 20578 34804 20580
rect 34748 20526 34750 20578
rect 34750 20526 34802 20578
rect 34802 20526 34804 20578
rect 34748 20524 34804 20526
rect 35756 20524 35812 20580
rect 35868 20188 35924 20244
rect 34636 19740 34692 19796
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34636 19180 34692 19236
rect 35420 19180 35476 19236
rect 32844 17778 32900 17780
rect 32844 17726 32846 17778
rect 32846 17726 32898 17778
rect 32898 17726 32900 17778
rect 32844 17724 32900 17726
rect 32284 17500 32340 17556
rect 30268 16994 30324 16996
rect 30268 16942 30270 16994
rect 30270 16942 30322 16994
rect 30322 16942 30324 16994
rect 30268 16940 30324 16942
rect 30604 16940 30660 16996
rect 30156 16770 30212 16772
rect 30156 16718 30158 16770
rect 30158 16718 30210 16770
rect 30210 16718 30212 16770
rect 30156 16716 30212 16718
rect 30156 16380 30212 16436
rect 32508 17612 32564 17668
rect 31276 16828 31332 16884
rect 31500 16882 31556 16884
rect 31500 16830 31502 16882
rect 31502 16830 31554 16882
rect 31554 16830 31556 16882
rect 31500 16828 31556 16830
rect 31724 16716 31780 16772
rect 30828 15484 30884 15540
rect 30604 15426 30660 15428
rect 30604 15374 30606 15426
rect 30606 15374 30658 15426
rect 30658 15374 30660 15426
rect 30604 15372 30660 15374
rect 30828 15314 30884 15316
rect 30828 15262 30830 15314
rect 30830 15262 30882 15314
rect 30882 15262 30884 15314
rect 30828 15260 30884 15262
rect 30716 15148 30772 15204
rect 30156 14476 30212 14532
rect 29932 13634 29988 13636
rect 29932 13582 29934 13634
rect 29934 13582 29986 13634
rect 29986 13582 29988 13634
rect 29932 13580 29988 13582
rect 29708 12178 29764 12180
rect 29708 12126 29710 12178
rect 29710 12126 29762 12178
rect 29762 12126 29764 12178
rect 29708 12124 29764 12126
rect 29148 10108 29204 10164
rect 28476 9772 28532 9828
rect 29372 9660 29428 9716
rect 29932 12962 29988 12964
rect 29932 12910 29934 12962
rect 29934 12910 29986 12962
rect 29986 12910 29988 12962
rect 29932 12908 29988 12910
rect 30380 13020 30436 13076
rect 32284 16380 32340 16436
rect 33068 17724 33124 17780
rect 33964 18450 34020 18452
rect 33964 18398 33966 18450
rect 33966 18398 34018 18450
rect 34018 18398 34020 18450
rect 33964 18396 34020 18398
rect 33516 17666 33572 17668
rect 33516 17614 33518 17666
rect 33518 17614 33570 17666
rect 33570 17614 33572 17666
rect 33516 17612 33572 17614
rect 34076 17836 34132 17892
rect 33964 17778 34020 17780
rect 33964 17726 33966 17778
rect 33966 17726 34018 17778
rect 34018 17726 34020 17778
rect 33964 17724 34020 17726
rect 33292 17554 33348 17556
rect 33292 17502 33294 17554
rect 33294 17502 33346 17554
rect 33346 17502 33348 17554
rect 33292 17500 33348 17502
rect 33516 17388 33572 17444
rect 33404 17164 33460 17220
rect 34076 17388 34132 17444
rect 33964 16994 34020 16996
rect 33964 16942 33966 16994
rect 33966 16942 34018 16994
rect 34018 16942 34020 16994
rect 33964 16940 34020 16942
rect 34412 18956 34468 19012
rect 34300 17554 34356 17556
rect 34300 17502 34302 17554
rect 34302 17502 34354 17554
rect 34354 17502 34356 17554
rect 34300 17500 34356 17502
rect 35868 18844 35924 18900
rect 34524 18284 34580 18340
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34412 17388 34468 17444
rect 33180 16828 33236 16884
rect 35420 17554 35476 17556
rect 35420 17502 35422 17554
rect 35422 17502 35474 17554
rect 35474 17502 35476 17554
rect 35420 17500 35476 17502
rect 34524 16828 34580 16884
rect 35532 17276 35588 17332
rect 35196 16716 35252 16772
rect 32060 15372 32116 15428
rect 31724 14028 31780 14084
rect 31500 13692 31556 13748
rect 31388 13468 31444 13524
rect 31052 12908 31108 12964
rect 30156 12290 30212 12292
rect 30156 12238 30158 12290
rect 30158 12238 30210 12290
rect 30210 12238 30212 12290
rect 30156 12236 30212 12238
rect 31612 13020 31668 13076
rect 31052 12290 31108 12292
rect 31052 12238 31054 12290
rect 31054 12238 31106 12290
rect 31106 12238 31108 12290
rect 31052 12236 31108 12238
rect 30044 11676 30100 11732
rect 30268 11676 30324 11732
rect 30940 11506 30996 11508
rect 30940 11454 30942 11506
rect 30942 11454 30994 11506
rect 30994 11454 30996 11506
rect 30940 11452 30996 11454
rect 29820 11228 29876 11284
rect 30044 11116 30100 11172
rect 30044 10668 30100 10724
rect 32284 15484 32340 15540
rect 31948 15090 32004 15092
rect 31948 15038 31950 15090
rect 31950 15038 32002 15090
rect 32002 15038 32004 15090
rect 31948 15036 32004 15038
rect 31836 13804 31892 13860
rect 31836 13356 31892 13412
rect 32508 14924 32564 14980
rect 32732 15260 32788 15316
rect 32732 14530 32788 14532
rect 32732 14478 32734 14530
rect 32734 14478 32786 14530
rect 32786 14478 32788 14530
rect 32732 14476 32788 14478
rect 32620 13916 32676 13972
rect 32508 13746 32564 13748
rect 32508 13694 32510 13746
rect 32510 13694 32562 13746
rect 32562 13694 32564 13746
rect 32508 13692 32564 13694
rect 32732 14140 32788 14196
rect 32732 13692 32788 13748
rect 32956 15372 33012 15428
rect 33068 15202 33124 15204
rect 33068 15150 33070 15202
rect 33070 15150 33122 15202
rect 33122 15150 33124 15202
rect 33068 15148 33124 15150
rect 33068 13746 33124 13748
rect 33068 13694 33070 13746
rect 33070 13694 33122 13746
rect 33122 13694 33124 13746
rect 33068 13692 33124 13694
rect 33404 16658 33460 16660
rect 33404 16606 33406 16658
rect 33406 16606 33458 16658
rect 33458 16606 33460 16658
rect 33404 16604 33460 16606
rect 33516 15314 33572 15316
rect 33516 15262 33518 15314
rect 33518 15262 33570 15314
rect 33570 15262 33572 15314
rect 33516 15260 33572 15262
rect 33852 15484 33908 15540
rect 33852 15148 33908 15204
rect 33516 14924 33572 14980
rect 33516 14700 33572 14756
rect 33292 13244 33348 13300
rect 33740 13858 33796 13860
rect 33740 13806 33742 13858
rect 33742 13806 33794 13858
rect 33794 13806 33796 13858
rect 33740 13804 33796 13806
rect 33516 13468 33572 13524
rect 33292 12962 33348 12964
rect 33292 12910 33294 12962
rect 33294 12910 33346 12962
rect 33346 12910 33348 12962
rect 33292 12908 33348 12910
rect 33404 12796 33460 12852
rect 31948 12124 32004 12180
rect 31276 11340 31332 11396
rect 28924 9042 28980 9044
rect 28924 8990 28926 9042
rect 28926 8990 28978 9042
rect 28978 8990 28980 9042
rect 28924 8988 28980 8990
rect 28588 8764 28644 8820
rect 28140 8316 28196 8372
rect 26572 8146 26628 8148
rect 26572 8094 26574 8146
rect 26574 8094 26626 8146
rect 26626 8094 26628 8146
rect 26572 8092 26628 8094
rect 27580 8034 27636 8036
rect 27580 7982 27582 8034
rect 27582 7982 27634 8034
rect 27634 7982 27636 8034
rect 27580 7980 27636 7982
rect 26124 7756 26180 7812
rect 26012 7420 26068 7476
rect 25676 4396 25732 4452
rect 28364 8258 28420 8260
rect 28364 8206 28366 8258
rect 28366 8206 28418 8258
rect 28418 8206 28420 8258
rect 28364 8204 28420 8206
rect 28700 8316 28756 8372
rect 29372 9324 29428 9380
rect 29148 8818 29204 8820
rect 29148 8766 29150 8818
rect 29150 8766 29202 8818
rect 29202 8766 29204 8818
rect 29148 8764 29204 8766
rect 28924 8204 28980 8260
rect 28476 8034 28532 8036
rect 28476 7982 28478 8034
rect 28478 7982 28530 8034
rect 28530 7982 28532 8034
rect 28476 7980 28532 7982
rect 27132 7420 27188 7476
rect 26460 7308 26516 7364
rect 26908 6524 26964 6580
rect 26572 5682 26628 5684
rect 26572 5630 26574 5682
rect 26574 5630 26626 5682
rect 26626 5630 26628 5682
rect 26572 5628 26628 5630
rect 27020 5628 27076 5684
rect 26460 5068 26516 5124
rect 26348 4844 26404 4900
rect 23100 4284 23156 4340
rect 23324 4226 23380 4228
rect 23324 4174 23326 4226
rect 23326 4174 23378 4226
rect 23378 4174 23380 4226
rect 23324 4172 23380 4174
rect 25452 4338 25508 4340
rect 25452 4286 25454 4338
rect 25454 4286 25506 4338
rect 25506 4286 25508 4338
rect 25452 4284 25508 4286
rect 25340 4226 25396 4228
rect 25340 4174 25342 4226
rect 25342 4174 25394 4226
rect 25394 4174 25396 4226
rect 25340 4172 25396 4174
rect 24556 4114 24612 4116
rect 24556 4062 24558 4114
rect 24558 4062 24610 4114
rect 24610 4062 24612 4114
rect 24556 4060 24612 4062
rect 26124 4114 26180 4116
rect 26124 4062 26126 4114
rect 26126 4062 26178 4114
rect 26178 4062 26180 4114
rect 26124 4060 26180 4062
rect 24444 3276 24500 3332
rect 26684 4450 26740 4452
rect 26684 4398 26686 4450
rect 26686 4398 26738 4450
rect 26738 4398 26740 4450
rect 26684 4396 26740 4398
rect 28476 7474 28532 7476
rect 28476 7422 28478 7474
rect 28478 7422 28530 7474
rect 28530 7422 28532 7474
rect 28476 7420 28532 7422
rect 29260 7420 29316 7476
rect 28028 6524 28084 6580
rect 29036 6578 29092 6580
rect 29036 6526 29038 6578
rect 29038 6526 29090 6578
rect 29090 6526 29092 6578
rect 29036 6524 29092 6526
rect 28588 6412 28644 6468
rect 27468 5628 27524 5684
rect 27580 5122 27636 5124
rect 27580 5070 27582 5122
rect 27582 5070 27634 5122
rect 27634 5070 27636 5122
rect 27580 5068 27636 5070
rect 27804 5906 27860 5908
rect 27804 5854 27806 5906
rect 27806 5854 27858 5906
rect 27858 5854 27860 5906
rect 27804 5852 27860 5854
rect 29820 9042 29876 9044
rect 29820 8990 29822 9042
rect 29822 8990 29874 9042
rect 29874 8990 29876 9042
rect 29820 8988 29876 8990
rect 30044 9042 30100 9044
rect 30044 8990 30046 9042
rect 30046 8990 30098 9042
rect 30098 8990 30100 9042
rect 30044 8988 30100 8990
rect 30156 8764 30212 8820
rect 29708 7980 29764 8036
rect 30268 7980 30324 8036
rect 29932 7420 29988 7476
rect 30940 9826 30996 9828
rect 30940 9774 30942 9826
rect 30942 9774 30994 9826
rect 30994 9774 30996 9826
rect 30940 9772 30996 9774
rect 31836 11788 31892 11844
rect 31388 11228 31444 11284
rect 31948 11676 32004 11732
rect 31724 11564 31780 11620
rect 32396 12290 32452 12292
rect 32396 12238 32398 12290
rect 32398 12238 32450 12290
rect 32450 12238 32452 12290
rect 32396 12236 32452 12238
rect 32844 12124 32900 12180
rect 32284 11564 32340 11620
rect 31836 11116 31892 11172
rect 31724 10834 31780 10836
rect 31724 10782 31726 10834
rect 31726 10782 31778 10834
rect 31778 10782 31780 10834
rect 31724 10780 31780 10782
rect 32508 11676 32564 11732
rect 32508 11116 32564 11172
rect 31388 10610 31444 10612
rect 31388 10558 31390 10610
rect 31390 10558 31442 10610
rect 31442 10558 31444 10610
rect 31388 10556 31444 10558
rect 32172 10610 32228 10612
rect 32172 10558 32174 10610
rect 32174 10558 32226 10610
rect 32226 10558 32228 10610
rect 32172 10556 32228 10558
rect 32172 10108 32228 10164
rect 31500 9266 31556 9268
rect 31500 9214 31502 9266
rect 31502 9214 31554 9266
rect 31554 9214 31556 9266
rect 31500 9212 31556 9214
rect 31052 9154 31108 9156
rect 31052 9102 31054 9154
rect 31054 9102 31106 9154
rect 31106 9102 31108 9154
rect 31052 9100 31108 9102
rect 30716 9042 30772 9044
rect 30716 8990 30718 9042
rect 30718 8990 30770 9042
rect 30770 8990 30772 9042
rect 30716 8988 30772 8990
rect 31500 8818 31556 8820
rect 31500 8766 31502 8818
rect 31502 8766 31554 8818
rect 31554 8766 31556 8818
rect 31500 8764 31556 8766
rect 34188 15036 34244 15092
rect 34524 15148 34580 15204
rect 34300 14588 34356 14644
rect 34636 14028 34692 14084
rect 34412 13916 34468 13972
rect 34748 13634 34804 13636
rect 34748 13582 34750 13634
rect 34750 13582 34802 13634
rect 34802 13582 34804 13634
rect 34748 13580 34804 13582
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35308 15820 35364 15876
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35532 14700 35588 14756
rect 35308 14476 35364 14532
rect 34972 13356 35028 13412
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35756 17442 35812 17444
rect 35756 17390 35758 17442
rect 35758 17390 35810 17442
rect 35810 17390 35812 17442
rect 35756 17388 35812 17390
rect 36764 21308 36820 21364
rect 35868 17276 35924 17332
rect 35980 18396 36036 18452
rect 35756 16994 35812 16996
rect 35756 16942 35758 16994
rect 35758 16942 35810 16994
rect 35810 16942 35812 16994
rect 35756 16940 35812 16942
rect 36092 18338 36148 18340
rect 36092 18286 36094 18338
rect 36094 18286 36146 18338
rect 36146 18286 36148 18338
rect 36092 18284 36148 18286
rect 36204 17948 36260 18004
rect 36092 17836 36148 17892
rect 37100 22258 37156 22260
rect 37100 22206 37102 22258
rect 37102 22206 37154 22258
rect 37154 22206 37156 22258
rect 37100 22204 37156 22206
rect 36988 21756 37044 21812
rect 37212 22092 37268 22148
rect 37324 21868 37380 21924
rect 37548 21756 37604 21812
rect 36988 20748 37044 20804
rect 36876 18508 36932 18564
rect 36988 20076 37044 20132
rect 36540 18226 36596 18228
rect 36540 18174 36542 18226
rect 36542 18174 36594 18226
rect 36594 18174 36596 18226
rect 36540 18172 36596 18174
rect 36316 17500 36372 17556
rect 36428 17388 36484 17444
rect 36540 16940 36596 16996
rect 36988 18284 37044 18340
rect 36652 16044 36708 16100
rect 36876 17500 36932 17556
rect 37324 20802 37380 20804
rect 37324 20750 37326 20802
rect 37326 20750 37378 20802
rect 37378 20750 37380 20802
rect 37324 20748 37380 20750
rect 37548 20636 37604 20692
rect 37436 19516 37492 19572
rect 37548 18562 37604 18564
rect 37548 18510 37550 18562
rect 37550 18510 37602 18562
rect 37602 18510 37604 18562
rect 37548 18508 37604 18510
rect 37212 17612 37268 17668
rect 37324 18172 37380 18228
rect 37772 25506 37828 25508
rect 37772 25454 37774 25506
rect 37774 25454 37826 25506
rect 37826 25454 37828 25506
rect 37772 25452 37828 25454
rect 37772 25228 37828 25284
rect 38220 25900 38276 25956
rect 38108 25452 38164 25508
rect 38220 25394 38276 25396
rect 38220 25342 38222 25394
rect 38222 25342 38274 25394
rect 38274 25342 38276 25394
rect 38220 25340 38276 25342
rect 37884 23884 37940 23940
rect 37772 23772 37828 23828
rect 38332 25228 38388 25284
rect 38556 23938 38612 23940
rect 38556 23886 38558 23938
rect 38558 23886 38610 23938
rect 38610 23886 38612 23938
rect 38556 23884 38612 23886
rect 37772 23436 37828 23492
rect 37884 21196 37940 21252
rect 37884 20188 37940 20244
rect 37660 18060 37716 18116
rect 37884 19516 37940 19572
rect 37548 16940 37604 16996
rect 37660 17164 37716 17220
rect 37436 16770 37492 16772
rect 37436 16718 37438 16770
rect 37438 16718 37490 16770
rect 37490 16718 37492 16770
rect 37436 16716 37492 16718
rect 36988 15820 37044 15876
rect 36652 14812 36708 14868
rect 35868 14476 35924 14532
rect 34860 13132 34916 13188
rect 34300 12796 34356 12852
rect 33964 11676 34020 11732
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 33068 11228 33124 11284
rect 33404 11004 33460 11060
rect 32732 9660 32788 9716
rect 36092 13356 36148 13412
rect 36316 12962 36372 12964
rect 36316 12910 36318 12962
rect 36318 12910 36370 12962
rect 36370 12910 36372 12962
rect 36316 12908 36372 12910
rect 36540 13020 36596 13076
rect 37324 16098 37380 16100
rect 37324 16046 37326 16098
rect 37326 16046 37378 16098
rect 37378 16046 37380 16098
rect 37324 16044 37380 16046
rect 37436 15820 37492 15876
rect 37324 15596 37380 15652
rect 37212 14364 37268 14420
rect 36428 12572 36484 12628
rect 35756 12124 35812 12180
rect 39004 31052 39060 31108
rect 38892 26572 38948 26628
rect 39116 30098 39172 30100
rect 39116 30046 39118 30098
rect 39118 30046 39170 30098
rect 39170 30046 39172 30098
rect 39116 30044 39172 30046
rect 39676 31554 39732 31556
rect 39676 31502 39678 31554
rect 39678 31502 39730 31554
rect 39730 31502 39732 31554
rect 39676 31500 39732 31502
rect 39676 30268 39732 30324
rect 39340 27692 39396 27748
rect 39116 27132 39172 27188
rect 40460 33458 40516 33460
rect 40460 33406 40462 33458
rect 40462 33406 40514 33458
rect 40514 33406 40516 33458
rect 40460 33404 40516 33406
rect 40460 32172 40516 32228
rect 40572 30268 40628 30324
rect 40796 34188 40852 34244
rect 41692 36370 41748 36372
rect 41692 36318 41694 36370
rect 41694 36318 41746 36370
rect 41746 36318 41748 36370
rect 41692 36316 41748 36318
rect 41468 35644 41524 35700
rect 42028 38722 42084 38724
rect 42028 38670 42030 38722
rect 42030 38670 42082 38722
rect 42082 38670 42084 38722
rect 42028 38668 42084 38670
rect 43484 45666 43540 45668
rect 43484 45614 43486 45666
rect 43486 45614 43538 45666
rect 43538 45614 43540 45666
rect 43484 45612 43540 45614
rect 44380 46674 44436 46676
rect 44380 46622 44382 46674
rect 44382 46622 44434 46674
rect 44434 46622 44436 46674
rect 44380 46620 44436 46622
rect 44268 46172 44324 46228
rect 43932 45890 43988 45892
rect 43932 45838 43934 45890
rect 43934 45838 43986 45890
rect 43986 45838 43988 45890
rect 43932 45836 43988 45838
rect 44380 45836 44436 45892
rect 43820 45500 43876 45556
rect 43820 44322 43876 44324
rect 43820 44270 43822 44322
rect 43822 44270 43874 44322
rect 43874 44270 43876 44322
rect 43820 44268 43876 44270
rect 43596 44156 43652 44212
rect 44268 44210 44324 44212
rect 44268 44158 44270 44210
rect 44270 44158 44322 44210
rect 44322 44158 44324 44210
rect 44268 44156 44324 44158
rect 44044 44098 44100 44100
rect 44044 44046 44046 44098
rect 44046 44046 44098 44098
rect 44098 44046 44100 44098
rect 44044 44044 44100 44046
rect 43932 43708 43988 43764
rect 44492 43596 44548 43652
rect 43372 43148 43428 43204
rect 44268 43260 44324 43316
rect 43596 42700 43652 42756
rect 43596 42364 43652 42420
rect 43260 42082 43316 42084
rect 43260 42030 43262 42082
rect 43262 42030 43314 42082
rect 43314 42030 43316 42082
rect 43260 42028 43316 42030
rect 44156 42140 44212 42196
rect 43036 41970 43092 41972
rect 43036 41918 43038 41970
rect 43038 41918 43090 41970
rect 43090 41918 43092 41970
rect 43036 41916 43092 41918
rect 42588 40460 42644 40516
rect 42700 40348 42756 40404
rect 42588 39340 42644 39396
rect 42252 38108 42308 38164
rect 41132 34354 41188 34356
rect 41132 34302 41134 34354
rect 41134 34302 41186 34354
rect 41186 34302 41188 34354
rect 41132 34300 41188 34302
rect 41020 33516 41076 33572
rect 41244 33404 41300 33460
rect 41468 33516 41524 33572
rect 40908 33180 40964 33236
rect 41020 32450 41076 32452
rect 41020 32398 41022 32450
rect 41022 32398 41074 32450
rect 41074 32398 41076 32450
rect 41020 32396 41076 32398
rect 40908 32172 40964 32228
rect 41356 31554 41412 31556
rect 41356 31502 41358 31554
rect 41358 31502 41410 31554
rect 41410 31502 41412 31554
rect 41356 31500 41412 31502
rect 41468 31388 41524 31444
rect 41244 30156 41300 30212
rect 40124 29708 40180 29764
rect 40460 29708 40516 29764
rect 40796 30044 40852 30100
rect 40348 29650 40404 29652
rect 40348 29598 40350 29650
rect 40350 29598 40402 29650
rect 40402 29598 40404 29650
rect 40348 29596 40404 29598
rect 40012 29484 40068 29540
rect 39900 28588 39956 28644
rect 40012 29148 40068 29204
rect 39900 27692 39956 27748
rect 41132 29708 41188 29764
rect 40460 28700 40516 28756
rect 40908 29484 40964 29540
rect 41468 30268 41524 30324
rect 41692 31778 41748 31780
rect 41692 31726 41694 31778
rect 41694 31726 41746 31778
rect 41746 31726 41748 31778
rect 41692 31724 41748 31726
rect 41916 37324 41972 37380
rect 41916 34860 41972 34916
rect 42700 38668 42756 38724
rect 42924 41132 42980 41188
rect 42924 40402 42980 40404
rect 42924 40350 42926 40402
rect 42926 40350 42978 40402
rect 42978 40350 42980 40402
rect 42924 40348 42980 40350
rect 43596 41468 43652 41524
rect 43372 40572 43428 40628
rect 42812 37772 42868 37828
rect 42476 36428 42532 36484
rect 42700 36988 42756 37044
rect 42028 34636 42084 34692
rect 42140 34188 42196 34244
rect 42140 33740 42196 33796
rect 42588 33458 42644 33460
rect 42588 33406 42590 33458
rect 42590 33406 42642 33458
rect 42642 33406 42644 33458
rect 42588 33404 42644 33406
rect 42476 33180 42532 33236
rect 42588 31724 42644 31780
rect 42252 31612 42308 31668
rect 41692 31276 41748 31332
rect 42364 31500 42420 31556
rect 41580 29820 41636 29876
rect 41244 28812 41300 28868
rect 41468 29260 41524 29316
rect 40908 28700 40964 28756
rect 41356 28588 41412 28644
rect 40348 28530 40404 28532
rect 40348 28478 40350 28530
rect 40350 28478 40402 28530
rect 40402 28478 40404 28530
rect 40348 28476 40404 28478
rect 38892 25394 38948 25396
rect 38892 25342 38894 25394
rect 38894 25342 38946 25394
rect 38946 25342 38948 25394
rect 38892 25340 38948 25342
rect 39004 23660 39060 23716
rect 38892 23378 38948 23380
rect 38892 23326 38894 23378
rect 38894 23326 38946 23378
rect 38946 23326 38948 23378
rect 38892 23324 38948 23326
rect 38220 23266 38276 23268
rect 38220 23214 38222 23266
rect 38222 23214 38274 23266
rect 38274 23214 38276 23266
rect 38220 23212 38276 23214
rect 38332 23154 38388 23156
rect 38332 23102 38334 23154
rect 38334 23102 38386 23154
rect 38386 23102 38388 23154
rect 38332 23100 38388 23102
rect 38892 22594 38948 22596
rect 38892 22542 38894 22594
rect 38894 22542 38946 22594
rect 38946 22542 38948 22594
rect 38892 22540 38948 22542
rect 37996 19068 38052 19124
rect 38108 21868 38164 21924
rect 38220 21474 38276 21476
rect 38220 21422 38222 21474
rect 38222 21422 38274 21474
rect 38274 21422 38276 21474
rect 38220 21420 38276 21422
rect 38332 20802 38388 20804
rect 38332 20750 38334 20802
rect 38334 20750 38386 20802
rect 38386 20750 38388 20802
rect 38332 20748 38388 20750
rect 38220 19964 38276 20020
rect 38668 20802 38724 20804
rect 38668 20750 38670 20802
rect 38670 20750 38722 20802
rect 38722 20750 38724 20802
rect 38668 20748 38724 20750
rect 38444 18956 38500 19012
rect 38556 19068 38612 19124
rect 38444 17666 38500 17668
rect 38444 17614 38446 17666
rect 38446 17614 38498 17666
rect 38498 17614 38500 17666
rect 38444 17612 38500 17614
rect 37996 17164 38052 17220
rect 37884 16828 37940 16884
rect 37996 15820 38052 15876
rect 39228 25676 39284 25732
rect 39564 25452 39620 25508
rect 39788 25564 39844 25620
rect 40236 26572 40292 26628
rect 40348 25676 40404 25732
rect 41132 25788 41188 25844
rect 40908 25564 40964 25620
rect 40796 25506 40852 25508
rect 40796 25454 40798 25506
rect 40798 25454 40850 25506
rect 40850 25454 40852 25506
rect 40796 25452 40852 25454
rect 40684 25340 40740 25396
rect 40012 24722 40068 24724
rect 40012 24670 40014 24722
rect 40014 24670 40066 24722
rect 40066 24670 40068 24722
rect 40012 24668 40068 24670
rect 40236 23772 40292 23828
rect 39116 23436 39172 23492
rect 39676 23100 39732 23156
rect 39228 22764 39284 22820
rect 39228 22428 39284 22484
rect 39228 22258 39284 22260
rect 39228 22206 39230 22258
rect 39230 22206 39282 22258
rect 39282 22206 39284 22258
rect 39228 22204 39284 22206
rect 39452 21420 39508 21476
rect 39340 21196 39396 21252
rect 39228 20524 39284 20580
rect 39228 19068 39284 19124
rect 39004 18060 39060 18116
rect 39004 17666 39060 17668
rect 39004 17614 39006 17666
rect 39006 17614 39058 17666
rect 39058 17614 39060 17666
rect 39004 17612 39060 17614
rect 39900 21868 39956 21924
rect 39676 20802 39732 20804
rect 39676 20750 39678 20802
rect 39678 20750 39730 20802
rect 39730 20750 39732 20802
rect 39676 20748 39732 20750
rect 39564 20636 39620 20692
rect 39676 20300 39732 20356
rect 39676 20076 39732 20132
rect 40348 23714 40404 23716
rect 40348 23662 40350 23714
rect 40350 23662 40402 23714
rect 40402 23662 40404 23714
rect 40348 23660 40404 23662
rect 40236 22316 40292 22372
rect 40236 21868 40292 21924
rect 40124 21756 40180 21812
rect 41020 23660 41076 23716
rect 41916 30268 41972 30324
rect 41916 29314 41972 29316
rect 41916 29262 41918 29314
rect 41918 29262 41970 29314
rect 41970 29262 41972 29314
rect 41916 29260 41972 29262
rect 41804 29202 41860 29204
rect 41804 29150 41806 29202
rect 41806 29150 41858 29202
rect 41858 29150 41860 29202
rect 41804 29148 41860 29150
rect 41692 28924 41748 28980
rect 41356 25452 41412 25508
rect 41916 25452 41972 25508
rect 42812 36428 42868 36484
rect 42924 35980 42980 36036
rect 43148 40012 43204 40068
rect 44044 41692 44100 41748
rect 44268 41746 44324 41748
rect 44268 41694 44270 41746
rect 44270 41694 44322 41746
rect 44322 41694 44324 41746
rect 44268 41692 44324 41694
rect 44492 42924 44548 42980
rect 44380 41580 44436 41636
rect 44268 41244 44324 41300
rect 43820 40460 43876 40516
rect 44828 47516 44884 47572
rect 45388 46060 45444 46116
rect 45276 45836 45332 45892
rect 44828 45666 44884 45668
rect 44828 45614 44830 45666
rect 44830 45614 44882 45666
rect 44882 45614 44884 45666
rect 44828 45612 44884 45614
rect 45724 47180 45780 47236
rect 46172 47234 46228 47236
rect 46172 47182 46174 47234
rect 46174 47182 46226 47234
rect 46226 47182 46228 47234
rect 46172 47180 46228 47182
rect 45836 46172 45892 46228
rect 45836 45948 45892 46004
rect 46844 47292 46900 47348
rect 45724 45164 45780 45220
rect 46732 45948 46788 46004
rect 46620 45164 46676 45220
rect 46060 44828 46116 44884
rect 45388 44716 45444 44772
rect 45948 44716 46004 44772
rect 44940 44268 44996 44324
rect 45836 44322 45892 44324
rect 45836 44270 45838 44322
rect 45838 44270 45890 44322
rect 45890 44270 45892 44322
rect 45836 44268 45892 44270
rect 45052 44210 45108 44212
rect 45052 44158 45054 44210
rect 45054 44158 45106 44210
rect 45106 44158 45108 44210
rect 45052 44156 45108 44158
rect 44828 44044 44884 44100
rect 44716 43708 44772 43764
rect 44828 43538 44884 43540
rect 44828 43486 44830 43538
rect 44830 43486 44882 43538
rect 44882 43486 44884 43538
rect 44828 43484 44884 43486
rect 46620 44604 46676 44660
rect 45052 43314 45108 43316
rect 45052 43262 45054 43314
rect 45054 43262 45106 43314
rect 45106 43262 45108 43314
rect 45052 43260 45108 43262
rect 44716 41970 44772 41972
rect 44716 41918 44718 41970
rect 44718 41918 44770 41970
rect 44770 41918 44772 41970
rect 44716 41916 44772 41918
rect 45388 42978 45444 42980
rect 45388 42926 45390 42978
rect 45390 42926 45442 42978
rect 45442 42926 45444 42978
rect 45388 42924 45444 42926
rect 46172 43372 46228 43428
rect 45836 43260 45892 43316
rect 46508 44322 46564 44324
rect 46508 44270 46510 44322
rect 46510 44270 46562 44322
rect 46562 44270 46564 44322
rect 46508 44268 46564 44270
rect 46508 43484 46564 43540
rect 45052 42642 45108 42644
rect 45052 42590 45054 42642
rect 45054 42590 45106 42642
rect 45106 42590 45108 42642
rect 45052 42588 45108 42590
rect 44940 42028 44996 42084
rect 45052 42364 45108 42420
rect 45276 41858 45332 41860
rect 45276 41806 45278 41858
rect 45278 41806 45330 41858
rect 45330 41806 45332 41858
rect 45276 41804 45332 41806
rect 43932 40124 43988 40180
rect 44716 40962 44772 40964
rect 44716 40910 44718 40962
rect 44718 40910 44770 40962
rect 44770 40910 44772 40962
rect 44716 40908 44772 40910
rect 43708 39676 43764 39732
rect 43484 39618 43540 39620
rect 43484 39566 43486 39618
rect 43486 39566 43538 39618
rect 43538 39566 43540 39618
rect 43484 39564 43540 39566
rect 43260 39506 43316 39508
rect 43260 39454 43262 39506
rect 43262 39454 43314 39506
rect 43314 39454 43316 39506
rect 43260 39452 43316 39454
rect 43372 39004 43428 39060
rect 43708 37996 43764 38052
rect 43484 37324 43540 37380
rect 45500 41580 45556 41636
rect 45388 41468 45444 41524
rect 45500 41132 45556 41188
rect 44156 40348 44212 40404
rect 44268 39228 44324 39284
rect 44940 40124 44996 40180
rect 45276 40572 45332 40628
rect 44828 39506 44884 39508
rect 44828 39454 44830 39506
rect 44830 39454 44882 39506
rect 44882 39454 44884 39506
rect 44828 39452 44884 39454
rect 44716 39394 44772 39396
rect 44716 39342 44718 39394
rect 44718 39342 44770 39394
rect 44770 39342 44772 39394
rect 44716 39340 44772 39342
rect 45388 39618 45444 39620
rect 45388 39566 45390 39618
rect 45390 39566 45442 39618
rect 45442 39566 45444 39618
rect 45388 39564 45444 39566
rect 45164 39228 45220 39284
rect 44156 38834 44212 38836
rect 44156 38782 44158 38834
rect 44158 38782 44210 38834
rect 44210 38782 44212 38834
rect 44156 38780 44212 38782
rect 44156 38162 44212 38164
rect 44156 38110 44158 38162
rect 44158 38110 44210 38162
rect 44210 38110 44212 38162
rect 44156 38108 44212 38110
rect 44604 38556 44660 38612
rect 44380 37996 44436 38052
rect 44044 36988 44100 37044
rect 43596 36876 43652 36932
rect 43148 36258 43204 36260
rect 43148 36206 43150 36258
rect 43150 36206 43202 36258
rect 43202 36206 43204 36258
rect 43148 36204 43204 36206
rect 43820 35084 43876 35140
rect 43932 34972 43988 35028
rect 43036 34130 43092 34132
rect 43036 34078 43038 34130
rect 43038 34078 43090 34130
rect 43090 34078 43092 34130
rect 43036 34076 43092 34078
rect 42812 32508 42868 32564
rect 43708 34130 43764 34132
rect 43708 34078 43710 34130
rect 43710 34078 43762 34130
rect 43762 34078 43764 34130
rect 43708 34076 43764 34078
rect 43932 34354 43988 34356
rect 43932 34302 43934 34354
rect 43934 34302 43986 34354
rect 43986 34302 43988 34354
rect 43932 34300 43988 34302
rect 44044 34188 44100 34244
rect 44380 35196 44436 35252
rect 43708 33852 43764 33908
rect 43372 33516 43428 33572
rect 43148 31836 43204 31892
rect 43484 32508 43540 32564
rect 43036 31500 43092 31556
rect 42924 31388 42980 31444
rect 42700 30828 42756 30884
rect 42588 30156 42644 30212
rect 43260 30380 43316 30436
rect 42700 29820 42756 29876
rect 42812 29932 42868 29988
rect 42924 29426 42980 29428
rect 42924 29374 42926 29426
rect 42926 29374 42978 29426
rect 42978 29374 42980 29426
rect 42924 29372 42980 29374
rect 42812 29260 42868 29316
rect 42140 28924 42196 28980
rect 42588 28476 42644 28532
rect 43820 31612 43876 31668
rect 43484 30940 43540 30996
rect 43372 30044 43428 30100
rect 44044 33740 44100 33796
rect 43932 30940 43988 30996
rect 43596 29820 43652 29876
rect 43148 28866 43204 28868
rect 43148 28814 43150 28866
rect 43150 28814 43202 28866
rect 43202 28814 43204 28866
rect 43148 28812 43204 28814
rect 43148 28530 43204 28532
rect 43148 28478 43150 28530
rect 43150 28478 43202 28530
rect 43202 28478 43204 28530
rect 43148 28476 43204 28478
rect 42028 25340 42084 25396
rect 42140 26460 42196 26516
rect 41468 25228 41524 25284
rect 41916 25116 41972 25172
rect 41580 24834 41636 24836
rect 41580 24782 41582 24834
rect 41582 24782 41634 24834
rect 41634 24782 41636 24834
rect 41580 24780 41636 24782
rect 41468 24556 41524 24612
rect 41804 24556 41860 24612
rect 42028 23996 42084 24052
rect 42028 23548 42084 23604
rect 40908 22540 40964 22596
rect 40684 22204 40740 22260
rect 40908 21532 40964 21588
rect 41356 21756 41412 21812
rect 40124 21196 40180 21252
rect 40460 20690 40516 20692
rect 40460 20638 40462 20690
rect 40462 20638 40514 20690
rect 40514 20638 40516 20690
rect 40460 20636 40516 20638
rect 40348 19628 40404 19684
rect 40236 18450 40292 18452
rect 40236 18398 40238 18450
rect 40238 18398 40290 18450
rect 40290 18398 40292 18450
rect 40236 18396 40292 18398
rect 40460 18284 40516 18340
rect 39788 17612 39844 17668
rect 39900 17836 39956 17892
rect 38892 17500 38948 17556
rect 38892 16940 38948 16996
rect 38668 16044 38724 16100
rect 38780 16604 38836 16660
rect 37660 15036 37716 15092
rect 37548 14530 37604 14532
rect 37548 14478 37550 14530
rect 37550 14478 37602 14530
rect 37602 14478 37604 14530
rect 37548 14476 37604 14478
rect 37324 13356 37380 13412
rect 37324 13020 37380 13076
rect 37100 12178 37156 12180
rect 37100 12126 37102 12178
rect 37102 12126 37154 12178
rect 37154 12126 37156 12178
rect 37100 12124 37156 12126
rect 37548 13132 37604 13188
rect 38108 14642 38164 14644
rect 38108 14590 38110 14642
rect 38110 14590 38162 14642
rect 38162 14590 38164 14642
rect 38108 14588 38164 14590
rect 37324 11788 37380 11844
rect 35532 11004 35588 11060
rect 35756 11228 35812 11284
rect 34076 10722 34132 10724
rect 34076 10670 34078 10722
rect 34078 10670 34130 10722
rect 34130 10670 34132 10722
rect 34076 10668 34132 10670
rect 33516 9884 33572 9940
rect 33516 9714 33572 9716
rect 33516 9662 33518 9714
rect 33518 9662 33570 9714
rect 33570 9662 33572 9714
rect 33516 9660 33572 9662
rect 34972 10722 35028 10724
rect 34972 10670 34974 10722
rect 34974 10670 35026 10722
rect 35026 10670 35028 10722
rect 34972 10668 35028 10670
rect 34412 10610 34468 10612
rect 34412 10558 34414 10610
rect 34414 10558 34466 10610
rect 34466 10558 34468 10610
rect 34412 10556 34468 10558
rect 34188 10108 34244 10164
rect 34524 9884 34580 9940
rect 33852 9154 33908 9156
rect 33852 9102 33854 9154
rect 33854 9102 33906 9154
rect 33906 9102 33908 9154
rect 33852 9100 33908 9102
rect 31612 8428 31668 8484
rect 30604 7474 30660 7476
rect 30604 7422 30606 7474
rect 30606 7422 30658 7474
rect 30658 7422 30660 7474
rect 30604 7420 30660 7422
rect 30716 8316 30772 8372
rect 32396 8818 32452 8820
rect 32396 8766 32398 8818
rect 32398 8766 32450 8818
rect 32450 8766 32452 8818
rect 32396 8764 32452 8766
rect 29596 5010 29652 5012
rect 29596 4958 29598 5010
rect 29598 4958 29650 5010
rect 29650 4958 29652 5010
rect 29596 4956 29652 4958
rect 30380 6524 30436 6580
rect 30492 6466 30548 6468
rect 30492 6414 30494 6466
rect 30494 6414 30546 6466
rect 30546 6414 30548 6466
rect 30492 6412 30548 6414
rect 31612 7644 31668 7700
rect 31052 7474 31108 7476
rect 31052 7422 31054 7474
rect 31054 7422 31106 7474
rect 31106 7422 31108 7474
rect 31052 7420 31108 7422
rect 30828 7196 30884 7252
rect 30828 6914 30884 6916
rect 30828 6862 30830 6914
rect 30830 6862 30882 6914
rect 30882 6862 30884 6914
rect 30828 6860 30884 6862
rect 30940 6748 30996 6804
rect 31276 5852 31332 5908
rect 31388 6188 31444 6244
rect 30268 4956 30324 5012
rect 28140 4898 28196 4900
rect 28140 4846 28142 4898
rect 28142 4846 28194 4898
rect 28194 4846 28196 4898
rect 28140 4844 28196 4846
rect 29708 4898 29764 4900
rect 29708 4846 29710 4898
rect 29710 4846 29762 4898
rect 29762 4846 29764 4898
rect 29708 4844 29764 4846
rect 29820 4732 29876 4788
rect 28028 4396 28084 4452
rect 31276 4956 31332 5012
rect 30716 4844 30772 4900
rect 31276 4732 31332 4788
rect 30268 4284 30324 4340
rect 28252 4226 28308 4228
rect 28252 4174 28254 4226
rect 28254 4174 28306 4226
rect 28306 4174 28308 4226
rect 28252 4172 28308 4174
rect 31052 4338 31108 4340
rect 31052 4286 31054 4338
rect 31054 4286 31106 4338
rect 31106 4286 31108 4338
rect 31052 4284 31108 4286
rect 31164 4226 31220 4228
rect 31164 4174 31166 4226
rect 31166 4174 31218 4226
rect 31218 4174 31220 4226
rect 31164 4172 31220 4174
rect 30492 3666 30548 3668
rect 30492 3614 30494 3666
rect 30494 3614 30546 3666
rect 30546 3614 30548 3666
rect 30492 3612 30548 3614
rect 31948 7420 32004 7476
rect 31836 6748 31892 6804
rect 32732 7532 32788 7588
rect 32284 6076 32340 6132
rect 32508 5852 32564 5908
rect 32396 5682 32452 5684
rect 32396 5630 32398 5682
rect 32398 5630 32450 5682
rect 32450 5630 32452 5682
rect 32396 5628 32452 5630
rect 31612 4956 31668 5012
rect 32284 4844 32340 4900
rect 31612 4450 31668 4452
rect 31612 4398 31614 4450
rect 31614 4398 31666 4450
rect 31666 4398 31668 4450
rect 31612 4396 31668 4398
rect 31612 3612 31668 3668
rect 29820 3388 29876 3444
rect 28364 3330 28420 3332
rect 28364 3278 28366 3330
rect 28366 3278 28418 3330
rect 28418 3278 28420 3330
rect 28364 3276 28420 3278
rect 32396 4620 32452 4676
rect 32060 3276 32116 3332
rect 32508 4450 32564 4452
rect 32508 4398 32510 4450
rect 32510 4398 32562 4450
rect 32562 4398 32564 4450
rect 32508 4396 32564 4398
rect 33740 8428 33796 8484
rect 34076 8428 34132 8484
rect 34524 9100 34580 9156
rect 35084 10556 35140 10612
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 33180 8146 33236 8148
rect 33180 8094 33182 8146
rect 33182 8094 33234 8146
rect 33234 8094 33236 8146
rect 33180 8092 33236 8094
rect 33292 7980 33348 8036
rect 33180 7586 33236 7588
rect 33180 7534 33182 7586
rect 33182 7534 33234 7586
rect 33234 7534 33236 7586
rect 33180 7532 33236 7534
rect 32956 7474 33012 7476
rect 32956 7422 32958 7474
rect 32958 7422 33010 7474
rect 33010 7422 33012 7474
rect 32956 7420 33012 7422
rect 33628 7586 33684 7588
rect 33628 7534 33630 7586
rect 33630 7534 33682 7586
rect 33682 7534 33684 7586
rect 33628 7532 33684 7534
rect 33964 8034 34020 8036
rect 33964 7982 33966 8034
rect 33966 7982 34018 8034
rect 34018 7982 34020 8034
rect 33964 7980 34020 7982
rect 33292 6748 33348 6804
rect 34188 7532 34244 7588
rect 36988 11004 37044 11060
rect 37100 11340 37156 11396
rect 36428 10892 36484 10948
rect 37324 11340 37380 11396
rect 36652 10722 36708 10724
rect 36652 10670 36654 10722
rect 36654 10670 36706 10722
rect 36706 10670 36708 10722
rect 36652 10668 36708 10670
rect 36316 10610 36372 10612
rect 36316 10558 36318 10610
rect 36318 10558 36370 10610
rect 36370 10558 36372 10610
rect 36316 10556 36372 10558
rect 35644 9938 35700 9940
rect 35644 9886 35646 9938
rect 35646 9886 35698 9938
rect 35698 9886 35700 9938
rect 35644 9884 35700 9886
rect 36428 9826 36484 9828
rect 36428 9774 36430 9826
rect 36430 9774 36482 9826
rect 36482 9774 36484 9826
rect 36428 9772 36484 9774
rect 37548 11394 37604 11396
rect 37548 11342 37550 11394
rect 37550 11342 37602 11394
rect 37602 11342 37604 11394
rect 37548 11340 37604 11342
rect 37548 10892 37604 10948
rect 37212 10108 37268 10164
rect 37100 9884 37156 9940
rect 38220 12738 38276 12740
rect 38220 12686 38222 12738
rect 38222 12686 38274 12738
rect 38274 12686 38276 12738
rect 38220 12684 38276 12686
rect 38444 15820 38500 15876
rect 38668 15874 38724 15876
rect 38668 15822 38670 15874
rect 38670 15822 38722 15874
rect 38722 15822 38724 15874
rect 38668 15820 38724 15822
rect 38556 15596 38612 15652
rect 39116 16492 39172 16548
rect 39452 16828 39508 16884
rect 38892 15538 38948 15540
rect 38892 15486 38894 15538
rect 38894 15486 38946 15538
rect 38946 15486 38948 15538
rect 38892 15484 38948 15486
rect 39340 15484 39396 15540
rect 39228 15426 39284 15428
rect 39228 15374 39230 15426
rect 39230 15374 39282 15426
rect 39282 15374 39284 15426
rect 39228 15372 39284 15374
rect 38780 15260 38836 15316
rect 39564 15820 39620 15876
rect 39676 15708 39732 15764
rect 40684 20524 40740 20580
rect 41020 20300 41076 20356
rect 40908 20188 40964 20244
rect 41356 20524 41412 20580
rect 41692 23436 41748 23492
rect 41804 23378 41860 23380
rect 41804 23326 41806 23378
rect 41806 23326 41858 23378
rect 41858 23326 41860 23378
rect 41804 23324 41860 23326
rect 42252 25116 42308 25172
rect 42140 22370 42196 22372
rect 42140 22318 42142 22370
rect 42142 22318 42194 22370
rect 42194 22318 42196 22370
rect 42140 22316 42196 22318
rect 42028 21532 42084 21588
rect 41468 21308 41524 21364
rect 41020 19740 41076 19796
rect 41356 19740 41412 19796
rect 41244 19404 41300 19460
rect 41132 17836 41188 17892
rect 40572 17500 40628 17556
rect 40348 16882 40404 16884
rect 40348 16830 40350 16882
rect 40350 16830 40402 16882
rect 40402 16830 40404 16882
rect 40348 16828 40404 16830
rect 38556 14924 38612 14980
rect 39340 15148 39396 15204
rect 38556 14530 38612 14532
rect 38556 14478 38558 14530
rect 38558 14478 38610 14530
rect 38610 14478 38612 14530
rect 38556 14476 38612 14478
rect 39228 15090 39284 15092
rect 39228 15038 39230 15090
rect 39230 15038 39282 15090
rect 39282 15038 39284 15090
rect 39228 15036 39284 15038
rect 39004 14812 39060 14868
rect 39004 14530 39060 14532
rect 39004 14478 39006 14530
rect 39006 14478 39058 14530
rect 39058 14478 39060 14530
rect 39004 14476 39060 14478
rect 38892 14418 38948 14420
rect 38892 14366 38894 14418
rect 38894 14366 38946 14418
rect 38946 14366 38948 14418
rect 38892 14364 38948 14366
rect 39788 15260 39844 15316
rect 39900 15426 39956 15428
rect 39900 15374 39902 15426
rect 39902 15374 39954 15426
rect 39954 15374 39956 15426
rect 39900 15372 39956 15374
rect 39564 14364 39620 14420
rect 40348 15820 40404 15876
rect 39788 14306 39844 14308
rect 39788 14254 39790 14306
rect 39790 14254 39842 14306
rect 39842 14254 39844 14306
rect 39788 14252 39844 14254
rect 40012 14306 40068 14308
rect 40012 14254 40014 14306
rect 40014 14254 40066 14306
rect 40066 14254 40068 14306
rect 40012 14252 40068 14254
rect 38668 12962 38724 12964
rect 38668 12910 38670 12962
rect 38670 12910 38722 12962
rect 38722 12910 38724 12962
rect 38668 12908 38724 12910
rect 39116 13244 39172 13300
rect 39004 12796 39060 12852
rect 39676 13858 39732 13860
rect 39676 13806 39678 13858
rect 39678 13806 39730 13858
rect 39730 13806 39732 13858
rect 39676 13804 39732 13806
rect 40236 14364 40292 14420
rect 40348 14140 40404 14196
rect 40460 14252 40516 14308
rect 40348 13916 40404 13972
rect 40236 13746 40292 13748
rect 40236 13694 40238 13746
rect 40238 13694 40290 13746
rect 40290 13694 40292 13746
rect 40236 13692 40292 13694
rect 40012 12684 40068 12740
rect 38332 11340 38388 11396
rect 39116 12348 39172 12404
rect 37884 9772 37940 9828
rect 38108 10892 38164 10948
rect 38220 9996 38276 10052
rect 38332 10108 38388 10164
rect 39564 12178 39620 12180
rect 39564 12126 39566 12178
rect 39566 12126 39618 12178
rect 39618 12126 39620 12178
rect 39564 12124 39620 12126
rect 39116 12012 39172 12068
rect 38668 9884 38724 9940
rect 38892 11900 38948 11956
rect 39004 9714 39060 9716
rect 39004 9662 39006 9714
rect 39006 9662 39058 9714
rect 39058 9662 39060 9714
rect 39004 9660 39060 9662
rect 39340 9996 39396 10052
rect 38444 8876 38500 8932
rect 34524 7980 34580 8036
rect 34748 7756 34804 7812
rect 35980 8316 36036 8372
rect 35308 8204 35364 8260
rect 35084 8146 35140 8148
rect 35084 8094 35086 8146
rect 35086 8094 35138 8146
rect 35138 8094 35140 8146
rect 35084 8092 35140 8094
rect 34860 7420 34916 7476
rect 34300 7250 34356 7252
rect 34300 7198 34302 7250
rect 34302 7198 34354 7250
rect 34354 7198 34356 7250
rect 34300 7196 34356 7198
rect 34524 6690 34580 6692
rect 34524 6638 34526 6690
rect 34526 6638 34578 6690
rect 34578 6638 34580 6690
rect 34524 6636 34580 6638
rect 32956 5122 33012 5124
rect 32956 5070 32958 5122
rect 32958 5070 33010 5122
rect 33010 5070 33012 5122
rect 32956 5068 33012 5070
rect 33852 4844 33908 4900
rect 33740 4620 33796 4676
rect 34300 6076 34356 6132
rect 34076 5628 34132 5684
rect 34188 5122 34244 5124
rect 34188 5070 34190 5122
rect 34190 5070 34242 5122
rect 34242 5070 34244 5122
rect 34188 5068 34244 5070
rect 34748 5122 34804 5124
rect 34748 5070 34750 5122
rect 34750 5070 34802 5122
rect 34802 5070 34804 5122
rect 34748 5068 34804 5070
rect 35868 8258 35924 8260
rect 35868 8206 35870 8258
rect 35870 8206 35922 8258
rect 35922 8206 35924 8258
rect 35868 8204 35924 8206
rect 37100 8258 37156 8260
rect 37100 8206 37102 8258
rect 37102 8206 37154 8258
rect 37154 8206 37156 8258
rect 37100 8204 37156 8206
rect 36316 8146 36372 8148
rect 36316 8094 36318 8146
rect 36318 8094 36370 8146
rect 36370 8094 36372 8146
rect 36316 8092 36372 8094
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35084 6860 35140 6916
rect 35756 6860 35812 6916
rect 35980 8034 36036 8036
rect 35980 7982 35982 8034
rect 35982 7982 36034 8034
rect 36034 7982 36036 8034
rect 35980 7980 36036 7982
rect 35644 6636 35700 6692
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35420 5122 35476 5124
rect 35420 5070 35422 5122
rect 35422 5070 35474 5122
rect 35474 5070 35476 5122
rect 35420 5068 35476 5070
rect 36092 6860 36148 6916
rect 36204 7644 36260 7700
rect 37548 7420 37604 7476
rect 37772 8092 37828 8148
rect 36204 6748 36260 6804
rect 36876 7196 36932 7252
rect 36092 6690 36148 6692
rect 36092 6638 36094 6690
rect 36094 6638 36146 6690
rect 36146 6638 36148 6690
rect 36092 6636 36148 6638
rect 35980 6524 36036 6580
rect 36428 6578 36484 6580
rect 36428 6526 36430 6578
rect 36430 6526 36482 6578
rect 36482 6526 36484 6578
rect 36428 6524 36484 6526
rect 36316 6188 36372 6244
rect 36092 5010 36148 5012
rect 36092 4958 36094 5010
rect 36094 4958 36146 5010
rect 36146 4958 36148 5010
rect 36092 4956 36148 4958
rect 34412 4620 34468 4676
rect 33740 4338 33796 4340
rect 33740 4286 33742 4338
rect 33742 4286 33794 4338
rect 33794 4286 33796 4338
rect 33740 4284 33796 4286
rect 35980 4620 36036 4676
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35196 3724 35252 3780
rect 33068 3388 33124 3444
rect 33404 3612 33460 3668
rect 32172 2828 32228 2884
rect 35084 3500 35140 3556
rect 36988 6690 37044 6692
rect 36988 6638 36990 6690
rect 36990 6638 37042 6690
rect 37042 6638 37044 6690
rect 36988 6636 37044 6638
rect 36876 6188 36932 6244
rect 36428 5628 36484 5684
rect 37212 4284 37268 4340
rect 36988 4060 37044 4116
rect 37548 6748 37604 6804
rect 37884 8034 37940 8036
rect 37884 7982 37886 8034
rect 37886 7982 37938 8034
rect 37938 7982 37940 8034
rect 37884 7980 37940 7982
rect 37884 7532 37940 7588
rect 37772 7420 37828 7476
rect 37884 4396 37940 4452
rect 38220 6748 38276 6804
rect 38556 7308 38612 7364
rect 38108 6076 38164 6132
rect 38332 6412 38388 6468
rect 38332 5906 38388 5908
rect 38332 5854 38334 5906
rect 38334 5854 38386 5906
rect 38386 5854 38388 5906
rect 38332 5852 38388 5854
rect 38892 8876 38948 8932
rect 39564 11788 39620 11844
rect 39788 11788 39844 11844
rect 40348 10332 40404 10388
rect 39788 9660 39844 9716
rect 39228 7980 39284 8036
rect 38668 6076 38724 6132
rect 38780 6690 38836 6692
rect 38780 6638 38782 6690
rect 38782 6638 38834 6690
rect 38834 6638 38836 6690
rect 38780 6636 38836 6638
rect 38780 5740 38836 5796
rect 39004 5906 39060 5908
rect 39004 5854 39006 5906
rect 39006 5854 39058 5906
rect 39058 5854 39060 5906
rect 39004 5852 39060 5854
rect 38220 5068 38276 5124
rect 38108 4396 38164 4452
rect 38780 4844 38836 4900
rect 38556 4114 38612 4116
rect 38556 4062 38558 4114
rect 38558 4062 38610 4114
rect 38610 4062 38612 4114
rect 38556 4060 38612 4062
rect 37436 3164 37492 3220
rect 39228 6018 39284 6020
rect 39228 5966 39230 6018
rect 39230 5966 39282 6018
rect 39282 5966 39284 6018
rect 39228 5964 39284 5966
rect 39564 7362 39620 7364
rect 39564 7310 39566 7362
rect 39566 7310 39618 7362
rect 39618 7310 39620 7362
rect 39564 7308 39620 7310
rect 39788 7474 39844 7476
rect 39788 7422 39790 7474
rect 39790 7422 39842 7474
rect 39842 7422 39844 7474
rect 39788 7420 39844 7422
rect 40460 9548 40516 9604
rect 41580 20130 41636 20132
rect 41580 20078 41582 20130
rect 41582 20078 41634 20130
rect 41634 20078 41636 20130
rect 41580 20076 41636 20078
rect 42028 20802 42084 20804
rect 42028 20750 42030 20802
rect 42030 20750 42082 20802
rect 42082 20750 42084 20802
rect 42028 20748 42084 20750
rect 41804 19404 41860 19460
rect 42028 19628 42084 19684
rect 41244 17388 41300 17444
rect 40908 16994 40964 16996
rect 40908 16942 40910 16994
rect 40910 16942 40962 16994
rect 40962 16942 40964 16994
rect 40908 16940 40964 16942
rect 41020 16716 41076 16772
rect 42700 26684 42756 26740
rect 43036 26850 43092 26852
rect 43036 26798 43038 26850
rect 43038 26798 43090 26850
rect 43090 26798 43092 26850
rect 43036 26796 43092 26798
rect 42924 26460 42980 26516
rect 43932 29932 43988 29988
rect 43708 28812 43764 28868
rect 45724 40796 45780 40852
rect 45948 41132 46004 41188
rect 46508 41916 46564 41972
rect 46396 41746 46452 41748
rect 46396 41694 46398 41746
rect 46398 41694 46450 41746
rect 46450 41694 46452 41746
rect 46396 41692 46452 41694
rect 45836 40348 45892 40404
rect 45724 39676 45780 39732
rect 46284 39394 46340 39396
rect 46284 39342 46286 39394
rect 46286 39342 46338 39394
rect 46338 39342 46340 39394
rect 46284 39340 46340 39342
rect 45948 38892 46004 38948
rect 46284 39004 46340 39060
rect 45724 38722 45780 38724
rect 45724 38670 45726 38722
rect 45726 38670 45778 38722
rect 45778 38670 45780 38722
rect 45724 38668 45780 38670
rect 45164 38556 45220 38612
rect 44828 37996 44884 38052
rect 45164 37378 45220 37380
rect 45164 37326 45166 37378
rect 45166 37326 45218 37378
rect 45218 37326 45220 37378
rect 45164 37324 45220 37326
rect 45500 37324 45556 37380
rect 45388 36876 45444 36932
rect 45276 36482 45332 36484
rect 45276 36430 45278 36482
rect 45278 36430 45330 36482
rect 45330 36430 45332 36482
rect 45276 36428 45332 36430
rect 47180 45948 47236 46004
rect 47180 44604 47236 44660
rect 47292 44492 47348 44548
rect 46956 43260 47012 43316
rect 47180 43426 47236 43428
rect 47180 43374 47182 43426
rect 47182 43374 47234 43426
rect 47234 43374 47236 43426
rect 47180 43372 47236 43374
rect 49084 47292 49140 47348
rect 48748 46956 48804 47012
rect 47740 46396 47796 46452
rect 47516 44268 47572 44324
rect 48412 45276 48468 45332
rect 49084 45890 49140 45892
rect 49084 45838 49086 45890
rect 49086 45838 49138 45890
rect 49138 45838 49140 45890
rect 49084 45836 49140 45838
rect 48636 43596 48692 43652
rect 47180 41970 47236 41972
rect 47180 41918 47182 41970
rect 47182 41918 47234 41970
rect 47234 41918 47236 41970
rect 47180 41916 47236 41918
rect 47964 43372 48020 43428
rect 47516 40796 47572 40852
rect 46844 40460 46900 40516
rect 47628 40348 47684 40404
rect 47292 40236 47348 40292
rect 46620 39116 46676 39172
rect 46732 40124 46788 40180
rect 46620 38892 46676 38948
rect 45612 36428 45668 36484
rect 45948 37212 46004 37268
rect 45164 36204 45220 36260
rect 45052 35084 45108 35140
rect 44268 34802 44324 34804
rect 44268 34750 44270 34802
rect 44270 34750 44322 34802
rect 44322 34750 44324 34802
rect 44268 34748 44324 34750
rect 44380 34354 44436 34356
rect 44380 34302 44382 34354
rect 44382 34302 44434 34354
rect 44434 34302 44436 34354
rect 44380 34300 44436 34302
rect 44268 32284 44324 32340
rect 44380 32396 44436 32452
rect 44268 31778 44324 31780
rect 44268 31726 44270 31778
rect 44270 31726 44322 31778
rect 44322 31726 44324 31778
rect 44268 31724 44324 31726
rect 44940 34748 44996 34804
rect 44716 34130 44772 34132
rect 44716 34078 44718 34130
rect 44718 34078 44770 34130
rect 44770 34078 44772 34130
rect 44716 34076 44772 34078
rect 44716 32562 44772 32564
rect 44716 32510 44718 32562
rect 44718 32510 44770 32562
rect 44770 32510 44772 32562
rect 44716 32508 44772 32510
rect 44604 31164 44660 31220
rect 45164 34076 45220 34132
rect 45276 34860 45332 34916
rect 45052 33740 45108 33796
rect 45164 33852 45220 33908
rect 45724 35868 45780 35924
rect 45836 35698 45892 35700
rect 45836 35646 45838 35698
rect 45838 35646 45890 35698
rect 45890 35646 45892 35698
rect 45836 35644 45892 35646
rect 45612 33964 45668 34020
rect 45276 33628 45332 33684
rect 45500 33740 45556 33796
rect 44940 32956 44996 33012
rect 44940 32786 44996 32788
rect 44940 32734 44942 32786
rect 44942 32734 44994 32786
rect 44994 32734 44996 32786
rect 44940 32732 44996 32734
rect 45164 33234 45220 33236
rect 45164 33182 45166 33234
rect 45166 33182 45218 33234
rect 45218 33182 45220 33234
rect 45164 33180 45220 33182
rect 45388 32508 45444 32564
rect 45836 33404 45892 33460
rect 47068 40012 47124 40068
rect 47068 39676 47124 39732
rect 47180 39618 47236 39620
rect 47180 39566 47182 39618
rect 47182 39566 47234 39618
rect 47234 39566 47236 39618
rect 47180 39564 47236 39566
rect 46956 39506 47012 39508
rect 46956 39454 46958 39506
rect 46958 39454 47010 39506
rect 47010 39454 47012 39506
rect 46956 39452 47012 39454
rect 47180 39340 47236 39396
rect 47068 38834 47124 38836
rect 47068 38782 47070 38834
rect 47070 38782 47122 38834
rect 47122 38782 47124 38834
rect 47068 38780 47124 38782
rect 46844 37324 46900 37380
rect 46620 36876 46676 36932
rect 47404 39452 47460 39508
rect 47404 39004 47460 39060
rect 47628 39506 47684 39508
rect 47628 39454 47630 39506
rect 47630 39454 47682 39506
rect 47682 39454 47684 39506
rect 47628 39452 47684 39454
rect 48076 43260 48132 43316
rect 48860 43426 48916 43428
rect 48860 43374 48862 43426
rect 48862 43374 48914 43426
rect 48914 43374 48916 43426
rect 48860 43372 48916 43374
rect 48636 42812 48692 42868
rect 48188 41858 48244 41860
rect 48188 41806 48190 41858
rect 48190 41806 48242 41858
rect 48242 41806 48244 41858
rect 48188 41804 48244 41806
rect 48860 40796 48916 40852
rect 48748 40348 48804 40404
rect 48748 40178 48804 40180
rect 48748 40126 48750 40178
rect 48750 40126 48802 40178
rect 48802 40126 48804 40178
rect 48748 40124 48804 40126
rect 47964 40012 48020 40068
rect 48188 39618 48244 39620
rect 48188 39566 48190 39618
rect 48190 39566 48242 39618
rect 48242 39566 48244 39618
rect 48188 39564 48244 39566
rect 47852 39340 47908 39396
rect 48076 38834 48132 38836
rect 48076 38782 48078 38834
rect 48078 38782 48130 38834
rect 48130 38782 48132 38834
rect 48076 38780 48132 38782
rect 48188 38722 48244 38724
rect 48188 38670 48190 38722
rect 48190 38670 48242 38722
rect 48242 38670 48244 38722
rect 48188 38668 48244 38670
rect 47964 36988 48020 37044
rect 47628 36204 47684 36260
rect 48972 40290 49028 40292
rect 48972 40238 48974 40290
rect 48974 40238 49026 40290
rect 49026 40238 49028 40290
rect 48972 40236 49028 40238
rect 49196 42866 49252 42868
rect 49196 42814 49198 42866
rect 49198 42814 49250 42866
rect 49250 42814 49252 42866
rect 49196 42812 49252 42814
rect 49196 41298 49252 41300
rect 49196 41246 49198 41298
rect 49198 41246 49250 41298
rect 49250 41246 49252 41298
rect 49196 41244 49252 41246
rect 48748 38946 48804 38948
rect 48748 38894 48750 38946
rect 48750 38894 48802 38946
rect 48802 38894 48804 38946
rect 48748 38892 48804 38894
rect 48748 37378 48804 37380
rect 48748 37326 48750 37378
rect 48750 37326 48802 37378
rect 48802 37326 48804 37378
rect 48748 37324 48804 37326
rect 48860 36988 48916 37044
rect 48412 36428 48468 36484
rect 47180 35196 47236 35252
rect 46956 34802 47012 34804
rect 46956 34750 46958 34802
rect 46958 34750 47010 34802
rect 47010 34750 47012 34802
rect 46956 34748 47012 34750
rect 46172 34018 46228 34020
rect 46172 33966 46174 34018
rect 46174 33966 46226 34018
rect 46226 33966 46228 34018
rect 46172 33964 46228 33966
rect 46508 33906 46564 33908
rect 46508 33854 46510 33906
rect 46510 33854 46562 33906
rect 46562 33854 46564 33906
rect 46508 33852 46564 33854
rect 45052 32284 45108 32340
rect 44940 31890 44996 31892
rect 44940 31838 44942 31890
rect 44942 31838 44994 31890
rect 44994 31838 44996 31890
rect 44940 31836 44996 31838
rect 44940 31052 44996 31108
rect 45724 32450 45780 32452
rect 45724 32398 45726 32450
rect 45726 32398 45778 32450
rect 45778 32398 45780 32450
rect 45724 32396 45780 32398
rect 45500 32172 45556 32228
rect 45724 31948 45780 32004
rect 44156 30156 44212 30212
rect 44044 28700 44100 28756
rect 44380 28588 44436 28644
rect 44716 29372 44772 29428
rect 44156 27746 44212 27748
rect 44156 27694 44158 27746
rect 44158 27694 44210 27746
rect 44210 27694 44212 27746
rect 44156 27692 44212 27694
rect 42476 26178 42532 26180
rect 42476 26126 42478 26178
rect 42478 26126 42530 26178
rect 42530 26126 42532 26178
rect 42476 26124 42532 26126
rect 42364 21532 42420 21588
rect 42588 24668 42644 24724
rect 42588 23042 42644 23044
rect 42588 22990 42590 23042
rect 42590 22990 42642 23042
rect 42642 22990 42644 23042
rect 42588 22988 42644 22990
rect 43484 26124 43540 26180
rect 43596 26684 43652 26740
rect 42924 25676 42980 25732
rect 42924 25228 42980 25284
rect 44044 26850 44100 26852
rect 44044 26798 44046 26850
rect 44046 26798 44098 26850
rect 44098 26798 44100 26850
rect 44044 26796 44100 26798
rect 43036 24332 43092 24388
rect 43148 23548 43204 23604
rect 42812 22988 42868 23044
rect 42588 22316 42644 22372
rect 42588 20748 42644 20804
rect 42364 20690 42420 20692
rect 42364 20638 42366 20690
rect 42366 20638 42418 20690
rect 42418 20638 42420 20690
rect 42364 20636 42420 20638
rect 42252 20188 42308 20244
rect 42476 19852 42532 19908
rect 42252 19740 42308 19796
rect 41916 18508 41972 18564
rect 42028 18450 42084 18452
rect 42028 18398 42030 18450
rect 42030 18398 42082 18450
rect 42082 18398 42084 18450
rect 42028 18396 42084 18398
rect 42812 20412 42868 20468
rect 43036 22764 43092 22820
rect 42700 19740 42756 19796
rect 43596 25394 43652 25396
rect 43596 25342 43598 25394
rect 43598 25342 43650 25394
rect 43650 25342 43652 25394
rect 43596 25340 43652 25342
rect 43820 25452 43876 25508
rect 44716 27858 44772 27860
rect 44716 27806 44718 27858
rect 44718 27806 44770 27858
rect 44770 27806 44772 27858
rect 44716 27804 44772 27806
rect 45052 30492 45108 30548
rect 45164 30268 45220 30324
rect 45276 30716 45332 30772
rect 45836 31724 45892 31780
rect 45612 31666 45668 31668
rect 45612 31614 45614 31666
rect 45614 31614 45666 31666
rect 45666 31614 45668 31666
rect 45612 31612 45668 31614
rect 45612 31218 45668 31220
rect 45612 31166 45614 31218
rect 45614 31166 45666 31218
rect 45666 31166 45668 31218
rect 45612 31164 45668 31166
rect 45500 29820 45556 29876
rect 45724 29986 45780 29988
rect 45724 29934 45726 29986
rect 45726 29934 45778 29986
rect 45778 29934 45780 29986
rect 45724 29932 45780 29934
rect 45612 29708 45668 29764
rect 46620 32562 46676 32564
rect 46620 32510 46622 32562
rect 46622 32510 46674 32562
rect 46674 32510 46676 32562
rect 46620 32508 46676 32510
rect 46284 31948 46340 32004
rect 46060 30994 46116 30996
rect 46060 30942 46062 30994
rect 46062 30942 46114 30994
rect 46114 30942 46116 30994
rect 46060 30940 46116 30942
rect 45948 29986 46004 29988
rect 45948 29934 45950 29986
rect 45950 29934 46002 29986
rect 46002 29934 46004 29986
rect 45948 29932 46004 29934
rect 46284 30882 46340 30884
rect 46284 30830 46286 30882
rect 46286 30830 46338 30882
rect 46338 30830 46340 30882
rect 46284 30828 46340 30830
rect 47068 33852 47124 33908
rect 47068 33458 47124 33460
rect 47068 33406 47070 33458
rect 47070 33406 47122 33458
rect 47122 33406 47124 33458
rect 47068 33404 47124 33406
rect 47404 34354 47460 34356
rect 47404 34302 47406 34354
rect 47406 34302 47458 34354
rect 47458 34302 47460 34354
rect 47404 34300 47460 34302
rect 46732 31836 46788 31892
rect 46508 31724 46564 31780
rect 46508 31500 46564 31556
rect 46620 31612 46676 31668
rect 46508 30492 46564 30548
rect 46396 30380 46452 30436
rect 46620 30268 46676 30324
rect 46396 30210 46452 30212
rect 46396 30158 46398 30210
rect 46398 30158 46450 30210
rect 46450 30158 46452 30210
rect 46396 30156 46452 30158
rect 46844 31388 46900 31444
rect 46844 30770 46900 30772
rect 46844 30718 46846 30770
rect 46846 30718 46898 30770
rect 46898 30718 46900 30770
rect 46844 30716 46900 30718
rect 45500 28700 45556 28756
rect 46060 28642 46116 28644
rect 46060 28590 46062 28642
rect 46062 28590 46114 28642
rect 46114 28590 46116 28642
rect 46060 28588 46116 28590
rect 45388 28476 45444 28532
rect 45052 27692 45108 27748
rect 44268 26236 44324 26292
rect 44268 25564 44324 25620
rect 43932 25282 43988 25284
rect 43932 25230 43934 25282
rect 43934 25230 43986 25282
rect 43986 25230 43988 25282
rect 43932 25228 43988 25230
rect 44828 25116 44884 25172
rect 43708 24892 43764 24948
rect 43372 24556 43428 24612
rect 43484 24668 43540 24724
rect 43484 23938 43540 23940
rect 43484 23886 43486 23938
rect 43486 23886 43538 23938
rect 43538 23886 43540 23938
rect 43484 23884 43540 23886
rect 43372 23436 43428 23492
rect 43372 22764 43428 22820
rect 43036 21532 43092 21588
rect 43148 20802 43204 20804
rect 43148 20750 43150 20802
rect 43150 20750 43202 20802
rect 43202 20750 43204 20802
rect 43148 20748 43204 20750
rect 43932 24556 43988 24612
rect 43596 22988 43652 23044
rect 45836 27804 45892 27860
rect 46732 29986 46788 29988
rect 46732 29934 46734 29986
rect 46734 29934 46786 29986
rect 46786 29934 46788 29986
rect 46732 29932 46788 29934
rect 46844 29708 46900 29764
rect 45276 26460 45332 26516
rect 46060 26514 46116 26516
rect 46060 26462 46062 26514
rect 46062 26462 46114 26514
rect 46114 26462 46116 26514
rect 46060 26460 46116 26462
rect 45724 26290 45780 26292
rect 45724 26238 45726 26290
rect 45726 26238 45778 26290
rect 45778 26238 45780 26290
rect 45724 26236 45780 26238
rect 44380 24610 44436 24612
rect 44380 24558 44382 24610
rect 44382 24558 44434 24610
rect 44434 24558 44436 24610
rect 44380 24556 44436 24558
rect 44828 23938 44884 23940
rect 44828 23886 44830 23938
rect 44830 23886 44882 23938
rect 44882 23886 44884 23938
rect 44828 23884 44884 23886
rect 44156 23660 44212 23716
rect 44940 23548 44996 23604
rect 44604 22652 44660 22708
rect 44156 22540 44212 22596
rect 42924 19628 42980 19684
rect 43036 19964 43092 20020
rect 42476 18956 42532 19012
rect 43036 19292 43092 19348
rect 42924 19010 42980 19012
rect 42924 18958 42926 19010
rect 42926 18958 42978 19010
rect 42978 18958 42980 19010
rect 42924 18956 42980 18958
rect 42364 18396 42420 18452
rect 42812 18396 42868 18452
rect 42140 18338 42196 18340
rect 42140 18286 42142 18338
rect 42142 18286 42194 18338
rect 42194 18286 42196 18338
rect 42140 18284 42196 18286
rect 41468 16882 41524 16884
rect 41468 16830 41470 16882
rect 41470 16830 41522 16882
rect 41522 16830 41524 16882
rect 41468 16828 41524 16830
rect 42588 18172 42644 18228
rect 41916 16604 41972 16660
rect 40572 15260 40628 15316
rect 40796 14924 40852 14980
rect 41132 15426 41188 15428
rect 41132 15374 41134 15426
rect 41134 15374 41186 15426
rect 41186 15374 41188 15426
rect 41132 15372 41188 15374
rect 41020 13970 41076 13972
rect 41020 13918 41022 13970
rect 41022 13918 41074 13970
rect 41074 13918 41076 13970
rect 41020 13916 41076 13918
rect 41692 15036 41748 15092
rect 41356 14642 41412 14644
rect 41356 14590 41358 14642
rect 41358 14590 41410 14642
rect 41410 14590 41412 14642
rect 41356 14588 41412 14590
rect 41244 13970 41300 13972
rect 41244 13918 41246 13970
rect 41246 13918 41298 13970
rect 41298 13918 41300 13970
rect 41244 13916 41300 13918
rect 42028 15092 42084 15148
rect 41468 13804 41524 13860
rect 41356 13746 41412 13748
rect 41356 13694 41358 13746
rect 41358 13694 41410 13746
rect 41410 13694 41412 13746
rect 41356 13692 41412 13694
rect 42252 14588 42308 14644
rect 42028 13804 42084 13860
rect 42140 13916 42196 13972
rect 41804 13468 41860 13524
rect 41580 13244 41636 13300
rect 41244 12572 41300 12628
rect 41244 12178 41300 12180
rect 41244 12126 41246 12178
rect 41246 12126 41298 12178
rect 41298 12126 41300 12178
rect 41244 12124 41300 12126
rect 41468 12178 41524 12180
rect 41468 12126 41470 12178
rect 41470 12126 41522 12178
rect 41522 12126 41524 12178
rect 41468 12124 41524 12126
rect 41020 12066 41076 12068
rect 41020 12014 41022 12066
rect 41022 12014 41074 12066
rect 41074 12014 41076 12066
rect 41020 12012 41076 12014
rect 41692 11788 41748 11844
rect 41244 10722 41300 10724
rect 41244 10670 41246 10722
rect 41246 10670 41298 10722
rect 41298 10670 41300 10722
rect 41244 10668 41300 10670
rect 41468 10386 41524 10388
rect 41468 10334 41470 10386
rect 41470 10334 41522 10386
rect 41522 10334 41524 10386
rect 41468 10332 41524 10334
rect 41244 10220 41300 10276
rect 41132 9938 41188 9940
rect 41132 9886 41134 9938
rect 41134 9886 41186 9938
rect 41186 9886 41188 9938
rect 41132 9884 41188 9886
rect 43036 18508 43092 18564
rect 42924 15986 42980 15988
rect 42924 15934 42926 15986
rect 42926 15934 42978 15986
rect 42978 15934 42980 15986
rect 42924 15932 42980 15934
rect 42812 13970 42868 13972
rect 42812 13918 42814 13970
rect 42814 13918 42866 13970
rect 42866 13918 42868 13970
rect 42812 13916 42868 13918
rect 42588 13468 42644 13524
rect 42812 13468 42868 13524
rect 41916 12684 41972 12740
rect 42028 12796 42084 12852
rect 41916 10444 41972 10500
rect 41804 10108 41860 10164
rect 42700 13244 42756 13300
rect 42364 13020 42420 13076
rect 42476 12684 42532 12740
rect 42588 12348 42644 12404
rect 42700 12236 42756 12292
rect 42812 12348 42868 12404
rect 42924 12012 42980 12068
rect 42476 11900 42532 11956
rect 43372 20578 43428 20580
rect 43372 20526 43374 20578
rect 43374 20526 43426 20578
rect 43426 20526 43428 20578
rect 43372 20524 43428 20526
rect 43260 20412 43316 20468
rect 43596 19964 43652 20020
rect 43260 19852 43316 19908
rect 43596 19180 43652 19236
rect 43484 18508 43540 18564
rect 43372 17948 43428 18004
rect 44044 20690 44100 20692
rect 44044 20638 44046 20690
rect 44046 20638 44098 20690
rect 44098 20638 44100 20690
rect 44044 20636 44100 20638
rect 44044 19852 44100 19908
rect 44268 19516 44324 19572
rect 44268 19068 44324 19124
rect 43932 18844 43988 18900
rect 44156 18844 44212 18900
rect 44268 18396 44324 18452
rect 44156 17388 44212 17444
rect 45836 25228 45892 25284
rect 47068 29484 47124 29540
rect 47628 34914 47684 34916
rect 47628 34862 47630 34914
rect 47630 34862 47682 34914
rect 47682 34862 47684 34914
rect 47628 34860 47684 34862
rect 47740 34636 47796 34692
rect 47628 34018 47684 34020
rect 47628 33966 47630 34018
rect 47630 33966 47682 34018
rect 47682 33966 47684 34018
rect 47628 33964 47684 33966
rect 47628 32562 47684 32564
rect 47628 32510 47630 32562
rect 47630 32510 47682 32562
rect 47682 32510 47684 32562
rect 47628 32508 47684 32510
rect 48188 35026 48244 35028
rect 48188 34974 48190 35026
rect 48190 34974 48242 35026
rect 48242 34974 48244 35026
rect 48188 34972 48244 34974
rect 48188 34636 48244 34692
rect 48076 32844 48132 32900
rect 48076 32674 48132 32676
rect 48076 32622 48078 32674
rect 48078 32622 48130 32674
rect 48130 32622 48132 32674
rect 48076 32620 48132 32622
rect 47852 32396 47908 32452
rect 48076 32396 48132 32452
rect 47740 31836 47796 31892
rect 48748 35922 48804 35924
rect 48748 35870 48750 35922
rect 48750 35870 48802 35922
rect 48802 35870 48804 35922
rect 48748 35868 48804 35870
rect 49196 38668 49252 38724
rect 49084 37266 49140 37268
rect 49084 37214 49086 37266
rect 49086 37214 49138 37266
rect 49138 37214 49140 37266
rect 49084 37212 49140 37214
rect 49084 36988 49140 37044
rect 49196 36594 49252 36596
rect 49196 36542 49198 36594
rect 49198 36542 49250 36594
rect 49250 36542 49252 36594
rect 49196 36540 49252 36542
rect 49084 36092 49140 36148
rect 48412 34188 48468 34244
rect 48300 31836 48356 31892
rect 48412 32508 48468 32564
rect 47516 31724 47572 31780
rect 48524 32396 48580 32452
rect 47292 30940 47348 30996
rect 47628 30994 47684 30996
rect 47628 30942 47630 30994
rect 47630 30942 47682 30994
rect 47682 30942 47684 30994
rect 47628 30940 47684 30942
rect 47404 30434 47460 30436
rect 47404 30382 47406 30434
rect 47406 30382 47458 30434
rect 47458 30382 47460 30434
rect 47404 30380 47460 30382
rect 47516 30268 47572 30324
rect 47404 30210 47460 30212
rect 47404 30158 47406 30210
rect 47406 30158 47458 30210
rect 47458 30158 47460 30210
rect 47404 30156 47460 30158
rect 47740 30268 47796 30324
rect 47404 29932 47460 29988
rect 47740 28866 47796 28868
rect 47740 28814 47742 28866
rect 47742 28814 47794 28866
rect 47794 28814 47796 28866
rect 47740 28812 47796 28814
rect 47404 28588 47460 28644
rect 48076 30604 48132 30660
rect 47964 30380 48020 30436
rect 48748 34748 48804 34804
rect 48748 34300 48804 34356
rect 49420 41244 49476 41300
rect 49308 36092 49364 36148
rect 49420 40796 49476 40852
rect 48860 33964 48916 34020
rect 48748 32674 48804 32676
rect 48748 32622 48750 32674
rect 48750 32622 48802 32674
rect 48802 32622 48804 32674
rect 48748 32620 48804 32622
rect 48188 30210 48244 30212
rect 48188 30158 48190 30210
rect 48190 30158 48242 30210
rect 48242 30158 48244 30210
rect 48188 30156 48244 30158
rect 48076 28642 48132 28644
rect 48076 28590 48078 28642
rect 48078 28590 48130 28642
rect 48130 28590 48132 28642
rect 48076 28588 48132 28590
rect 48524 30604 48580 30660
rect 48636 30492 48692 30548
rect 46620 27692 46676 27748
rect 46508 27634 46564 27636
rect 46508 27582 46510 27634
rect 46510 27582 46562 27634
rect 46562 27582 46564 27634
rect 46508 27580 46564 27582
rect 46508 26514 46564 26516
rect 46508 26462 46510 26514
rect 46510 26462 46562 26514
rect 46562 26462 46564 26514
rect 46508 26460 46564 26462
rect 47068 26962 47124 26964
rect 47068 26910 47070 26962
rect 47070 26910 47122 26962
rect 47122 26910 47124 26962
rect 47068 26908 47124 26910
rect 46620 26402 46676 26404
rect 46620 26350 46622 26402
rect 46622 26350 46674 26402
rect 46674 26350 46676 26402
rect 46620 26348 46676 26350
rect 46844 26402 46900 26404
rect 46844 26350 46846 26402
rect 46846 26350 46898 26402
rect 46898 26350 46900 26402
rect 46844 26348 46900 26350
rect 46732 26178 46788 26180
rect 46732 26126 46734 26178
rect 46734 26126 46786 26178
rect 46786 26126 46788 26178
rect 46732 26124 46788 26126
rect 47068 26290 47124 26292
rect 47068 26238 47070 26290
rect 47070 26238 47122 26290
rect 47122 26238 47124 26290
rect 47068 26236 47124 26238
rect 46396 25228 46452 25284
rect 46284 24834 46340 24836
rect 46284 24782 46286 24834
rect 46286 24782 46338 24834
rect 46338 24782 46340 24834
rect 46284 24780 46340 24782
rect 45836 24668 45892 24724
rect 46172 24610 46228 24612
rect 46172 24558 46174 24610
rect 46174 24558 46226 24610
rect 46226 24558 46228 24610
rect 46172 24556 46228 24558
rect 45500 23660 45556 23716
rect 46060 23436 46116 23492
rect 45388 22540 45444 22596
rect 44940 22482 44996 22484
rect 44940 22430 44942 22482
rect 44942 22430 44994 22482
rect 44994 22430 44996 22482
rect 44940 22428 44996 22430
rect 46956 25676 47012 25732
rect 47180 24946 47236 24948
rect 47180 24894 47182 24946
rect 47182 24894 47234 24946
rect 47234 24894 47236 24946
rect 47180 24892 47236 24894
rect 47068 24444 47124 24500
rect 45948 22370 46004 22372
rect 45948 22318 45950 22370
rect 45950 22318 46002 22370
rect 46002 22318 46004 22370
rect 45948 22316 46004 22318
rect 45500 22146 45556 22148
rect 45500 22094 45502 22146
rect 45502 22094 45554 22146
rect 45554 22094 45556 22146
rect 45500 22092 45556 22094
rect 46844 21810 46900 21812
rect 46844 21758 46846 21810
rect 46846 21758 46898 21810
rect 46898 21758 46900 21810
rect 46844 21756 46900 21758
rect 47516 26908 47572 26964
rect 48076 27132 48132 27188
rect 47628 26572 47684 26628
rect 47516 26460 47572 26516
rect 47516 25340 47572 25396
rect 47852 26348 47908 26404
rect 47740 25116 47796 25172
rect 47628 24332 47684 24388
rect 48860 30434 48916 30436
rect 48860 30382 48862 30434
rect 48862 30382 48914 30434
rect 48914 30382 48916 30434
rect 48860 30380 48916 30382
rect 48748 30268 48804 30324
rect 48860 29538 48916 29540
rect 48860 29486 48862 29538
rect 48862 29486 48914 29538
rect 48914 29486 48916 29538
rect 48860 29484 48916 29486
rect 48412 27580 48468 27636
rect 48748 27634 48804 27636
rect 48748 27582 48750 27634
rect 48750 27582 48802 27634
rect 48802 27582 48804 27634
rect 48748 27580 48804 27582
rect 49084 32284 49140 32340
rect 49196 31890 49252 31892
rect 49196 31838 49198 31890
rect 49198 31838 49250 31890
rect 49250 31838 49252 31890
rect 49196 31836 49252 31838
rect 49308 30940 49364 30996
rect 49084 30044 49140 30100
rect 48972 27692 49028 27748
rect 49084 29484 49140 29540
rect 48860 27132 48916 27188
rect 49196 27580 49252 27636
rect 49196 27186 49252 27188
rect 49196 27134 49198 27186
rect 49198 27134 49250 27186
rect 49250 27134 49252 27186
rect 49196 27132 49252 27134
rect 49644 40012 49700 40068
rect 49532 39564 49588 39620
rect 49532 36540 49588 36596
rect 49532 30380 49588 30436
rect 48748 26572 48804 26628
rect 48188 26236 48244 26292
rect 48860 26178 48916 26180
rect 48860 26126 48862 26178
rect 48862 26126 48914 26178
rect 48914 26126 48916 26178
rect 48860 26124 48916 26126
rect 48748 25676 48804 25732
rect 48188 25564 48244 25620
rect 48188 25340 48244 25396
rect 47852 24668 47908 24724
rect 47852 23772 47908 23828
rect 48076 24722 48132 24724
rect 48076 24670 48078 24722
rect 48078 24670 48130 24722
rect 48130 24670 48132 24722
rect 48076 24668 48132 24670
rect 48748 24498 48804 24500
rect 48748 24446 48750 24498
rect 48750 24446 48802 24498
rect 48802 24446 48804 24498
rect 48748 24444 48804 24446
rect 48300 24332 48356 24388
rect 48524 23826 48580 23828
rect 48524 23774 48526 23826
rect 48526 23774 48578 23826
rect 48578 23774 48580 23826
rect 48524 23772 48580 23774
rect 49084 25618 49140 25620
rect 49084 25566 49086 25618
rect 49086 25566 49138 25618
rect 49138 25566 49140 25618
rect 49084 25564 49140 25566
rect 49196 24050 49252 24052
rect 49196 23998 49198 24050
rect 49198 23998 49250 24050
rect 49250 23998 49252 24050
rect 49196 23996 49252 23998
rect 48076 23324 48132 23380
rect 47292 22092 47348 22148
rect 47740 21810 47796 21812
rect 47740 21758 47742 21810
rect 47742 21758 47794 21810
rect 47794 21758 47796 21810
rect 47740 21756 47796 21758
rect 45724 20802 45780 20804
rect 45724 20750 45726 20802
rect 45726 20750 45778 20802
rect 45778 20750 45780 20802
rect 45724 20748 45780 20750
rect 44828 20524 44884 20580
rect 44940 20076 44996 20132
rect 45052 19964 45108 20020
rect 45164 20076 45220 20132
rect 45052 19740 45108 19796
rect 45724 20018 45780 20020
rect 45724 19966 45726 20018
rect 45726 19966 45778 20018
rect 45778 19966 45780 20018
rect 45724 19964 45780 19966
rect 45612 19906 45668 19908
rect 45612 19854 45614 19906
rect 45614 19854 45666 19906
rect 45666 19854 45668 19906
rect 45612 19852 45668 19854
rect 45500 19234 45556 19236
rect 45500 19182 45502 19234
rect 45502 19182 45554 19234
rect 45554 19182 45556 19234
rect 45500 19180 45556 19182
rect 44604 16604 44660 16660
rect 44716 17612 44772 17668
rect 45724 18284 45780 18340
rect 46284 20076 46340 20132
rect 46060 19852 46116 19908
rect 45948 18508 46004 18564
rect 44716 16882 44772 16884
rect 44716 16830 44718 16882
rect 44718 16830 44770 16882
rect 44770 16830 44772 16882
rect 44716 16828 44772 16830
rect 44492 16492 44548 16548
rect 43484 13580 43540 13636
rect 43820 15932 43876 15988
rect 43596 12796 43652 12852
rect 43708 13356 43764 13412
rect 43372 12348 43428 12404
rect 43260 12236 43316 12292
rect 43484 12178 43540 12180
rect 43484 12126 43486 12178
rect 43486 12126 43538 12178
rect 43538 12126 43540 12178
rect 43484 12124 43540 12126
rect 43148 11676 43204 11732
rect 43484 11788 43540 11844
rect 42028 9996 42084 10052
rect 42924 10668 42980 10724
rect 41692 9884 41748 9940
rect 41356 9324 41412 9380
rect 42028 9772 42084 9828
rect 42140 9324 42196 9380
rect 41468 8988 41524 9044
rect 40908 8316 40964 8372
rect 40012 7756 40068 7812
rect 40124 7644 40180 7700
rect 39788 6860 39844 6916
rect 39452 6524 39508 6580
rect 41356 8428 41412 8484
rect 41132 7362 41188 7364
rect 41132 7310 41134 7362
rect 41134 7310 41186 7362
rect 41186 7310 41188 7362
rect 41132 7308 41188 7310
rect 41244 7196 41300 7252
rect 40348 5740 40404 5796
rect 41020 5740 41076 5796
rect 41916 7644 41972 7700
rect 41580 7474 41636 7476
rect 41580 7422 41582 7474
rect 41582 7422 41634 7474
rect 41634 7422 41636 7474
rect 41580 7420 41636 7422
rect 42140 8146 42196 8148
rect 42140 8094 42142 8146
rect 42142 8094 42194 8146
rect 42194 8094 42196 8146
rect 42140 8092 42196 8094
rect 42588 10498 42644 10500
rect 42588 10446 42590 10498
rect 42590 10446 42642 10498
rect 42642 10446 42644 10498
rect 42588 10444 42644 10446
rect 42588 9996 42644 10052
rect 42476 9436 42532 9492
rect 42476 9212 42532 9268
rect 42588 8930 42644 8932
rect 42588 8878 42590 8930
rect 42590 8878 42642 8930
rect 42642 8878 42644 8930
rect 42588 8876 42644 8878
rect 42812 7980 42868 8036
rect 42588 7756 42644 7812
rect 42476 6802 42532 6804
rect 42476 6750 42478 6802
rect 42478 6750 42530 6802
rect 42530 6750 42532 6802
rect 42476 6748 42532 6750
rect 42140 6578 42196 6580
rect 42140 6526 42142 6578
rect 42142 6526 42194 6578
rect 42194 6526 42196 6578
rect 42140 6524 42196 6526
rect 42364 6466 42420 6468
rect 42364 6414 42366 6466
rect 42366 6414 42418 6466
rect 42418 6414 42420 6466
rect 42364 6412 42420 6414
rect 41356 5740 41412 5796
rect 39788 4844 39844 4900
rect 39340 3724 39396 3780
rect 40572 4508 40628 4564
rect 39788 3554 39844 3556
rect 39788 3502 39790 3554
rect 39790 3502 39842 3554
rect 39842 3502 39844 3554
rect 39788 3500 39844 3502
rect 41020 5010 41076 5012
rect 41020 4958 41022 5010
rect 41022 4958 41074 5010
rect 41074 4958 41076 5010
rect 41020 4956 41076 4958
rect 40796 3666 40852 3668
rect 40796 3614 40798 3666
rect 40798 3614 40850 3666
rect 40850 3614 40852 3666
rect 40796 3612 40852 3614
rect 43036 7196 43092 7252
rect 44940 16492 44996 16548
rect 44828 14924 44884 14980
rect 44268 13580 44324 13636
rect 44492 13804 44548 13860
rect 44156 13468 44212 13524
rect 44044 12796 44100 12852
rect 43708 11900 43764 11956
rect 43596 11564 43652 11620
rect 43484 11228 43540 11284
rect 43820 11282 43876 11284
rect 43820 11230 43822 11282
rect 43822 11230 43874 11282
rect 43874 11230 43876 11282
rect 43820 11228 43876 11230
rect 44268 11954 44324 11956
rect 44268 11902 44270 11954
rect 44270 11902 44322 11954
rect 44322 11902 44324 11954
rect 44268 11900 44324 11902
rect 44268 11618 44324 11620
rect 44268 11566 44270 11618
rect 44270 11566 44322 11618
rect 44322 11566 44324 11618
rect 44268 11564 44324 11566
rect 44044 10668 44100 10724
rect 43708 10444 43764 10500
rect 43372 10332 43428 10388
rect 43372 7980 43428 8036
rect 43036 6860 43092 6916
rect 43484 6860 43540 6916
rect 43484 6524 43540 6580
rect 43036 6412 43092 6468
rect 42924 5794 42980 5796
rect 42924 5742 42926 5794
rect 42926 5742 42978 5794
rect 42978 5742 42980 5794
rect 42924 5740 42980 5742
rect 43260 6466 43316 6468
rect 43260 6414 43262 6466
rect 43262 6414 43314 6466
rect 43314 6414 43316 6466
rect 43260 6412 43316 6414
rect 43148 5234 43204 5236
rect 43148 5182 43150 5234
rect 43150 5182 43202 5234
rect 43202 5182 43204 5234
rect 43148 5180 43204 5182
rect 43484 4732 43540 4788
rect 43820 6188 43876 6244
rect 44044 5964 44100 6020
rect 44268 5964 44324 6020
rect 44044 5180 44100 5236
rect 45052 15874 45108 15876
rect 45052 15822 45054 15874
rect 45054 15822 45106 15874
rect 45106 15822 45108 15874
rect 45052 15820 45108 15822
rect 45836 17442 45892 17444
rect 45836 17390 45838 17442
rect 45838 17390 45890 17442
rect 45890 17390 45892 17442
rect 45836 17388 45892 17390
rect 45948 16716 46004 16772
rect 45388 14530 45444 14532
rect 45388 14478 45390 14530
rect 45390 14478 45442 14530
rect 45442 14478 45444 14530
rect 45388 14476 45444 14478
rect 46172 18956 46228 19012
rect 46284 17666 46340 17668
rect 46284 17614 46286 17666
rect 46286 17614 46338 17666
rect 46338 17614 46340 17666
rect 46284 17612 46340 17614
rect 46732 21586 46788 21588
rect 46732 21534 46734 21586
rect 46734 21534 46786 21586
rect 46786 21534 46788 21586
rect 46732 21532 46788 21534
rect 47516 21586 47572 21588
rect 47516 21534 47518 21586
rect 47518 21534 47570 21586
rect 47570 21534 47572 21586
rect 47516 21532 47572 21534
rect 48636 21532 48692 21588
rect 46844 20748 46900 20804
rect 46508 18562 46564 18564
rect 46508 18510 46510 18562
rect 46510 18510 46562 18562
rect 46562 18510 46564 18562
rect 46508 18508 46564 18510
rect 46732 19964 46788 20020
rect 46620 18284 46676 18340
rect 47068 20188 47124 20244
rect 47852 19292 47908 19348
rect 47852 18956 47908 19012
rect 46396 17052 46452 17108
rect 46060 14924 46116 14980
rect 44828 13580 44884 13636
rect 44604 10668 44660 10724
rect 44492 10108 44548 10164
rect 44716 11676 44772 11732
rect 44940 13468 44996 13524
rect 45836 14252 45892 14308
rect 45164 13020 45220 13076
rect 45500 13132 45556 13188
rect 48748 20188 48804 20244
rect 48748 19852 48804 19908
rect 48748 18844 48804 18900
rect 47852 17836 47908 17892
rect 47516 16770 47572 16772
rect 47516 16718 47518 16770
rect 47518 16718 47570 16770
rect 47570 16718 47572 16770
rect 47516 16716 47572 16718
rect 47964 17106 48020 17108
rect 47964 17054 47966 17106
rect 47966 17054 48018 17106
rect 48018 17054 48020 17106
rect 47964 17052 48020 17054
rect 47068 16492 47124 16548
rect 48636 17836 48692 17892
rect 47068 16156 47124 16212
rect 46732 14476 46788 14532
rect 46732 13916 46788 13972
rect 46060 12962 46116 12964
rect 46060 12910 46062 12962
rect 46062 12910 46114 12962
rect 46114 12910 46116 12962
rect 46060 12908 46116 12910
rect 46172 12738 46228 12740
rect 46172 12686 46174 12738
rect 46174 12686 46226 12738
rect 46226 12686 46228 12738
rect 46172 12684 46228 12686
rect 45388 12572 45444 12628
rect 45164 12460 45220 12516
rect 44604 9772 44660 9828
rect 45388 11228 45444 11284
rect 46284 12348 46340 12404
rect 46508 12460 46564 12516
rect 47740 14588 47796 14644
rect 46956 13692 47012 13748
rect 46844 13132 46900 13188
rect 48412 16210 48468 16212
rect 48412 16158 48414 16210
rect 48414 16158 48466 16210
rect 48466 16158 48468 16210
rect 48412 16156 48468 16158
rect 49420 21644 49476 21700
rect 49084 20130 49140 20132
rect 49084 20078 49086 20130
rect 49086 20078 49138 20130
rect 49138 20078 49140 20130
rect 49084 20076 49140 20078
rect 49196 19346 49252 19348
rect 49196 19294 49198 19346
rect 49198 19294 49250 19346
rect 49250 19294 49252 19346
rect 49196 19292 49252 19294
rect 49196 17836 49252 17892
rect 49084 16604 49140 16660
rect 48860 15260 48916 15316
rect 49084 14812 49140 14868
rect 49196 14642 49252 14644
rect 49196 14590 49198 14642
rect 49198 14590 49250 14642
rect 49250 14590 49252 14642
rect 49196 14588 49252 14590
rect 48860 13858 48916 13860
rect 48860 13806 48862 13858
rect 48862 13806 48914 13858
rect 48914 13806 48916 13858
rect 48860 13804 48916 13806
rect 48076 13746 48132 13748
rect 48076 13694 48078 13746
rect 48078 13694 48130 13746
rect 48130 13694 48132 13746
rect 48076 13692 48132 13694
rect 47964 13468 48020 13524
rect 47068 12684 47124 12740
rect 45836 12124 45892 12180
rect 45948 12066 46004 12068
rect 45948 12014 45950 12066
rect 45950 12014 46002 12066
rect 46002 12014 46004 12066
rect 45948 12012 46004 12014
rect 45388 10556 45444 10612
rect 45276 10332 45332 10388
rect 44828 9938 44884 9940
rect 44828 9886 44830 9938
rect 44830 9886 44882 9938
rect 44882 9886 44884 9938
rect 44828 9884 44884 9886
rect 45052 9826 45108 9828
rect 45052 9774 45054 9826
rect 45054 9774 45106 9826
rect 45106 9774 45108 9826
rect 45052 9772 45108 9774
rect 46060 10610 46116 10612
rect 46060 10558 46062 10610
rect 46062 10558 46114 10610
rect 46114 10558 46116 10610
rect 46060 10556 46116 10558
rect 45836 9602 45892 9604
rect 45836 9550 45838 9602
rect 45838 9550 45890 9602
rect 45890 9550 45892 9602
rect 45836 9548 45892 9550
rect 45500 8764 45556 8820
rect 44828 6636 44884 6692
rect 44828 6188 44884 6244
rect 44716 6076 44772 6132
rect 44380 5180 44436 5236
rect 43932 4732 43988 4788
rect 44156 4844 44212 4900
rect 44380 4450 44436 4452
rect 44380 4398 44382 4450
rect 44382 4398 44434 4450
rect 44434 4398 44436 4450
rect 44380 4396 44436 4398
rect 44492 3836 44548 3892
rect 43036 3442 43092 3444
rect 43036 3390 43038 3442
rect 43038 3390 43090 3442
rect 43090 3390 43092 3442
rect 43036 3388 43092 3390
rect 42364 3276 42420 3332
rect 44044 3554 44100 3556
rect 44044 3502 44046 3554
rect 44046 3502 44098 3554
rect 44098 3502 44100 3554
rect 44044 3500 44100 3502
rect 45724 8034 45780 8036
rect 45724 7982 45726 8034
rect 45726 7982 45778 8034
rect 45778 7982 45780 8034
rect 45724 7980 45780 7982
rect 45612 7532 45668 7588
rect 45948 8876 46004 8932
rect 45948 8428 46004 8484
rect 46508 9212 46564 9268
rect 46732 10722 46788 10724
rect 46732 10670 46734 10722
rect 46734 10670 46786 10722
rect 46786 10670 46788 10722
rect 46732 10668 46788 10670
rect 47068 12012 47124 12068
rect 46956 10444 47012 10500
rect 46844 10386 46900 10388
rect 46844 10334 46846 10386
rect 46846 10334 46898 10386
rect 46898 10334 46900 10386
rect 46844 10332 46900 10334
rect 47068 9938 47124 9940
rect 47068 9886 47070 9938
rect 47070 9886 47122 9938
rect 47122 9886 47124 9938
rect 47068 9884 47124 9886
rect 47516 12348 47572 12404
rect 47740 12236 47796 12292
rect 47852 13020 47908 13076
rect 47628 11676 47684 11732
rect 47964 12908 48020 12964
rect 48300 13020 48356 13076
rect 47964 11564 48020 11620
rect 47292 11340 47348 11396
rect 47292 10220 47348 10276
rect 48076 10780 48132 10836
rect 47628 10332 47684 10388
rect 47852 9324 47908 9380
rect 46396 9100 46452 9156
rect 46396 8428 46452 8484
rect 45948 7644 46004 7700
rect 45388 7196 45444 7252
rect 45164 6412 45220 6468
rect 45164 5852 45220 5908
rect 45276 6524 45332 6580
rect 45052 5628 45108 5684
rect 44940 4844 44996 4900
rect 45388 6466 45444 6468
rect 45388 6414 45390 6466
rect 45390 6414 45442 6466
rect 45442 6414 45444 6466
rect 45388 6412 45444 6414
rect 45388 6188 45444 6244
rect 45612 6524 45668 6580
rect 46284 6524 46340 6580
rect 46396 7980 46452 8036
rect 45724 6076 45780 6132
rect 45500 5964 45556 6020
rect 46620 7644 46676 7700
rect 46844 8764 46900 8820
rect 46508 6636 46564 6692
rect 47068 9042 47124 9044
rect 47068 8990 47070 9042
rect 47070 8990 47122 9042
rect 47122 8990 47124 9042
rect 47068 8988 47124 8990
rect 48076 9100 48132 9156
rect 46956 7532 47012 7588
rect 47852 9042 47908 9044
rect 47852 8990 47854 9042
rect 47854 8990 47906 9042
rect 47906 8990 47908 9042
rect 47852 8988 47908 8990
rect 47628 8764 47684 8820
rect 48524 13468 48580 13524
rect 48748 12348 48804 12404
rect 49644 20076 49700 20132
rect 49084 12850 49140 12852
rect 49084 12798 49086 12850
rect 49086 12798 49138 12850
rect 49138 12798 49140 12850
rect 49084 12796 49140 12798
rect 49644 12460 49700 12516
rect 49196 12236 49252 12292
rect 49084 12178 49140 12180
rect 49084 12126 49086 12178
rect 49086 12126 49138 12178
rect 49138 12126 49140 12178
rect 49084 12124 49140 12126
rect 48748 11564 48804 11620
rect 49084 11676 49140 11732
rect 49196 11340 49252 11396
rect 49420 12124 49476 12180
rect 48972 10722 49028 10724
rect 48972 10670 48974 10722
rect 48974 10670 49026 10722
rect 49026 10670 49028 10722
rect 48972 10668 49028 10670
rect 48524 10444 48580 10500
rect 48412 7532 48468 7588
rect 47516 7420 47572 7476
rect 47404 6748 47460 6804
rect 47292 6636 47348 6692
rect 46060 5234 46116 5236
rect 46060 5182 46062 5234
rect 46062 5182 46114 5234
rect 46114 5182 46116 5234
rect 46060 5180 46116 5182
rect 44828 4508 44884 4564
rect 45948 4844 46004 4900
rect 44828 3500 44884 3556
rect 43932 3164 43988 3220
rect 45612 2828 45668 2884
rect 46956 5964 47012 6020
rect 46508 4172 46564 4228
rect 46844 5852 46900 5908
rect 47740 6188 47796 6244
rect 48860 9884 48916 9940
rect 49084 9324 49140 9380
rect 48748 9154 48804 9156
rect 48748 9102 48750 9154
rect 48750 9102 48802 9154
rect 48802 9102 48804 9154
rect 48748 9100 48804 9102
rect 48748 8876 48804 8932
rect 48860 8092 48916 8148
rect 48748 7250 48804 7252
rect 48748 7198 48750 7250
rect 48750 7198 48802 7250
rect 48802 7198 48804 7250
rect 48748 7196 48804 7198
rect 48188 5964 48244 6020
rect 47628 5628 47684 5684
rect 47516 4956 47572 5012
rect 47740 4226 47796 4228
rect 47740 4174 47742 4226
rect 47742 4174 47794 4226
rect 47794 4174 47796 4226
rect 47740 4172 47796 4174
rect 47628 3724 47684 3780
rect 48076 3836 48132 3892
rect 48972 7420 49028 7476
rect 49196 8988 49252 9044
rect 49196 7644 49252 7700
rect 49644 10668 49700 10724
rect 49308 7420 49364 7476
rect 49532 10220 49588 10276
rect 48972 6412 49028 6468
rect 49196 6300 49252 6356
rect 48972 6188 49028 6244
rect 48748 4732 48804 4788
rect 48636 3724 48692 3780
rect 48748 3666 48804 3668
rect 48748 3614 48750 3666
rect 48750 3614 48802 3666
rect 48802 3614 48804 3666
rect 48748 3612 48804 3614
rect 48076 3330 48132 3332
rect 48076 3278 48078 3330
rect 48078 3278 48130 3330
rect 48130 3278 48132 3330
rect 48076 3276 48132 3278
rect 49308 6076 49364 6132
rect 49196 4620 49252 4676
rect 48972 2716 49028 2772
rect 49196 2268 49252 2324
<< metal3 >>
rect 50200 48916 51000 48944
rect 48178 48860 48188 48916
rect 48244 48860 51000 48916
rect 50200 48832 51000 48860
rect 33730 47964 33740 48020
rect 33796 47964 48188 48020
rect 48244 47964 48254 48020
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 40012 47628 42364 47684
rect 42420 47628 45388 47684
rect 45444 47628 47516 47684
rect 47572 47628 47582 47684
rect 40012 47460 40068 47628
rect 40562 47516 40572 47572
rect 40628 47516 44828 47572
rect 44884 47516 44894 47572
rect 37762 47404 37772 47460
rect 37828 47404 40012 47460
rect 40068 47404 40078 47460
rect 41234 47404 41244 47460
rect 41300 47404 41916 47460
rect 41972 47404 41982 47460
rect 42130 47404 42140 47460
rect 42196 47404 44156 47460
rect 44212 47404 44222 47460
rect 15810 47292 15820 47348
rect 15876 47292 19852 47348
rect 19908 47292 19918 47348
rect 38770 47292 38780 47348
rect 38836 47292 46844 47348
rect 46900 47292 49084 47348
rect 49140 47292 49150 47348
rect 35186 47180 35196 47236
rect 35252 47180 35980 47236
rect 36036 47180 36046 47236
rect 36866 47180 36876 47236
rect 36932 47180 40348 47236
rect 40404 47180 41020 47236
rect 41076 47180 41086 47236
rect 41346 47180 41356 47236
rect 41412 47180 45724 47236
rect 45780 47180 46172 47236
rect 46228 47180 46238 47236
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 32274 46956 32284 47012
rect 32340 46956 48748 47012
rect 48804 46956 48814 47012
rect 6290 46844 6300 46900
rect 6356 46844 11900 46900
rect 11956 46844 11966 46900
rect 34178 46844 34188 46900
rect 34244 46844 37772 46900
rect 37828 46844 37838 46900
rect 6626 46732 6636 46788
rect 6692 46732 8428 46788
rect 8484 46732 9548 46788
rect 9604 46732 9614 46788
rect 23874 46620 23884 46676
rect 23940 46620 25228 46676
rect 25284 46620 25294 46676
rect 32162 46620 32172 46676
rect 32228 46620 34412 46676
rect 34468 46620 34478 46676
rect 41010 46620 41020 46676
rect 41076 46620 41356 46676
rect 41412 46620 44380 46676
rect 44436 46620 44446 46676
rect 3378 46508 3388 46564
rect 3444 46508 7084 46564
rect 7140 46508 7150 46564
rect 7298 46508 7308 46564
rect 7364 46508 8092 46564
rect 8148 46508 8158 46564
rect 24994 46396 25004 46452
rect 25060 46396 47740 46452
rect 47796 46396 47806 46452
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 30258 46172 30268 46228
rect 30324 46172 32060 46228
rect 32116 46172 32126 46228
rect 41682 46172 41692 46228
rect 41748 46172 44268 46228
rect 44324 46172 45836 46228
rect 45892 46172 45902 46228
rect 41570 46060 41580 46116
rect 41636 46060 45388 46116
rect 45444 46060 45454 46116
rect 28914 45948 28924 46004
rect 28980 45948 31948 46004
rect 32004 45948 32014 46004
rect 43026 45948 43036 46004
rect 43092 45948 45836 46004
rect 45892 45948 46732 46004
rect 46788 45948 47180 46004
rect 47236 45948 47246 46004
rect 6290 45836 6300 45892
rect 6356 45836 7756 45892
rect 7812 45836 7822 45892
rect 26562 45836 26572 45892
rect 26628 45836 27356 45892
rect 27412 45836 27422 45892
rect 27570 45836 27580 45892
rect 27636 45836 29148 45892
rect 29204 45836 29214 45892
rect 30594 45836 30604 45892
rect 30660 45836 31276 45892
rect 31332 45836 31342 45892
rect 41794 45836 41804 45892
rect 41860 45836 42588 45892
rect 42644 45836 43932 45892
rect 43988 45836 43998 45892
rect 44370 45836 44380 45892
rect 44436 45836 45276 45892
rect 45332 45836 49084 45892
rect 49140 45836 49150 45892
rect 3042 45724 3052 45780
rect 3108 45724 4396 45780
rect 4452 45724 4462 45780
rect 4946 45724 4956 45780
rect 5012 45724 7196 45780
rect 7252 45724 7262 45780
rect 26674 45724 26684 45780
rect 26740 45724 28028 45780
rect 28084 45724 28094 45780
rect 6038 45612 6076 45668
rect 6132 45612 7308 45668
rect 7364 45612 7374 45668
rect 43474 45612 43484 45668
rect 43540 45612 44828 45668
rect 44884 45612 44894 45668
rect 43026 45500 43036 45556
rect 43092 45500 43820 45556
rect 43876 45500 43886 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 41458 45388 41468 45444
rect 41524 45388 43652 45444
rect 43596 45332 43652 45388
rect 26450 45276 26460 45332
rect 26516 45276 26796 45332
rect 26852 45276 28140 45332
rect 28196 45276 28206 45332
rect 43596 45276 48412 45332
rect 48468 45276 48478 45332
rect 18386 45164 18396 45220
rect 18452 45164 21644 45220
rect 21700 45164 21710 45220
rect 26898 45164 26908 45220
rect 26964 45164 27916 45220
rect 27972 45164 29932 45220
rect 29988 45164 32956 45220
rect 33012 45164 33022 45220
rect 33394 45164 33404 45220
rect 33460 45164 35196 45220
rect 35252 45164 37100 45220
rect 37156 45164 37166 45220
rect 45714 45164 45724 45220
rect 45780 45164 46620 45220
rect 46676 45164 46686 45220
rect 28588 45108 28644 45164
rect 7186 45052 7196 45108
rect 7252 45052 7756 45108
rect 7812 45052 8988 45108
rect 9044 45052 9054 45108
rect 25554 45052 25564 45108
rect 25620 45052 27020 45108
rect 27076 45052 27086 45108
rect 28578 45052 28588 45108
rect 28644 45052 28654 45108
rect 30930 45052 30940 45108
rect 30996 45052 32172 45108
rect 32228 45052 32238 45108
rect 33618 45052 33628 45108
rect 33684 45052 35084 45108
rect 35140 45052 36204 45108
rect 36260 45052 37212 45108
rect 37268 45052 37278 45108
rect 5170 44940 5180 44996
rect 5236 44940 5852 44996
rect 5908 44940 6748 44996
rect 6804 44940 6814 44996
rect 30594 44940 30604 44996
rect 30660 44940 32396 44996
rect 32452 44940 34188 44996
rect 34244 44940 34254 44996
rect 41346 44940 41356 44996
rect 41412 44940 42700 44996
rect 42756 44940 43260 44996
rect 43316 44940 43326 44996
rect 31266 44828 31276 44884
rect 31332 44828 31724 44884
rect 31780 44828 33852 44884
rect 33908 44828 33918 44884
rect 35074 44828 35084 44884
rect 35140 44828 37324 44884
rect 37380 44828 37390 44884
rect 42578 44828 42588 44884
rect 42644 44828 46060 44884
rect 46116 44828 46126 44884
rect 45378 44716 45388 44772
rect 45444 44716 45948 44772
rect 46004 44716 46014 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 38322 44604 38332 44660
rect 38388 44604 38668 44660
rect 46610 44604 46620 44660
rect 46676 44604 47180 44660
rect 47236 44604 47246 44660
rect 30818 44492 30828 44548
rect 30884 44492 35868 44548
rect 35924 44492 35934 44548
rect 38612 44436 38668 44604
rect 50200 44576 51000 44688
rect 42466 44492 42476 44548
rect 42532 44492 47292 44548
rect 47348 44492 47358 44548
rect 18498 44380 18508 44436
rect 18564 44380 21980 44436
rect 22036 44380 22046 44436
rect 24546 44380 24556 44436
rect 24612 44380 25228 44436
rect 25284 44380 25294 44436
rect 26674 44380 26684 44436
rect 26740 44380 27916 44436
rect 27972 44380 27982 44436
rect 32498 44380 32508 44436
rect 32564 44380 33740 44436
rect 33796 44380 33806 44436
rect 34738 44380 34748 44436
rect 34804 44380 36988 44436
rect 37044 44380 37054 44436
rect 37202 44380 37212 44436
rect 37268 44380 38332 44436
rect 38388 44380 38398 44436
rect 38612 44380 41132 44436
rect 41188 44380 41198 44436
rect 42354 44380 42364 44436
rect 42420 44380 46564 44436
rect 46508 44324 46564 44380
rect 4610 44268 4620 44324
rect 4676 44268 5740 44324
rect 5796 44268 5806 44324
rect 16482 44268 16492 44324
rect 16548 44268 18396 44324
rect 18452 44268 18462 44324
rect 42914 44268 42924 44324
rect 42980 44268 43820 44324
rect 43876 44268 43886 44324
rect 44044 44268 44940 44324
rect 44996 44268 45006 44324
rect 45798 44268 45836 44324
rect 45892 44268 45902 44324
rect 46498 44268 46508 44324
rect 46564 44268 47516 44324
rect 47572 44268 47582 44324
rect 44044 44212 44100 44268
rect 20290 44156 20300 44212
rect 20356 44156 22316 44212
rect 22372 44156 22382 44212
rect 39890 44156 39900 44212
rect 39956 44156 43596 44212
rect 43652 44156 44100 44212
rect 44258 44156 44268 44212
rect 44324 44156 45052 44212
rect 45108 44156 45118 44212
rect 21634 44044 21644 44100
rect 21700 44044 22428 44100
rect 22484 44044 25900 44100
rect 25956 44044 25966 44100
rect 27122 44044 27132 44100
rect 27188 44044 27916 44100
rect 27972 44044 28252 44100
rect 28308 44044 28318 44100
rect 33170 44044 33180 44100
rect 33236 44044 33740 44100
rect 33796 44044 33806 44100
rect 38612 44044 40460 44100
rect 40516 44044 44044 44100
rect 44100 44044 44828 44100
rect 44884 44044 44894 44100
rect 5842 43932 5852 43988
rect 5908 43932 6188 43988
rect 6244 43932 6254 43988
rect 6402 43932 6412 43988
rect 6468 43932 7084 43988
rect 7140 43932 7150 43988
rect 35970 43932 35980 43988
rect 36036 43932 36988 43988
rect 37044 43932 37054 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 38612 43876 38668 44044
rect 6038 43820 6076 43876
rect 6132 43820 6142 43876
rect 37090 43820 37100 43876
rect 37156 43820 38668 43876
rect 41010 43820 41020 43876
rect 41076 43820 41468 43876
rect 41524 43820 41534 43876
rect 5730 43708 5740 43764
rect 5796 43708 7644 43764
rect 7700 43708 7710 43764
rect 32946 43708 32956 43764
rect 33012 43708 33740 43764
rect 33796 43708 33806 43764
rect 43922 43708 43932 43764
rect 43988 43708 44716 43764
rect 44772 43708 44782 43764
rect 3490 43596 3500 43652
rect 3556 43596 4676 43652
rect 4834 43596 4844 43652
rect 4900 43596 5628 43652
rect 5684 43596 7420 43652
rect 7476 43596 7486 43652
rect 23090 43596 23100 43652
rect 23156 43596 23660 43652
rect 23716 43596 23726 43652
rect 34850 43596 34860 43652
rect 34916 43596 35420 43652
rect 35476 43596 35980 43652
rect 36036 43596 36046 43652
rect 44482 43596 44492 43652
rect 44548 43596 48636 43652
rect 48692 43596 48702 43652
rect 4620 43540 4676 43596
rect 3042 43484 3052 43540
rect 3108 43484 3948 43540
rect 4004 43484 4014 43540
rect 4620 43484 7084 43540
rect 7140 43484 8540 43540
rect 8596 43484 8606 43540
rect 8866 43484 8876 43540
rect 8932 43484 10444 43540
rect 10500 43484 11228 43540
rect 11284 43484 12012 43540
rect 12068 43484 12078 43540
rect 27794 43484 27804 43540
rect 27860 43484 28028 43540
rect 28084 43484 29932 43540
rect 29988 43484 29998 43540
rect 31602 43484 31612 43540
rect 31668 43484 32620 43540
rect 32676 43484 32686 43540
rect 35186 43484 35196 43540
rect 35252 43484 35756 43540
rect 35812 43484 35822 43540
rect 36530 43484 36540 43540
rect 36596 43484 38332 43540
rect 38388 43484 38398 43540
rect 44818 43484 44828 43540
rect 44884 43484 46508 43540
rect 46564 43484 46574 43540
rect 8540 43428 8596 43484
rect 3266 43372 3276 43428
rect 3332 43372 7532 43428
rect 7588 43372 7598 43428
rect 8540 43372 9772 43428
rect 9828 43372 10780 43428
rect 10836 43372 10846 43428
rect 24546 43372 24556 43428
rect 24612 43372 27580 43428
rect 27636 43372 27646 43428
rect 28130 43372 28140 43428
rect 28196 43372 29148 43428
rect 29204 43372 29214 43428
rect 31938 43372 31948 43428
rect 32004 43372 33068 43428
rect 33124 43372 33134 43428
rect 33506 43372 33516 43428
rect 33572 43372 35084 43428
rect 35140 43372 35150 43428
rect 35634 43372 35644 43428
rect 35700 43372 37212 43428
rect 37268 43372 37278 43428
rect 41682 43372 41692 43428
rect 41748 43372 42588 43428
rect 42644 43372 42654 43428
rect 46162 43372 46172 43428
rect 46228 43372 47180 43428
rect 47236 43372 47246 43428
rect 47954 43372 47964 43428
rect 48020 43372 48860 43428
rect 48916 43372 48926 43428
rect 2482 43260 2492 43316
rect 2548 43260 3836 43316
rect 3892 43260 3902 43316
rect 4162 43260 4172 43316
rect 4228 43260 8092 43316
rect 8148 43260 8158 43316
rect 8418 43260 8428 43316
rect 8484 43260 10444 43316
rect 10500 43260 10510 43316
rect 27346 43260 27356 43316
rect 27412 43260 28364 43316
rect 28420 43260 29372 43316
rect 29428 43260 29438 43316
rect 30370 43260 30380 43316
rect 30436 43260 30828 43316
rect 30884 43260 36652 43316
rect 36708 43260 37100 43316
rect 37156 43260 37772 43316
rect 37828 43260 37838 43316
rect 42130 43260 42140 43316
rect 42196 43260 42206 43316
rect 44258 43260 44268 43316
rect 44324 43260 45052 43316
rect 45108 43260 45118 43316
rect 45826 43260 45836 43316
rect 45892 43260 46956 43316
rect 47012 43260 48076 43316
rect 48132 43260 48142 43316
rect 42140 43204 42196 43260
rect 4946 43148 4956 43204
rect 5012 43148 5292 43204
rect 5348 43148 8204 43204
rect 8260 43148 8270 43204
rect 25890 43148 25900 43204
rect 25956 43148 27692 43204
rect 27748 43148 27758 43204
rect 28914 43148 28924 43204
rect 28980 43148 31836 43204
rect 31892 43148 31902 43204
rect 32274 43148 32284 43204
rect 32340 43148 32676 43204
rect 37538 43148 37548 43204
rect 37604 43148 38108 43204
rect 38164 43148 38174 43204
rect 38658 43148 38668 43204
rect 38724 43148 40348 43204
rect 40404 43148 43372 43204
rect 43428 43148 43438 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 6300 43092 6356 43148
rect 6290 43036 6300 43092
rect 6356 43036 6366 43092
rect 28242 43036 28252 43092
rect 28308 43036 29036 43092
rect 29092 43036 31164 43092
rect 31220 43036 31230 43092
rect 6402 42924 6412 42980
rect 6468 42924 6860 42980
rect 6916 42924 11564 42980
rect 11620 42924 11630 42980
rect 20178 42924 20188 42980
rect 20244 42924 21532 42980
rect 21588 42924 22876 42980
rect 22932 42924 22942 42980
rect 27906 42924 27916 42980
rect 27972 42924 28476 42980
rect 28532 42924 29148 42980
rect 29204 42924 29214 42980
rect 5058 42812 5068 42868
rect 5124 42812 6076 42868
rect 6132 42812 8428 42868
rect 8484 42812 8494 42868
rect 9874 42812 9884 42868
rect 9940 42812 10836 42868
rect 19170 42812 19180 42868
rect 19236 42812 21196 42868
rect 21252 42812 21868 42868
rect 21924 42812 21934 42868
rect 26898 42812 26908 42868
rect 26964 42812 27244 42868
rect 27300 42812 29260 42868
rect 29316 42812 29326 42868
rect 10780 42756 10836 42812
rect 32620 42756 32676 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 35858 42924 35868 42980
rect 35924 42924 37548 42980
rect 37604 42924 37614 42980
rect 38612 42924 38780 42980
rect 38836 42924 38846 42980
rect 44482 42924 44492 42980
rect 44548 42924 45388 42980
rect 45444 42924 45454 42980
rect 34738 42812 34748 42868
rect 34804 42812 34972 42868
rect 35028 42812 35038 42868
rect 8866 42700 8876 42756
rect 8932 42700 10332 42756
rect 10388 42700 10398 42756
rect 10770 42700 10780 42756
rect 10836 42700 11452 42756
rect 11508 42700 12124 42756
rect 12180 42700 12190 42756
rect 22306 42700 22316 42756
rect 22372 42700 26796 42756
rect 8194 42588 8204 42644
rect 8260 42588 10220 42644
rect 10276 42588 10286 42644
rect 15138 42588 15148 42644
rect 15204 42588 16492 42644
rect 16548 42588 16558 42644
rect 20066 42588 20076 42644
rect 20132 42588 22204 42644
rect 22260 42588 22270 42644
rect 22530 42588 22540 42644
rect 22596 42588 22988 42644
rect 23044 42588 23436 42644
rect 23492 42588 23502 42644
rect 18246 42476 18284 42532
rect 18340 42476 18350 42532
rect 18610 42476 18620 42532
rect 18676 42476 19068 42532
rect 19124 42476 19134 42532
rect 22082 42476 22092 42532
rect 22148 42476 23100 42532
rect 23156 42476 23166 42532
rect 23314 42476 23324 42532
rect 23380 42476 25452 42532
rect 25508 42476 25518 42532
rect 26852 42476 26908 42756
rect 30594 42700 30604 42756
rect 30660 42700 31948 42756
rect 32004 42700 32014 42756
rect 32610 42700 32620 42756
rect 32676 42700 32686 42756
rect 33842 42700 33852 42756
rect 33908 42700 35308 42756
rect 35364 42700 35374 42756
rect 38612 42644 38668 42924
rect 48626 42812 48636 42868
rect 48692 42812 49196 42868
rect 49252 42812 49262 42868
rect 41794 42700 41804 42756
rect 41860 42700 42476 42756
rect 42532 42700 42542 42756
rect 42802 42700 42812 42756
rect 42868 42700 43596 42756
rect 43652 42700 43662 42756
rect 31042 42588 31052 42644
rect 31108 42588 32452 42644
rect 32396 42532 32452 42588
rect 38332 42588 39116 42644
rect 39172 42588 39182 42644
rect 42690 42588 42700 42644
rect 42756 42588 45052 42644
rect 45108 42588 45118 42644
rect 26964 42476 26974 42532
rect 31602 42476 31612 42532
rect 31668 42476 32172 42532
rect 32228 42476 32238 42532
rect 32396 42476 32732 42532
rect 32788 42476 32798 42532
rect 33058 42476 33068 42532
rect 33124 42476 33740 42532
rect 33796 42476 33806 42532
rect 36390 42476 36428 42532
rect 36484 42476 36494 42532
rect 23324 42420 23380 42476
rect 21634 42364 21644 42420
rect 21700 42364 23380 42420
rect 26908 42420 26964 42476
rect 38332 42420 38388 42588
rect 38546 42476 38556 42532
rect 38612 42476 40348 42532
rect 40404 42476 40414 42532
rect 26908 42364 38444 42420
rect 38500 42364 38510 42420
rect 43586 42364 43596 42420
rect 43652 42364 45052 42420
rect 45108 42364 45118 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 27906 42252 27916 42308
rect 27972 42252 37660 42308
rect 37716 42252 40796 42308
rect 40852 42252 40862 42308
rect 7970 42140 7980 42196
rect 8036 42140 8316 42196
rect 8372 42140 9660 42196
rect 9716 42140 9726 42196
rect 18722 42140 18732 42196
rect 18788 42140 18798 42196
rect 31154 42140 31164 42196
rect 31220 42140 31612 42196
rect 31668 42140 31678 42196
rect 31826 42140 31836 42196
rect 31892 42140 32396 42196
rect 32452 42140 32956 42196
rect 33012 42140 33022 42196
rect 34402 42140 34412 42196
rect 34468 42140 35868 42196
rect 35924 42140 35934 42196
rect 36866 42140 36876 42196
rect 36932 42140 37660 42196
rect 37716 42140 38668 42196
rect 38724 42140 39676 42196
rect 39732 42140 41244 42196
rect 41300 42140 41310 42196
rect 41804 42140 44156 42196
rect 44212 42140 44222 42196
rect 18732 41972 18788 42140
rect 27906 42028 27916 42084
rect 27972 42028 30492 42084
rect 30548 42028 30558 42084
rect 30706 42028 30716 42084
rect 30772 42028 31276 42084
rect 31332 42028 31342 42084
rect 36194 42028 36204 42084
rect 36260 42028 37436 42084
rect 37492 42028 37502 42084
rect 6626 41916 6636 41972
rect 6692 41916 8652 41972
rect 8708 41916 12684 41972
rect 12740 41916 18284 41972
rect 18340 41916 23436 41972
rect 23492 41916 25228 41972
rect 25284 41916 25294 41972
rect 29474 41916 29484 41972
rect 29540 41916 31388 41972
rect 31444 41916 31454 41972
rect 38098 41916 38108 41972
rect 38164 41916 38444 41972
rect 38500 41916 39228 41972
rect 39284 41916 39294 41972
rect 39452 41916 40292 41972
rect 39452 41860 39508 41916
rect 40236 41860 40292 41916
rect 41804 41860 41860 42140
rect 43250 42028 43260 42084
rect 43316 42028 44940 42084
rect 44996 42028 45006 42084
rect 43026 41916 43036 41972
rect 43092 41916 44716 41972
rect 44772 41916 44782 41972
rect 46498 41916 46508 41972
rect 46564 41916 47180 41972
rect 47236 41916 47246 41972
rect 16370 41804 16380 41860
rect 16436 41804 16940 41860
rect 16996 41804 17500 41860
rect 17556 41804 17566 41860
rect 24098 41804 24108 41860
rect 24164 41804 27244 41860
rect 27300 41804 27310 41860
rect 32386 41804 32396 41860
rect 32452 41804 33516 41860
rect 33572 41804 33582 41860
rect 34738 41804 34748 41860
rect 34804 41804 35084 41860
rect 35140 41804 35150 41860
rect 38210 41804 38220 41860
rect 38276 41804 39508 41860
rect 40226 41804 40236 41860
rect 40292 41804 40302 41860
rect 41794 41804 41804 41860
rect 41860 41804 41870 41860
rect 44044 41804 45276 41860
rect 45332 41804 45342 41860
rect 48150 41804 48188 41860
rect 48244 41804 48254 41860
rect 44044 41748 44100 41804
rect 18610 41692 18620 41748
rect 18676 41692 19292 41748
rect 19348 41692 19358 41748
rect 23100 41692 23548 41748
rect 23604 41692 30156 41748
rect 30212 41692 30222 41748
rect 33282 41692 33292 41748
rect 33348 41692 34188 41748
rect 34244 41692 34254 41748
rect 34850 41692 34860 41748
rect 34916 41692 37100 41748
rect 37156 41692 37166 41748
rect 37874 41692 37884 41748
rect 37940 41692 39676 41748
rect 39732 41692 39742 41748
rect 42354 41692 42364 41748
rect 42420 41692 44044 41748
rect 44100 41692 44110 41748
rect 44258 41692 44268 41748
rect 44324 41692 46396 41748
rect 46452 41692 46462 41748
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 23100 41524 23156 41692
rect 38546 41580 38556 41636
rect 38612 41580 39340 41636
rect 39396 41580 41132 41636
rect 41188 41580 41198 41636
rect 42242 41580 42252 41636
rect 42308 41580 44380 41636
rect 44436 41580 45500 41636
rect 45556 41580 45566 41636
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 23090 41468 23100 41524
rect 23156 41468 23166 41524
rect 43586 41468 43596 41524
rect 43652 41468 45388 41524
rect 45444 41468 45454 41524
rect 34290 41356 34300 41412
rect 34356 41356 36204 41412
rect 36260 41356 36270 41412
rect 16370 41244 16380 41300
rect 16436 41244 18844 41300
rect 18900 41244 20636 41300
rect 20692 41244 20702 41300
rect 28578 41244 28588 41300
rect 28644 41244 29372 41300
rect 29428 41244 29438 41300
rect 34066 41244 34076 41300
rect 34132 41244 34916 41300
rect 44258 41244 44268 41300
rect 44324 41244 49196 41300
rect 49252 41244 49420 41300
rect 49476 41244 49486 41300
rect 34860 41188 34916 41244
rect 9986 41132 9996 41188
rect 10052 41132 12460 41188
rect 12516 41132 13580 41188
rect 13636 41132 13646 41188
rect 16706 41132 16716 41188
rect 16772 41132 17612 41188
rect 17668 41132 18172 41188
rect 18228 41132 18238 41188
rect 24098 41132 24108 41188
rect 24164 41132 24780 41188
rect 24836 41132 25228 41188
rect 25284 41132 25294 41188
rect 31826 41132 31836 41188
rect 31892 41132 33628 41188
rect 33684 41132 33694 41188
rect 34850 41132 34860 41188
rect 34916 41132 35532 41188
rect 35588 41132 39004 41188
rect 39060 41132 39070 41188
rect 40450 41132 40460 41188
rect 40516 41132 41244 41188
rect 41300 41132 42140 41188
rect 42196 41132 42924 41188
rect 42980 41132 42990 41188
rect 45490 41132 45500 41188
rect 45556 41132 45948 41188
rect 46004 41132 46014 41188
rect 9874 41020 9884 41076
rect 9940 41020 11676 41076
rect 11732 41020 11742 41076
rect 17042 41020 17052 41076
rect 17108 41020 18732 41076
rect 18788 41020 18798 41076
rect 19730 41020 19740 41076
rect 19796 41020 21308 41076
rect 21364 41020 21374 41076
rect 30818 41020 30828 41076
rect 30884 41020 32284 41076
rect 32340 41020 32350 41076
rect 35186 41020 35196 41076
rect 35252 41020 35756 41076
rect 35812 41020 36876 41076
rect 36932 41020 36942 41076
rect 10546 40908 10556 40964
rect 10612 40908 12796 40964
rect 12852 40908 12862 40964
rect 17490 40908 17500 40964
rect 17556 40908 18508 40964
rect 18564 40908 18574 40964
rect 19954 40908 19964 40964
rect 20020 40908 20412 40964
rect 20468 40908 20478 40964
rect 33058 40908 33068 40964
rect 33124 40908 35420 40964
rect 35476 40908 35486 40964
rect 37090 40908 37100 40964
rect 37156 40908 38780 40964
rect 38836 40908 38846 40964
rect 42354 40908 42364 40964
rect 42420 40908 44716 40964
rect 44772 40908 44782 40964
rect 17500 40796 18284 40852
rect 18340 40796 18350 40852
rect 21298 40796 21308 40852
rect 21364 40796 22652 40852
rect 22708 40796 22718 40852
rect 25890 40796 25900 40852
rect 25956 40796 28196 40852
rect 33842 40796 33852 40852
rect 33908 40796 34860 40852
rect 34916 40796 34926 40852
rect 35186 40796 35196 40852
rect 35252 40796 38220 40852
rect 38276 40796 38286 40852
rect 45714 40796 45724 40852
rect 45780 40796 47516 40852
rect 47572 40796 47582 40852
rect 48850 40796 48860 40852
rect 48916 40796 49420 40852
rect 49476 40796 49486 40852
rect 17500 40740 17556 40796
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 28140 40740 28196 40796
rect 16594 40684 16604 40740
rect 16660 40684 17500 40740
rect 17556 40684 17566 40740
rect 17938 40684 17948 40740
rect 18004 40684 18014 40740
rect 26898 40684 26908 40740
rect 26964 40684 27692 40740
rect 27748 40684 27758 40740
rect 28130 40684 28140 40740
rect 28196 40684 37548 40740
rect 37604 40684 37614 40740
rect 6178 40572 6188 40628
rect 6244 40572 7756 40628
rect 7812 40572 8316 40628
rect 8372 40572 8382 40628
rect 4498 40460 4508 40516
rect 4564 40460 5068 40516
rect 5124 40460 5134 40516
rect 5394 40460 5404 40516
rect 5460 40460 5470 40516
rect 7634 40460 7644 40516
rect 7700 40460 8204 40516
rect 8260 40460 9548 40516
rect 9604 40460 9614 40516
rect 5404 40404 5460 40460
rect 2930 40348 2940 40404
rect 2996 40348 3724 40404
rect 3780 40348 3790 40404
rect 4610 40348 4620 40404
rect 4676 40348 6300 40404
rect 6356 40348 6366 40404
rect 17948 40292 18004 40684
rect 18610 40572 18620 40628
rect 18676 40572 20076 40628
rect 20132 40572 20142 40628
rect 26338 40572 26348 40628
rect 26404 40572 27580 40628
rect 27636 40572 27646 40628
rect 33282 40572 33292 40628
rect 33348 40572 34524 40628
rect 34580 40572 34590 40628
rect 38658 40572 38668 40628
rect 38724 40572 41020 40628
rect 41076 40572 41086 40628
rect 43362 40572 43372 40628
rect 43428 40572 45276 40628
rect 45332 40572 45342 40628
rect 22082 40460 22092 40516
rect 22148 40460 22428 40516
rect 22484 40460 25452 40516
rect 25508 40460 25518 40516
rect 30146 40460 30156 40516
rect 30212 40460 36092 40516
rect 36148 40460 36158 40516
rect 39442 40460 39452 40516
rect 39508 40460 41804 40516
rect 41860 40460 41870 40516
rect 42578 40460 42588 40516
rect 42644 40460 43820 40516
rect 43876 40460 43886 40516
rect 46834 40460 46844 40516
rect 46900 40460 49028 40516
rect 41804 40404 41860 40460
rect 48972 40404 49028 40460
rect 50200 40404 51000 40432
rect 18834 40348 18844 40404
rect 18900 40348 19740 40404
rect 19796 40348 19806 40404
rect 20290 40348 20300 40404
rect 20356 40348 21980 40404
rect 22036 40348 22046 40404
rect 34402 40348 34412 40404
rect 34468 40348 34972 40404
rect 35028 40348 35038 40404
rect 36418 40348 36428 40404
rect 36484 40348 37324 40404
rect 37380 40348 37390 40404
rect 37874 40348 37884 40404
rect 37940 40348 38108 40404
rect 38164 40348 39676 40404
rect 39732 40348 39742 40404
rect 41804 40348 42700 40404
rect 42756 40348 42766 40404
rect 42914 40348 42924 40404
rect 42980 40348 44156 40404
rect 44212 40348 45836 40404
rect 45892 40348 45902 40404
rect 47618 40348 47628 40404
rect 47684 40348 48748 40404
rect 48804 40348 48814 40404
rect 48972 40348 51000 40404
rect 50200 40320 51000 40348
rect 16146 40236 16156 40292
rect 16212 40236 18004 40292
rect 19954 40236 19964 40292
rect 20020 40236 20524 40292
rect 20580 40236 20590 40292
rect 24434 40236 24444 40292
rect 24500 40236 25788 40292
rect 25844 40236 25854 40292
rect 33954 40236 33964 40292
rect 34020 40236 36204 40292
rect 36260 40236 36540 40292
rect 36596 40236 36606 40292
rect 40898 40236 40908 40292
rect 40964 40236 41468 40292
rect 41524 40236 41534 40292
rect 47282 40236 47292 40292
rect 47348 40236 48972 40292
rect 49028 40236 49038 40292
rect 8866 40124 8876 40180
rect 8932 40124 9436 40180
rect 9492 40124 9502 40180
rect 18162 40124 18172 40180
rect 18228 40124 21420 40180
rect 21476 40124 21486 40180
rect 26786 40124 26796 40180
rect 26852 40124 27804 40180
rect 27860 40124 27870 40180
rect 35186 40124 35196 40180
rect 35252 40124 36988 40180
rect 37044 40124 37054 40180
rect 41906 40124 41916 40180
rect 41972 40124 43932 40180
rect 43988 40124 44940 40180
rect 44996 40124 45006 40180
rect 46722 40124 46732 40180
rect 46788 40124 48748 40180
rect 48804 40124 48814 40180
rect 5058 40012 5068 40068
rect 5124 40012 6076 40068
rect 6132 40012 6748 40068
rect 6804 40012 6814 40068
rect 17724 40012 17948 40068
rect 18004 40012 18014 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 17724 39956 17780 40012
rect 17714 39900 17724 39956
rect 17780 39900 17790 39956
rect 8530 39676 8540 39732
rect 8596 39676 8606 39732
rect 8540 39620 8596 39676
rect 4946 39564 4956 39620
rect 5012 39564 7532 39620
rect 7588 39564 7598 39620
rect 7746 39564 7756 39620
rect 7812 39564 9324 39620
rect 9380 39564 9390 39620
rect 14018 39564 14028 39620
rect 14084 39564 15036 39620
rect 15092 39564 15102 39620
rect 5842 39452 5852 39508
rect 5908 39452 8092 39508
rect 8148 39452 8540 39508
rect 8596 39452 8606 39508
rect 10210 39452 10220 39508
rect 10276 39452 11452 39508
rect 11508 39452 11518 39508
rect 14914 39452 14924 39508
rect 14980 39452 16156 39508
rect 16212 39452 16222 39508
rect 17042 39452 17052 39508
rect 17108 39452 17724 39508
rect 17780 39452 17790 39508
rect 18172 39396 18228 40124
rect 43148 40068 43204 40124
rect 43138 40012 43148 40068
rect 43204 40012 43214 40068
rect 47058 40012 47068 40068
rect 47124 40012 47964 40068
rect 48020 40012 49644 40068
rect 49700 40012 49710 40068
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 21186 39900 21196 39956
rect 21252 39900 22204 39956
rect 22260 39900 22270 39956
rect 24658 39900 24668 39956
rect 24724 39900 25676 39956
rect 25732 39900 26572 39956
rect 26628 39900 26638 39956
rect 20290 39788 20300 39844
rect 20356 39788 21084 39844
rect 21140 39788 21150 39844
rect 34626 39788 34636 39844
rect 34692 39788 35308 39844
rect 35364 39788 35374 39844
rect 39778 39788 39788 39844
rect 39844 39788 41244 39844
rect 41300 39788 41310 39844
rect 39218 39676 39228 39732
rect 39284 39676 41356 39732
rect 41412 39676 41422 39732
rect 43698 39676 43708 39732
rect 43764 39676 45724 39732
rect 45780 39676 47068 39732
rect 47124 39676 47134 39732
rect 20066 39564 20076 39620
rect 20132 39564 20636 39620
rect 20692 39564 20702 39620
rect 26226 39564 26236 39620
rect 26292 39564 26908 39620
rect 35522 39564 35532 39620
rect 35588 39564 35980 39620
rect 36036 39564 37212 39620
rect 37268 39564 37278 39620
rect 37538 39564 37548 39620
rect 37604 39564 41300 39620
rect 43474 39564 43484 39620
rect 43540 39564 45388 39620
rect 45444 39564 45454 39620
rect 46396 39564 47180 39620
rect 47236 39564 48188 39620
rect 48244 39564 49532 39620
rect 49588 39564 49598 39620
rect 26852 39508 26908 39564
rect 18610 39452 18620 39508
rect 18676 39452 21756 39508
rect 21812 39452 21822 39508
rect 26852 39452 28588 39508
rect 28644 39452 29372 39508
rect 29428 39452 29438 39508
rect 30370 39452 30380 39508
rect 30436 39452 30828 39508
rect 30884 39452 30894 39508
rect 36306 39452 36316 39508
rect 36372 39452 37324 39508
rect 37380 39452 37390 39508
rect 37548 39452 38892 39508
rect 38948 39452 38958 39508
rect 37548 39396 37604 39452
rect 2930 39340 2940 39396
rect 2996 39340 5740 39396
rect 5796 39340 5806 39396
rect 15474 39340 15484 39396
rect 15540 39340 16716 39396
rect 16772 39340 16782 39396
rect 17490 39340 17500 39396
rect 17556 39340 18228 39396
rect 19058 39340 19068 39396
rect 19124 39340 20188 39396
rect 20244 39340 20972 39396
rect 21028 39340 21038 39396
rect 21522 39340 21532 39396
rect 21588 39340 22652 39396
rect 22708 39340 25676 39396
rect 25732 39340 26348 39396
rect 26404 39340 26414 39396
rect 28466 39340 28476 39396
rect 28532 39340 29484 39396
rect 29540 39340 29550 39396
rect 32274 39340 32284 39396
rect 32340 39340 35644 39396
rect 35700 39340 36428 39396
rect 36484 39340 37604 39396
rect 38322 39340 38332 39396
rect 38388 39340 39228 39396
rect 39284 39340 39294 39396
rect 17574 39228 17612 39284
rect 17668 39228 17678 39284
rect 38994 39228 39004 39284
rect 39060 39228 41020 39284
rect 41076 39228 41086 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 41244 39172 41300 39564
rect 46396 39508 46452 39564
rect 43250 39452 43260 39508
rect 43316 39452 44828 39508
rect 44884 39452 46452 39508
rect 46946 39452 46956 39508
rect 47012 39452 47404 39508
rect 47460 39452 47628 39508
rect 47684 39452 47694 39508
rect 42578 39340 42588 39396
rect 42644 39340 44716 39396
rect 44772 39340 44782 39396
rect 46246 39340 46284 39396
rect 46340 39340 46350 39396
rect 47170 39340 47180 39396
rect 47236 39340 47852 39396
rect 47908 39340 47918 39396
rect 44258 39228 44268 39284
rect 44324 39228 45164 39284
rect 45220 39228 45230 39284
rect 35858 39116 35868 39172
rect 35924 39116 37660 39172
rect 37716 39116 40684 39172
rect 40740 39116 40750 39172
rect 41122 39116 41132 39172
rect 41188 39116 41804 39172
rect 41860 39116 46620 39172
rect 46676 39116 46686 39172
rect 8978 39004 8988 39060
rect 9044 39004 9884 39060
rect 9940 39004 9950 39060
rect 26114 39004 26124 39060
rect 26180 39004 26908 39060
rect 26964 39004 27356 39060
rect 27412 39004 27422 39060
rect 30034 39004 30044 39060
rect 30100 39004 32172 39060
rect 32228 39004 32238 39060
rect 37538 39004 37548 39060
rect 37604 39004 38332 39060
rect 38388 39004 43372 39060
rect 43428 39004 43438 39060
rect 46274 39004 46284 39060
rect 46340 39004 47404 39060
rect 47460 39004 47470 39060
rect 5954 38892 5964 38948
rect 6020 38892 7084 38948
rect 7140 38892 7150 38948
rect 23762 38892 23772 38948
rect 23828 38892 25788 38948
rect 25844 38892 29820 38948
rect 29876 38892 29886 38948
rect 35410 38892 35420 38948
rect 35476 38892 39228 38948
rect 39284 38892 39294 38948
rect 40002 38892 40012 38948
rect 40068 38892 45948 38948
rect 46004 38892 46014 38948
rect 46610 38892 46620 38948
rect 46676 38892 48748 38948
rect 48804 38892 48814 38948
rect 40012 38836 40068 38892
rect 6962 38780 6972 38836
rect 7028 38780 9548 38836
rect 9604 38780 9614 38836
rect 23314 38780 23324 38836
rect 23380 38780 23884 38836
rect 23940 38780 23950 38836
rect 24434 38780 24444 38836
rect 24500 38780 25340 38836
rect 25396 38780 25406 38836
rect 26786 38780 26796 38836
rect 26852 38780 28140 38836
rect 28196 38780 32956 38836
rect 33012 38780 33852 38836
rect 33908 38780 33918 38836
rect 38882 38780 38892 38836
rect 38948 38780 40068 38836
rect 44146 38780 44156 38836
rect 44212 38780 47068 38836
rect 47124 38780 48076 38836
rect 48132 38780 48142 38836
rect 24444 38724 24500 38780
rect 2930 38668 2940 38724
rect 2996 38668 5292 38724
rect 5348 38668 5358 38724
rect 13906 38668 13916 38724
rect 13972 38668 15708 38724
rect 15764 38668 15774 38724
rect 23996 38668 24500 38724
rect 25340 38724 25396 38780
rect 25340 38668 27692 38724
rect 27748 38668 27758 38724
rect 27916 38668 34300 38724
rect 34356 38668 35252 38724
rect 23996 38612 24052 38668
rect 27916 38612 27972 38668
rect 35196 38612 35252 38668
rect 36092 38668 36764 38724
rect 36820 38668 36830 38724
rect 39106 38668 39116 38724
rect 39172 38668 40236 38724
rect 40292 38668 40302 38724
rect 40460 38668 42028 38724
rect 42084 38668 42094 38724
rect 42690 38668 42700 38724
rect 42756 38668 45724 38724
rect 45780 38668 45790 38724
rect 48178 38668 48188 38724
rect 48244 38668 49196 38724
rect 49252 38668 49262 38724
rect 8754 38556 8764 38612
rect 8820 38556 9996 38612
rect 10052 38556 10062 38612
rect 15474 38556 15484 38612
rect 15540 38556 15932 38612
rect 15988 38556 15998 38612
rect 20290 38556 20300 38612
rect 20356 38556 20524 38612
rect 20580 38556 20590 38612
rect 23986 38556 23996 38612
rect 24052 38556 24062 38612
rect 27122 38556 27132 38612
rect 27188 38556 27972 38612
rect 30594 38556 30604 38612
rect 30660 38556 31724 38612
rect 31780 38556 31790 38612
rect 33170 38556 33180 38612
rect 33236 38556 33852 38612
rect 33908 38556 33918 38612
rect 35196 38556 35812 38612
rect 35756 38500 35812 38556
rect 36092 38500 36148 38668
rect 40460 38612 40516 38668
rect 38882 38556 38892 38612
rect 38948 38556 40516 38612
rect 44594 38556 44604 38612
rect 44660 38556 45164 38612
rect 45220 38556 45230 38612
rect 25554 38444 25564 38500
rect 25620 38444 26908 38500
rect 35746 38444 35756 38500
rect 35812 38444 35822 38500
rect 36082 38444 36092 38500
rect 36148 38444 36158 38500
rect 36418 38444 36428 38500
rect 36484 38444 37884 38500
rect 37940 38444 40348 38500
rect 40404 38444 40414 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 26852 38276 26908 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 37622 38332 37660 38388
rect 37716 38332 37726 38388
rect 12674 38220 12684 38276
rect 12740 38220 13580 38276
rect 13636 38220 13646 38276
rect 26852 38220 28812 38276
rect 28868 38220 29596 38276
rect 29652 38220 36876 38276
rect 36932 38220 36942 38276
rect 18162 38108 18172 38164
rect 18228 38108 18732 38164
rect 18788 38108 18798 38164
rect 20962 38108 20972 38164
rect 21028 38108 21644 38164
rect 21700 38108 22764 38164
rect 22820 38108 22830 38164
rect 28578 38108 28588 38164
rect 28644 38108 30212 38164
rect 34850 38108 34860 38164
rect 34916 38108 35196 38164
rect 35252 38108 35262 38164
rect 35522 38108 35532 38164
rect 35588 38108 36988 38164
rect 37044 38108 37054 38164
rect 42242 38108 42252 38164
rect 42308 38108 44156 38164
rect 44212 38108 44222 38164
rect 30156 38052 30212 38108
rect 2706 37996 2716 38052
rect 2772 37996 5628 38052
rect 5684 37996 10556 38052
rect 10612 37996 10622 38052
rect 15138 37996 15148 38052
rect 15204 37996 15596 38052
rect 15652 37996 15932 38052
rect 15988 37996 16380 38052
rect 16436 37996 16940 38052
rect 16996 37996 17006 38052
rect 17154 37996 17164 38052
rect 17220 37996 17724 38052
rect 17780 37996 18284 38052
rect 18340 37996 18350 38052
rect 21858 37996 21868 38052
rect 21924 37996 22428 38052
rect 22484 37996 22494 38052
rect 28466 37996 28476 38052
rect 28532 37996 29372 38052
rect 29428 37996 29438 38052
rect 30146 37996 30156 38052
rect 30212 37996 30604 38052
rect 30660 37996 30670 38052
rect 33954 37996 33964 38052
rect 34020 37996 36204 38052
rect 36260 37996 36270 38052
rect 40226 37996 40236 38052
rect 40292 37996 43708 38052
rect 43764 37996 44380 38052
rect 44436 37996 44828 38052
rect 44884 37996 44894 38052
rect 20066 37884 20076 37940
rect 20132 37884 22540 37940
rect 22596 37884 22606 37940
rect 24658 37884 24668 37940
rect 24724 37884 25452 37940
rect 25508 37884 25518 37940
rect 28242 37884 28252 37940
rect 28308 37884 32284 37940
rect 32340 37884 32350 37940
rect 32722 37884 32732 37940
rect 32788 37884 34860 37940
rect 34916 37884 34926 37940
rect 35746 37884 35756 37940
rect 35812 37884 38892 37940
rect 38948 37884 38958 37940
rect 41010 37884 41020 37940
rect 41076 37884 41580 37940
rect 41636 37884 41646 37940
rect 10770 37772 10780 37828
rect 10836 37772 11788 37828
rect 11844 37772 11854 37828
rect 15026 37772 15036 37828
rect 15092 37772 16156 37828
rect 16212 37772 16222 37828
rect 17266 37772 17276 37828
rect 17332 37772 17948 37828
rect 18004 37772 18508 37828
rect 18564 37772 18574 37828
rect 21746 37772 21756 37828
rect 21812 37772 22204 37828
rect 22260 37772 22270 37828
rect 27682 37772 27692 37828
rect 27748 37772 27916 37828
rect 27972 37772 29372 37828
rect 29428 37772 29438 37828
rect 30482 37772 30492 37828
rect 30548 37772 30558 37828
rect 32498 37772 32508 37828
rect 32564 37772 35868 37828
rect 35924 37772 35934 37828
rect 41234 37772 41244 37828
rect 41300 37772 42812 37828
rect 42868 37772 42878 37828
rect 15362 37660 15372 37716
rect 15428 37660 15820 37716
rect 15876 37660 17388 37716
rect 17444 37660 17454 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 30492 37492 30548 37772
rect 32050 37660 32060 37716
rect 32116 37660 35980 37716
rect 36036 37660 36046 37716
rect 38882 37660 38892 37716
rect 38948 37660 39900 37716
rect 39956 37660 39966 37716
rect 34934 37548 34972 37604
rect 35028 37548 35038 37604
rect 18946 37436 18956 37492
rect 19012 37436 19628 37492
rect 19684 37436 19694 37492
rect 26338 37436 26348 37492
rect 26404 37436 27132 37492
rect 27188 37436 27198 37492
rect 28242 37436 28252 37492
rect 28308 37436 28318 37492
rect 29810 37436 29820 37492
rect 29876 37436 31052 37492
rect 31108 37436 31118 37492
rect 31714 37436 31724 37492
rect 31780 37436 32396 37492
rect 32452 37436 32462 37492
rect 38994 37436 39004 37492
rect 39060 37436 39676 37492
rect 39732 37436 39742 37492
rect 28252 37380 28308 37436
rect 6402 37324 6412 37380
rect 6468 37324 8540 37380
rect 8596 37324 8606 37380
rect 15586 37324 15596 37380
rect 15652 37324 17388 37380
rect 17444 37324 17454 37380
rect 25666 37324 25676 37380
rect 25732 37324 28308 37380
rect 30370 37324 30380 37380
rect 30436 37324 30716 37380
rect 30772 37324 30782 37380
rect 36866 37324 36876 37380
rect 36932 37324 39564 37380
rect 39620 37324 39630 37380
rect 40898 37324 40908 37380
rect 40964 37324 41916 37380
rect 41972 37324 41982 37380
rect 43474 37324 43484 37380
rect 43540 37324 45164 37380
rect 45220 37324 45500 37380
rect 45556 37324 46844 37380
rect 46900 37324 48748 37380
rect 48804 37324 48814 37380
rect 4946 37212 4956 37268
rect 5012 37212 6076 37268
rect 6132 37212 6142 37268
rect 18274 37212 18284 37268
rect 18340 37212 19292 37268
rect 19348 37212 19358 37268
rect 20514 37212 20524 37268
rect 20580 37212 23100 37268
rect 23156 37212 23166 37268
rect 23314 37212 23324 37268
rect 23380 37212 23884 37268
rect 23940 37212 25228 37268
rect 25284 37212 25294 37268
rect 25890 37212 25900 37268
rect 25956 37212 26796 37268
rect 26852 37212 27356 37268
rect 27412 37212 27422 37268
rect 30146 37212 30156 37268
rect 30212 37212 34076 37268
rect 34132 37212 34142 37268
rect 38434 37212 38444 37268
rect 38500 37212 40012 37268
rect 40068 37212 40078 37268
rect 45938 37212 45948 37268
rect 46004 37212 49084 37268
rect 49140 37212 49150 37268
rect 14914 37100 14924 37156
rect 14980 37100 16268 37156
rect 16324 37100 16334 37156
rect 24546 37100 24556 37156
rect 24612 37100 25564 37156
rect 25620 37100 25630 37156
rect 29922 37100 29932 37156
rect 29988 37100 30492 37156
rect 30548 37100 30558 37156
rect 32274 37100 32284 37156
rect 32340 37100 34412 37156
rect 34468 37100 34478 37156
rect 39890 37100 39900 37156
rect 39956 37100 40908 37156
rect 40964 37100 40974 37156
rect 6514 36988 6524 37044
rect 6580 36988 8316 37044
rect 8372 36988 8382 37044
rect 20066 36988 20076 37044
rect 20132 36988 21868 37044
rect 21924 36988 21934 37044
rect 27570 36988 27580 37044
rect 27636 36988 31052 37044
rect 31108 36988 31948 37044
rect 32004 36988 33068 37044
rect 33124 36988 33134 37044
rect 42690 36988 42700 37044
rect 42756 36988 44044 37044
rect 44100 36988 44110 37044
rect 47954 36988 47964 37044
rect 48020 36988 48860 37044
rect 48916 36988 49084 37044
rect 49140 36988 49150 37044
rect 33068 36932 33124 36988
rect 22530 36876 22540 36932
rect 22596 36876 23324 36932
rect 23380 36876 24668 36932
rect 24724 36876 26236 36932
rect 26292 36876 26302 36932
rect 30594 36876 30604 36932
rect 30660 36876 31276 36932
rect 31332 36876 31342 36932
rect 33068 36876 33628 36932
rect 33684 36876 33694 36932
rect 43586 36876 43596 36932
rect 43652 36876 45388 36932
rect 45444 36876 46620 36932
rect 46676 36876 46686 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 2258 36652 2268 36708
rect 2324 36652 2828 36708
rect 2884 36652 3388 36708
rect 16818 36652 16828 36708
rect 16884 36652 17612 36708
rect 17668 36652 17678 36708
rect 22194 36652 22204 36708
rect 22260 36652 22876 36708
rect 22932 36652 22942 36708
rect 34962 36652 34972 36708
rect 35028 36652 35644 36708
rect 35700 36652 35710 36708
rect 3332 36596 3388 36652
rect 3332 36540 4620 36596
rect 4676 36540 4686 36596
rect 8082 36540 8092 36596
rect 8148 36540 10220 36596
rect 10276 36540 11228 36596
rect 11284 36540 11294 36596
rect 20514 36540 20524 36596
rect 20580 36540 21980 36596
rect 22036 36540 22316 36596
rect 22372 36540 22382 36596
rect 29474 36540 29484 36596
rect 29540 36540 31276 36596
rect 31332 36540 31342 36596
rect 34066 36540 34076 36596
rect 34132 36540 40908 36596
rect 40964 36540 40974 36596
rect 49186 36540 49196 36596
rect 49252 36540 49532 36596
rect 49588 36540 49598 36596
rect 9202 36428 9212 36484
rect 9268 36428 9884 36484
rect 9940 36428 9950 36484
rect 10546 36428 10556 36484
rect 10612 36428 11564 36484
rect 11620 36428 11630 36484
rect 30342 36428 30380 36484
rect 30436 36428 30446 36484
rect 33282 36428 33292 36484
rect 33348 36428 35980 36484
rect 36036 36428 36652 36484
rect 36708 36428 36718 36484
rect 41468 36428 42476 36484
rect 42532 36428 42812 36484
rect 42868 36428 42878 36484
rect 45266 36428 45276 36484
rect 45332 36428 45612 36484
rect 45668 36428 48412 36484
rect 48468 36428 48478 36484
rect 10556 36372 10612 36428
rect 41468 36372 41524 36428
rect 8866 36316 8876 36372
rect 8932 36316 9660 36372
rect 9716 36316 10612 36372
rect 12674 36316 12684 36372
rect 12740 36316 13804 36372
rect 13860 36316 13870 36372
rect 32498 36316 32508 36372
rect 32564 36316 34300 36372
rect 34356 36316 34366 36372
rect 37314 36316 37324 36372
rect 37380 36316 41524 36372
rect 41682 36316 41692 36372
rect 41748 36316 41758 36372
rect 41692 36260 41748 36316
rect 9202 36204 9212 36260
rect 9268 36204 11452 36260
rect 11508 36204 11518 36260
rect 13682 36204 13692 36260
rect 13748 36204 15596 36260
rect 15652 36204 15662 36260
rect 19506 36204 19516 36260
rect 19572 36204 21644 36260
rect 21700 36204 21710 36260
rect 22642 36204 22652 36260
rect 22708 36204 24108 36260
rect 24164 36204 24174 36260
rect 24546 36204 24556 36260
rect 24612 36204 32620 36260
rect 32676 36204 32686 36260
rect 37874 36204 37884 36260
rect 37940 36204 41748 36260
rect 43138 36204 43148 36260
rect 43204 36204 45164 36260
rect 45220 36204 47628 36260
rect 47684 36204 49140 36260
rect 49084 36148 49140 36204
rect 50200 36148 51000 36176
rect 49074 36092 49084 36148
rect 49140 36092 49150 36148
rect 49298 36092 49308 36148
rect 49364 36092 51000 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50200 36064 51000 36092
rect 22418 35980 22428 36036
rect 22484 35980 24556 36036
rect 24612 35980 24622 36036
rect 40114 35980 40124 36036
rect 40180 35980 42924 36036
rect 42980 35980 42990 36036
rect 14802 35868 14812 35924
rect 14868 35868 16716 35924
rect 16772 35868 16782 35924
rect 22866 35868 22876 35924
rect 22932 35868 23996 35924
rect 24052 35868 24062 35924
rect 37986 35868 37996 35924
rect 38052 35868 40236 35924
rect 40292 35868 40302 35924
rect 45714 35868 45724 35924
rect 45780 35868 48748 35924
rect 48804 35868 48814 35924
rect 14130 35756 14140 35812
rect 14196 35756 15260 35812
rect 15316 35756 15326 35812
rect 22082 35756 22092 35812
rect 22148 35756 23548 35812
rect 23604 35756 23614 35812
rect 27346 35756 27356 35812
rect 27412 35756 28028 35812
rect 28084 35756 28094 35812
rect 29362 35756 29372 35812
rect 29428 35756 33852 35812
rect 33908 35756 33918 35812
rect 37538 35756 37548 35812
rect 37604 35756 38668 35812
rect 38724 35756 38734 35812
rect 39666 35756 39676 35812
rect 39732 35756 41356 35812
rect 41412 35756 41422 35812
rect 7410 35644 7420 35700
rect 7476 35644 8316 35700
rect 8372 35644 8382 35700
rect 8642 35644 8652 35700
rect 8708 35644 9660 35700
rect 9716 35644 9726 35700
rect 21634 35644 21644 35700
rect 21700 35644 22540 35700
rect 22596 35644 22606 35700
rect 27570 35644 27580 35700
rect 27636 35644 28588 35700
rect 28644 35644 29148 35700
rect 29204 35644 30268 35700
rect 30324 35644 30334 35700
rect 31154 35644 31164 35700
rect 31220 35644 31612 35700
rect 31668 35644 33404 35700
rect 33460 35644 33470 35700
rect 34178 35644 34188 35700
rect 34244 35644 36988 35700
rect 37044 35644 38556 35700
rect 38612 35644 41468 35700
rect 41524 35644 45836 35700
rect 45892 35644 45902 35700
rect 8652 35588 8708 35644
rect 6290 35532 6300 35588
rect 6356 35532 6636 35588
rect 6692 35532 7196 35588
rect 7252 35532 8708 35588
rect 37538 35532 37548 35588
rect 37604 35532 39452 35588
rect 39508 35532 39518 35588
rect 17602 35420 17612 35476
rect 17668 35420 22316 35476
rect 22372 35420 22382 35476
rect 32610 35420 32620 35476
rect 32676 35420 33740 35476
rect 33796 35420 35588 35476
rect 38658 35420 38668 35476
rect 38724 35420 40348 35476
rect 40404 35420 40414 35476
rect 35532 35364 35588 35420
rect 21634 35308 21644 35364
rect 21700 35308 23324 35364
rect 23380 35308 23390 35364
rect 28354 35308 28364 35364
rect 28420 35308 29260 35364
rect 29316 35308 29326 35364
rect 32246 35308 32284 35364
rect 32340 35308 32350 35364
rect 35532 35308 38668 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 38612 35252 38668 35308
rect 1922 35196 1932 35252
rect 1988 35196 3052 35252
rect 3108 35196 3500 35252
rect 3556 35196 3566 35252
rect 8978 35196 8988 35252
rect 9044 35196 10444 35252
rect 10500 35196 11788 35252
rect 11844 35196 12684 35252
rect 12740 35196 12750 35252
rect 18162 35196 18172 35252
rect 18228 35196 18844 35252
rect 18900 35196 18910 35252
rect 21522 35196 21532 35252
rect 21588 35196 23660 35252
rect 23716 35196 23726 35252
rect 29138 35196 29148 35252
rect 29204 35196 29708 35252
rect 29764 35196 29774 35252
rect 38612 35196 39676 35252
rect 39732 35196 39742 35252
rect 40226 35196 40236 35252
rect 40292 35196 40348 35252
rect 40404 35196 40414 35252
rect 44370 35196 44380 35252
rect 44436 35196 47180 35252
rect 47236 35196 47246 35252
rect 21532 35140 21588 35196
rect 2482 35084 2492 35140
rect 2548 35084 3668 35140
rect 7970 35084 7980 35140
rect 8036 35084 9324 35140
rect 9380 35084 9772 35140
rect 9828 35084 9838 35140
rect 17042 35084 17052 35140
rect 17108 35084 18060 35140
rect 18116 35084 21588 35140
rect 27458 35084 27468 35140
rect 27524 35084 28700 35140
rect 28756 35084 28766 35140
rect 29922 35084 29932 35140
rect 29988 35084 30268 35140
rect 30324 35084 30334 35140
rect 32162 35084 32172 35140
rect 32228 35084 32844 35140
rect 32900 35084 35532 35140
rect 35588 35084 35598 35140
rect 37202 35084 37212 35140
rect 37268 35084 38892 35140
rect 38948 35084 38958 35140
rect 39890 35084 39900 35140
rect 39956 35084 43820 35140
rect 43876 35084 45052 35140
rect 45108 35084 45118 35140
rect 3612 35028 3668 35084
rect 3154 34972 3164 35028
rect 3220 34972 3388 35028
rect 3444 34972 3454 35028
rect 3602 34972 3612 35028
rect 3668 34972 3678 35028
rect 5058 34972 5068 35028
rect 5124 34972 6188 35028
rect 6244 34972 6254 35028
rect 7298 34972 7308 35028
rect 7364 34972 8540 35028
rect 8596 34972 8606 35028
rect 13010 34972 13020 35028
rect 13076 34972 14252 35028
rect 14308 34972 14318 35028
rect 17826 34972 17836 35028
rect 17892 34972 20412 35028
rect 20468 34972 21308 35028
rect 21364 34972 21374 35028
rect 31714 34972 31724 35028
rect 31780 34972 32620 35028
rect 32676 34972 32686 35028
rect 37314 34972 37324 35028
rect 37380 34972 39340 35028
rect 39396 34972 39406 35028
rect 43922 34972 43932 35028
rect 43988 34972 48188 35028
rect 48244 34972 48254 35028
rect 3378 34860 3388 34916
rect 3444 34860 5628 34916
rect 5684 34860 5694 34916
rect 16930 34860 16940 34916
rect 16996 34860 18172 34916
rect 18228 34860 20972 34916
rect 21028 34860 22988 34916
rect 23044 34860 23054 34916
rect 29474 34860 29484 34916
rect 29540 34860 30044 34916
rect 30100 34860 30110 34916
rect 40226 34860 40236 34916
rect 40292 34860 41020 34916
rect 41076 34860 41916 34916
rect 41972 34860 41982 34916
rect 45266 34860 45276 34916
rect 45332 34860 47628 34916
rect 47684 34860 47694 34916
rect 2706 34748 2716 34804
rect 2772 34748 3836 34804
rect 3892 34748 5740 34804
rect 5796 34748 5806 34804
rect 38098 34748 38108 34804
rect 38164 34748 39788 34804
rect 39844 34748 39854 34804
rect 44258 34748 44268 34804
rect 44324 34748 44940 34804
rect 44996 34748 45006 34804
rect 46946 34748 46956 34804
rect 47012 34748 48748 34804
rect 48804 34748 48814 34804
rect 2258 34636 2268 34692
rect 2324 34636 2940 34692
rect 2996 34636 3006 34692
rect 3378 34636 3388 34692
rect 3444 34636 3724 34692
rect 3780 34636 3790 34692
rect 4508 34580 4564 34748
rect 4722 34636 4732 34692
rect 4788 34636 5852 34692
rect 5908 34636 5918 34692
rect 9314 34636 9324 34692
rect 9380 34636 10556 34692
rect 10612 34636 10622 34692
rect 42018 34636 42028 34692
rect 42084 34636 47740 34692
rect 47796 34636 48188 34692
rect 48244 34636 48254 34692
rect 4508 34524 4844 34580
rect 4900 34524 4910 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4050 34412 4060 34468
rect 4116 34412 4564 34468
rect 4508 34356 4564 34412
rect 2258 34300 2268 34356
rect 2324 34300 2716 34356
rect 2772 34300 2782 34356
rect 4498 34300 4508 34356
rect 4564 34300 6300 34356
rect 6356 34300 6366 34356
rect 7858 34300 7868 34356
rect 7924 34300 10108 34356
rect 10164 34300 10174 34356
rect 28018 34300 28028 34356
rect 28084 34300 28588 34356
rect 28644 34300 28654 34356
rect 29250 34300 29260 34356
rect 29316 34300 29326 34356
rect 29474 34300 29484 34356
rect 29540 34300 29820 34356
rect 29876 34300 30156 34356
rect 30212 34300 30222 34356
rect 30454 34300 30492 34356
rect 30548 34300 30558 34356
rect 41122 34300 41132 34356
rect 41188 34300 43932 34356
rect 43988 34300 44380 34356
rect 44436 34300 44446 34356
rect 47394 34300 47404 34356
rect 47460 34300 48748 34356
rect 48804 34300 48814 34356
rect 29260 34244 29316 34300
rect 17714 34188 17724 34244
rect 17780 34188 20860 34244
rect 20916 34188 21532 34244
rect 21588 34188 23548 34244
rect 23604 34188 25228 34244
rect 25284 34188 25294 34244
rect 29260 34188 30604 34244
rect 30660 34188 30670 34244
rect 37426 34188 37436 34244
rect 37492 34188 40796 34244
rect 40852 34188 42140 34244
rect 42196 34188 42206 34244
rect 44034 34188 44044 34244
rect 44100 34188 48412 34244
rect 48468 34188 48478 34244
rect 29484 34132 29540 34188
rect 2034 34076 2044 34132
rect 2100 34076 3164 34132
rect 3220 34076 3230 34132
rect 15922 34076 15932 34132
rect 15988 34076 16380 34132
rect 16436 34076 17388 34132
rect 17444 34076 17454 34132
rect 27234 34076 27244 34132
rect 27300 34076 27804 34132
rect 27860 34076 28364 34132
rect 28420 34076 28430 34132
rect 29474 34076 29484 34132
rect 29540 34076 29550 34132
rect 29922 34076 29932 34132
rect 29988 34076 30940 34132
rect 30996 34076 31006 34132
rect 31826 34076 31836 34132
rect 31892 34076 33068 34132
rect 33124 34076 33134 34132
rect 43026 34076 43036 34132
rect 43092 34076 43708 34132
rect 43764 34076 43774 34132
rect 44706 34076 44716 34132
rect 44772 34076 45164 34132
rect 45220 34076 46508 34132
rect 46564 34076 46574 34132
rect 11218 33964 11228 34020
rect 11284 33964 12124 34020
rect 12180 33964 12684 34020
rect 12740 33964 12750 34020
rect 18610 33964 18620 34020
rect 18676 33964 20412 34020
rect 20468 33964 20478 34020
rect 33954 33964 33964 34020
rect 34020 33964 36988 34020
rect 37044 33964 37054 34020
rect 45602 33964 45612 34020
rect 45668 33964 46172 34020
rect 46228 33964 46238 34020
rect 47618 33964 47628 34020
rect 47684 33964 48860 34020
rect 48916 33964 48926 34020
rect 2930 33852 2940 33908
rect 2996 33852 4284 33908
rect 4340 33852 4350 33908
rect 39554 33852 39564 33908
rect 39620 33852 43708 33908
rect 43764 33852 43774 33908
rect 45154 33852 45164 33908
rect 45220 33852 46508 33908
rect 46564 33852 47068 33908
rect 47124 33852 47134 33908
rect 42130 33740 42140 33796
rect 42196 33740 44044 33796
rect 44100 33740 44110 33796
rect 45042 33740 45052 33796
rect 45108 33740 45500 33796
rect 45556 33740 45566 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 43596 33628 45276 33684
rect 45332 33628 45342 33684
rect 43596 33572 43652 33628
rect 17154 33516 17164 33572
rect 17220 33516 17836 33572
rect 17892 33516 17902 33572
rect 23426 33516 23436 33572
rect 23492 33516 24332 33572
rect 24388 33516 24398 33572
rect 27570 33516 27580 33572
rect 27636 33516 32060 33572
rect 32116 33516 35084 33572
rect 35140 33516 35150 33572
rect 41010 33516 41020 33572
rect 41076 33516 41468 33572
rect 41524 33516 43372 33572
rect 43428 33516 43652 33572
rect 5058 33404 5068 33460
rect 5124 33404 5964 33460
rect 6020 33404 6030 33460
rect 19394 33404 19404 33460
rect 19460 33404 20188 33460
rect 20244 33404 20254 33460
rect 29698 33404 29708 33460
rect 29764 33404 30156 33460
rect 30212 33404 30222 33460
rect 34738 33404 34748 33460
rect 34804 33404 36428 33460
rect 36484 33404 36494 33460
rect 39890 33404 39900 33460
rect 39956 33404 40460 33460
rect 40516 33404 40526 33460
rect 41234 33404 41244 33460
rect 41300 33404 42588 33460
rect 42644 33404 42654 33460
rect 45826 33404 45836 33460
rect 45892 33404 47068 33460
rect 47124 33404 47134 33460
rect 9090 33292 9100 33348
rect 9156 33292 11004 33348
rect 11060 33292 11070 33348
rect 12562 33292 12572 33348
rect 12628 33292 13132 33348
rect 13188 33292 13468 33348
rect 13524 33292 13534 33348
rect 17490 33292 17500 33348
rect 17556 33292 18172 33348
rect 18228 33292 19348 33348
rect 28578 33292 28588 33348
rect 28644 33292 29260 33348
rect 29316 33292 29596 33348
rect 29652 33292 29662 33348
rect 32386 33292 32396 33348
rect 32452 33292 33516 33348
rect 33572 33292 33582 33348
rect 19292 33236 19348 33292
rect 7298 33180 7308 33236
rect 7364 33180 7374 33236
rect 7746 33180 7756 33236
rect 7812 33180 8316 33236
rect 8372 33180 8382 33236
rect 9426 33180 9436 33236
rect 9492 33180 10556 33236
rect 10612 33180 10622 33236
rect 13794 33180 13804 33236
rect 13860 33180 15708 33236
rect 15764 33180 15774 33236
rect 16146 33180 16156 33236
rect 16212 33180 17612 33236
rect 17668 33180 17678 33236
rect 19282 33180 19292 33236
rect 19348 33180 19358 33236
rect 33282 33180 33292 33236
rect 33348 33180 34300 33236
rect 34356 33180 34366 33236
rect 37762 33180 37772 33236
rect 37828 33180 40908 33236
rect 40964 33180 40974 33236
rect 42466 33180 42476 33236
rect 42532 33180 45164 33236
rect 45220 33180 45230 33236
rect 7308 33124 7364 33180
rect 7308 33068 8876 33124
rect 8932 33068 10892 33124
rect 10948 33068 11564 33124
rect 11620 33068 11630 33124
rect 15362 33068 15372 33124
rect 15428 33068 17388 33124
rect 17444 33068 17724 33124
rect 17780 33068 18060 33124
rect 18116 33068 18126 33124
rect 18274 33068 18284 33124
rect 18340 33068 19068 33124
rect 19124 33068 19134 33124
rect 19404 33068 20412 33124
rect 20468 33068 20478 33124
rect 25666 33068 25676 33124
rect 25732 33068 26796 33124
rect 26852 33068 26862 33124
rect 31126 33068 31164 33124
rect 31220 33068 31836 33124
rect 31892 33068 31902 33124
rect 7308 33012 7364 33068
rect 19404 33012 19460 33068
rect 44940 33012 44996 33180
rect 6962 32956 6972 33012
rect 7028 32956 7364 33012
rect 14578 32956 14588 33012
rect 14644 32956 16380 33012
rect 16436 32956 16446 33012
rect 19394 32956 19404 33012
rect 19460 32956 19470 33012
rect 30706 32956 30716 33012
rect 30772 32956 32284 33012
rect 32340 32956 32350 33012
rect 37986 32956 37996 33012
rect 38052 32956 39228 33012
rect 39284 32956 39294 33012
rect 44930 32956 44940 33012
rect 44996 32956 45006 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 48038 32844 48076 32900
rect 48132 32844 48142 32900
rect 15698 32732 15708 32788
rect 15764 32732 18508 32788
rect 18564 32732 18574 32788
rect 18722 32732 18732 32788
rect 18788 32732 19068 32788
rect 19124 32732 19134 32788
rect 19506 32732 19516 32788
rect 19572 32732 20076 32788
rect 20132 32732 20142 32788
rect 27906 32732 27916 32788
rect 27972 32732 28700 32788
rect 28756 32732 28766 32788
rect 32274 32732 32284 32788
rect 32340 32732 33180 32788
rect 33236 32732 34300 32788
rect 34356 32732 34366 32788
rect 44930 32732 44940 32788
rect 44996 32732 48020 32788
rect 47964 32676 48020 32732
rect 10098 32620 10108 32676
rect 10164 32620 10780 32676
rect 10836 32620 11228 32676
rect 11284 32620 11294 32676
rect 18610 32620 18620 32676
rect 18676 32620 18956 32676
rect 19012 32620 20412 32676
rect 20468 32620 20478 32676
rect 26898 32620 26908 32676
rect 26964 32620 28364 32676
rect 28420 32620 28430 32676
rect 28914 32620 28924 32676
rect 28980 32620 29708 32676
rect 29764 32620 29774 32676
rect 47964 32620 48076 32676
rect 48132 32620 48748 32676
rect 48804 32620 48814 32676
rect 9762 32508 9772 32564
rect 9828 32508 11116 32564
rect 11172 32508 11676 32564
rect 11732 32508 11742 32564
rect 16594 32508 16604 32564
rect 16660 32508 17276 32564
rect 17332 32508 17342 32564
rect 18834 32508 18844 32564
rect 18900 32508 19516 32564
rect 19572 32508 20300 32564
rect 20356 32508 20366 32564
rect 27122 32508 27132 32564
rect 27188 32508 31500 32564
rect 31556 32508 37548 32564
rect 37604 32508 37614 32564
rect 37986 32508 37996 32564
rect 38052 32508 38556 32564
rect 38612 32508 38892 32564
rect 38948 32508 38958 32564
rect 42802 32508 42812 32564
rect 42868 32508 43484 32564
rect 43540 32508 44716 32564
rect 44772 32508 45388 32564
rect 45444 32508 46452 32564
rect 46610 32508 46620 32564
rect 46676 32508 47628 32564
rect 47684 32508 48412 32564
rect 48468 32508 48478 32564
rect 46396 32452 46452 32508
rect 1922 32396 1932 32452
rect 1988 32396 3052 32452
rect 3108 32396 3118 32452
rect 16818 32396 16828 32452
rect 16884 32396 20860 32452
rect 20916 32396 20926 32452
rect 33170 32396 33180 32452
rect 33236 32396 34412 32452
rect 34468 32396 34478 32452
rect 36194 32396 36204 32452
rect 36260 32396 36988 32452
rect 37044 32396 37054 32452
rect 38434 32396 38444 32452
rect 38500 32396 41020 32452
rect 41076 32396 41086 32452
rect 44370 32396 44380 32452
rect 44436 32396 45724 32452
rect 45780 32396 45790 32452
rect 46396 32396 47852 32452
rect 47908 32396 47918 32452
rect 48066 32396 48076 32452
rect 48132 32396 48524 32452
rect 48580 32396 48590 32452
rect 28466 32284 28476 32340
rect 28532 32284 29260 32340
rect 29316 32284 29326 32340
rect 44258 32284 44268 32340
rect 44324 32284 45052 32340
rect 45108 32284 49084 32340
rect 49140 32284 49150 32340
rect 17602 32172 17612 32228
rect 17668 32172 18060 32228
rect 18116 32172 18126 32228
rect 40450 32172 40460 32228
rect 40516 32172 40908 32228
rect 40964 32172 40974 32228
rect 45462 32172 45500 32228
rect 45556 32172 45566 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 17266 32060 17276 32116
rect 17332 32060 18172 32116
rect 18228 32060 18238 32116
rect 23874 32060 23884 32116
rect 23940 32060 31164 32116
rect 31220 32060 31230 32116
rect 33618 32060 33628 32116
rect 33684 32060 34076 32116
rect 34132 32060 34142 32116
rect 1810 31948 1820 32004
rect 1876 31948 2156 32004
rect 2212 31948 5516 32004
rect 5572 31948 5964 32004
rect 6020 31948 6030 32004
rect 8754 31948 8764 32004
rect 8820 31948 9884 32004
rect 9940 31948 9950 32004
rect 17826 31948 17836 32004
rect 17892 31948 18396 32004
rect 18452 31948 18462 32004
rect 21186 31948 21196 32004
rect 21252 31948 21924 32004
rect 27458 31948 27468 32004
rect 27524 31948 28028 32004
rect 28084 31948 28094 32004
rect 45714 31948 45724 32004
rect 45780 31948 46284 32004
rect 46340 31948 46350 32004
rect 2258 31836 2268 31892
rect 2324 31836 4620 31892
rect 4676 31836 4956 31892
rect 5012 31836 5628 31892
rect 5684 31836 5694 31892
rect 9762 31836 9772 31892
rect 9828 31836 10780 31892
rect 10836 31836 10846 31892
rect 16818 31836 16828 31892
rect 16884 31836 17500 31892
rect 17556 31836 19180 31892
rect 19236 31836 19246 31892
rect 21868 31780 21924 31948
rect 50200 31892 51000 31920
rect 25778 31836 25788 31892
rect 25844 31836 28476 31892
rect 28532 31836 28542 31892
rect 31602 31836 31612 31892
rect 31668 31836 31948 31892
rect 32004 31836 32014 31892
rect 33730 31836 33740 31892
rect 33796 31836 35868 31892
rect 35924 31836 35934 31892
rect 43138 31836 43148 31892
rect 43204 31836 44772 31892
rect 44930 31836 44940 31892
rect 44996 31836 46732 31892
rect 46788 31836 46798 31892
rect 47730 31836 47740 31892
rect 47796 31836 47806 31892
rect 48290 31836 48300 31892
rect 48356 31836 49196 31892
rect 49252 31836 49262 31892
rect 49420 31836 51000 31892
rect 44716 31780 44772 31836
rect 47740 31780 47796 31836
rect 49420 31780 49476 31836
rect 50200 31808 51000 31836
rect 9202 31724 9212 31780
rect 9268 31724 12572 31780
rect 12628 31724 13580 31780
rect 13636 31724 18172 31780
rect 18228 31724 18238 31780
rect 19394 31724 19404 31780
rect 19460 31724 20412 31780
rect 20468 31724 20478 31780
rect 21858 31724 21868 31780
rect 21924 31724 31388 31780
rect 31444 31724 31454 31780
rect 35970 31724 35980 31780
rect 36036 31724 38108 31780
rect 38164 31724 38174 31780
rect 41682 31724 41692 31780
rect 41748 31724 42588 31780
rect 42644 31724 44268 31780
rect 44324 31724 44334 31780
rect 44716 31724 45836 31780
rect 45892 31724 45902 31780
rect 46498 31724 46508 31780
rect 46564 31724 47516 31780
rect 47572 31724 47582 31780
rect 47740 31724 49476 31780
rect 9314 31612 9324 31668
rect 9380 31612 9996 31668
rect 10052 31612 10062 31668
rect 19842 31612 19852 31668
rect 19908 31612 20524 31668
rect 20580 31612 20590 31668
rect 27906 31612 27916 31668
rect 27972 31612 29372 31668
rect 29428 31612 29438 31668
rect 30034 31612 30044 31668
rect 30100 31612 30716 31668
rect 30772 31612 30782 31668
rect 31490 31612 31500 31668
rect 31556 31612 31836 31668
rect 31892 31612 32620 31668
rect 32676 31612 32686 31668
rect 37314 31612 37324 31668
rect 37380 31612 38892 31668
rect 38948 31612 39340 31668
rect 39396 31612 39406 31668
rect 42242 31612 42252 31668
rect 42308 31612 43820 31668
rect 43876 31612 43886 31668
rect 45602 31612 45612 31668
rect 45668 31612 46620 31668
rect 46676 31612 46686 31668
rect 18946 31500 18956 31556
rect 19012 31500 19628 31556
rect 19684 31500 20748 31556
rect 20804 31500 20814 31556
rect 29810 31500 29820 31556
rect 29876 31500 30940 31556
rect 30996 31500 31006 31556
rect 36306 31500 36316 31556
rect 36372 31500 37436 31556
rect 37492 31500 37502 31556
rect 38322 31500 38332 31556
rect 38388 31500 39396 31556
rect 39666 31500 39676 31556
rect 39732 31500 40796 31556
rect 40852 31500 40862 31556
rect 41346 31500 41356 31556
rect 41412 31500 42364 31556
rect 42420 31500 42430 31556
rect 43026 31500 43036 31556
rect 43092 31500 46508 31556
rect 46564 31500 46574 31556
rect 18274 31388 18284 31444
rect 18340 31388 19180 31444
rect 19236 31388 19246 31444
rect 20178 31388 20188 31444
rect 20244 31388 20636 31444
rect 20692 31388 21140 31444
rect 21522 31388 21532 31444
rect 21588 31388 23884 31444
rect 23940 31388 23950 31444
rect 34178 31388 34188 31444
rect 34244 31388 34748 31444
rect 34804 31388 36092 31444
rect 36148 31388 38220 31444
rect 38276 31388 38286 31444
rect 38612 31388 39116 31444
rect 39172 31388 39182 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 21084 31332 21140 31388
rect 20514 31276 20524 31332
rect 20580 31276 20590 31332
rect 21084 31276 29596 31332
rect 29652 31276 30940 31332
rect 30996 31276 31164 31332
rect 31220 31276 31230 31332
rect 33814 31276 33852 31332
rect 33908 31276 33918 31332
rect 34066 31276 34076 31332
rect 34132 31276 34524 31332
rect 34580 31276 35084 31332
rect 35140 31276 35756 31332
rect 35812 31276 38444 31332
rect 38500 31276 38510 31332
rect 20524 31220 20580 31276
rect 38612 31220 38668 31388
rect 39340 31332 39396 31500
rect 41458 31388 41468 31444
rect 41524 31388 42924 31444
rect 42980 31388 46844 31444
rect 46900 31388 46910 31444
rect 38882 31276 38892 31332
rect 38948 31276 41692 31332
rect 41748 31276 41758 31332
rect 8306 31164 8316 31220
rect 8372 31164 9548 31220
rect 9604 31164 10668 31220
rect 10724 31164 10734 31220
rect 16706 31164 16716 31220
rect 16772 31164 17388 31220
rect 17444 31164 18508 31220
rect 18564 31164 18574 31220
rect 20524 31164 21532 31220
rect 21588 31164 21598 31220
rect 26114 31164 26124 31220
rect 26180 31164 38668 31220
rect 44594 31164 44604 31220
rect 44660 31164 45612 31220
rect 45668 31164 45678 31220
rect 6290 31052 6300 31108
rect 6356 31052 8204 31108
rect 8260 31052 8270 31108
rect 8642 31052 8652 31108
rect 8708 31052 9212 31108
rect 9268 31052 10444 31108
rect 10500 31052 10510 31108
rect 17714 31052 17724 31108
rect 17780 31052 18284 31108
rect 18340 31052 18350 31108
rect 20290 31052 20300 31108
rect 20356 31052 21308 31108
rect 21364 31052 21374 31108
rect 30482 31052 30492 31108
rect 30548 31052 31948 31108
rect 32004 31052 32014 31108
rect 34402 31052 34412 31108
rect 34468 31052 36652 31108
rect 36708 31052 37212 31108
rect 37268 31052 37278 31108
rect 38658 31052 38668 31108
rect 38724 31052 39004 31108
rect 39060 31052 39070 31108
rect 44930 31052 44940 31108
rect 44996 31052 47684 31108
rect 47628 30996 47684 31052
rect 2594 30940 2604 30996
rect 2660 30940 3500 30996
rect 3556 30940 4060 30996
rect 4116 30940 4126 30996
rect 12114 30940 12124 30996
rect 12180 30940 13020 30996
rect 13076 30940 13086 30996
rect 13804 30940 16044 30996
rect 16100 30940 16110 30996
rect 21410 30940 21420 30996
rect 21476 30940 24556 30996
rect 24612 30940 24622 30996
rect 31714 30940 31724 30996
rect 31780 30940 32060 30996
rect 32116 30940 33180 30996
rect 33236 30940 33246 30996
rect 34178 30940 34188 30996
rect 34244 30940 34524 30996
rect 34580 30940 35308 30996
rect 35364 30940 35374 30996
rect 43474 30940 43484 30996
rect 43540 30940 43932 30996
rect 43988 30940 43998 30996
rect 46050 30940 46060 30996
rect 46116 30940 47292 30996
rect 47348 30940 47358 30996
rect 47618 30940 47628 30996
rect 47684 30940 49308 30996
rect 49364 30940 49374 30996
rect 6850 30828 6860 30884
rect 6916 30828 7532 30884
rect 7588 30828 7598 30884
rect 13804 30772 13860 30940
rect 43932 30884 43988 30940
rect 18834 30828 18844 30884
rect 18900 30828 19628 30884
rect 19684 30828 22764 30884
rect 22820 30828 22830 30884
rect 29138 30828 29148 30884
rect 29204 30828 31948 30884
rect 32004 30828 40460 30884
rect 40516 30828 42700 30884
rect 42756 30828 42766 30884
rect 43932 30828 46284 30884
rect 46340 30828 46350 30884
rect 5954 30716 5964 30772
rect 6020 30716 6412 30772
rect 6468 30716 7196 30772
rect 7252 30716 7262 30772
rect 13794 30716 13804 30772
rect 13860 30716 13870 30772
rect 16258 30716 16268 30772
rect 16324 30716 17724 30772
rect 17780 30716 18620 30772
rect 18676 30716 18686 30772
rect 28690 30716 28700 30772
rect 28756 30716 29932 30772
rect 29988 30716 29998 30772
rect 34402 30716 34412 30772
rect 34468 30716 35196 30772
rect 35252 30716 35262 30772
rect 45266 30716 45276 30772
rect 45332 30716 46844 30772
rect 46900 30716 46910 30772
rect 48066 30604 48076 30660
rect 48132 30604 48524 30660
rect 48580 30604 48590 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 7186 30492 7196 30548
rect 7252 30492 8316 30548
rect 8372 30492 8382 30548
rect 10210 30492 10220 30548
rect 10276 30492 14476 30548
rect 14532 30492 14542 30548
rect 36530 30492 36540 30548
rect 36596 30492 37548 30548
rect 37604 30492 37614 30548
rect 45042 30492 45052 30548
rect 45108 30492 46508 30548
rect 46564 30492 48636 30548
rect 48692 30492 48702 30548
rect 36540 30436 36596 30492
rect 3042 30380 3052 30436
rect 3108 30380 7868 30436
rect 7924 30380 7934 30436
rect 23426 30380 23436 30436
rect 23492 30380 27692 30436
rect 27748 30380 28140 30436
rect 28196 30380 28206 30436
rect 33842 30380 33852 30436
rect 33908 30380 36596 30436
rect 42588 30380 43260 30436
rect 43316 30380 43326 30436
rect 46386 30380 46396 30436
rect 46452 30380 47404 30436
rect 47460 30380 47470 30436
rect 47954 30380 47964 30436
rect 48020 30380 48860 30436
rect 48916 30380 49532 30436
rect 49588 30380 49598 30436
rect 8306 30268 8316 30324
rect 8372 30268 9996 30324
rect 10052 30268 10062 30324
rect 13906 30268 13916 30324
rect 13972 30268 17500 30324
rect 17556 30268 17566 30324
rect 26236 30268 27468 30324
rect 27524 30268 27534 30324
rect 30706 30268 30716 30324
rect 30772 30268 31836 30324
rect 31892 30268 31902 30324
rect 38098 30268 38108 30324
rect 38164 30268 39676 30324
rect 39732 30268 39742 30324
rect 40562 30268 40572 30324
rect 40628 30268 40638 30324
rect 41458 30268 41468 30324
rect 41524 30268 41916 30324
rect 41972 30268 41982 30324
rect 26236 30212 26292 30268
rect 40572 30212 40628 30268
rect 42588 30212 42644 30380
rect 42812 30268 45164 30324
rect 45220 30268 45230 30324
rect 46610 30268 46620 30324
rect 46676 30268 47516 30324
rect 47572 30268 47582 30324
rect 47730 30268 47740 30324
rect 47796 30268 48748 30324
rect 48804 30268 48814 30324
rect 23202 30156 23212 30212
rect 23268 30156 24220 30212
rect 24276 30156 24286 30212
rect 26226 30156 26236 30212
rect 26292 30156 26302 30212
rect 27346 30156 27356 30212
rect 27412 30156 30268 30212
rect 30324 30156 30334 30212
rect 31042 30156 31052 30212
rect 31108 30156 31164 30212
rect 31220 30156 31724 30212
rect 31780 30156 31790 30212
rect 33394 30156 33404 30212
rect 33460 30156 35196 30212
rect 35252 30156 35262 30212
rect 35420 30156 37884 30212
rect 37940 30156 38220 30212
rect 38276 30156 38286 30212
rect 40572 30156 41244 30212
rect 41300 30156 41310 30212
rect 42578 30156 42588 30212
rect 42644 30156 42654 30212
rect 4946 30044 4956 30100
rect 5012 30044 5292 30100
rect 5348 30044 5358 30100
rect 18386 30044 18396 30100
rect 18452 30044 23548 30100
rect 23604 30044 24668 30100
rect 24724 30044 24734 30100
rect 26236 29988 26292 30156
rect 35420 30100 35476 30156
rect 28466 30044 28476 30100
rect 28532 30044 30716 30100
rect 30772 30044 30782 30100
rect 31714 30044 31724 30100
rect 31780 30044 35476 30100
rect 36418 30044 36428 30100
rect 36484 30044 39116 30100
rect 39172 30044 39182 30100
rect 40226 30044 40236 30100
rect 40292 30044 40796 30100
rect 40852 30044 40862 30100
rect 42812 29988 42868 30268
rect 44146 30156 44156 30212
rect 44212 30156 46396 30212
rect 46452 30156 47404 30212
rect 47460 30156 47470 30212
rect 48066 30156 48076 30212
rect 48132 30156 48188 30212
rect 48244 30156 48254 30212
rect 43362 30044 43372 30100
rect 43428 30044 46004 30100
rect 46274 30044 46284 30100
rect 46340 30044 49084 30100
rect 49140 30044 49150 30100
rect 45948 29988 46004 30044
rect 15026 29932 15036 29988
rect 15092 29932 15708 29988
rect 15764 29932 15774 29988
rect 20066 29932 20076 29988
rect 20132 29932 21196 29988
rect 21252 29932 21262 29988
rect 22418 29932 22428 29988
rect 22484 29932 24220 29988
rect 24276 29932 24780 29988
rect 24836 29932 25004 29988
rect 25060 29932 26292 29988
rect 26898 29932 26908 29988
rect 26964 29932 28588 29988
rect 28644 29932 28654 29988
rect 29698 29932 29708 29988
rect 29764 29932 30492 29988
rect 30548 29932 30558 29988
rect 30818 29932 30828 29988
rect 30884 29932 33964 29988
rect 34020 29932 34030 29988
rect 37650 29932 37660 29988
rect 37716 29932 38108 29988
rect 38164 29932 38174 29988
rect 42802 29932 42812 29988
rect 42868 29932 42878 29988
rect 43922 29932 43932 29988
rect 43988 29932 45724 29988
rect 45780 29932 45790 29988
rect 45938 29932 45948 29988
rect 46004 29932 46014 29988
rect 46722 29932 46732 29988
rect 46788 29932 47404 29988
rect 47460 29932 47470 29988
rect 29708 29876 29764 29932
rect 21634 29820 21644 29876
rect 21700 29820 22652 29876
rect 22708 29820 23772 29876
rect 23828 29820 23838 29876
rect 27906 29820 27916 29876
rect 27972 29820 29764 29876
rect 33964 29876 34020 29932
rect 33964 29820 41580 29876
rect 41636 29820 41646 29876
rect 42690 29820 42700 29876
rect 42756 29820 43596 29876
rect 43652 29820 43662 29876
rect 45462 29820 45500 29876
rect 45556 29820 45566 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 42700 29764 42756 29820
rect 21410 29708 21420 29764
rect 21476 29708 23884 29764
rect 23940 29708 23950 29764
rect 33282 29708 33292 29764
rect 33348 29708 34860 29764
rect 34916 29708 34926 29764
rect 36978 29708 36988 29764
rect 37044 29708 37660 29764
rect 37716 29708 37726 29764
rect 40114 29708 40124 29764
rect 40180 29708 40460 29764
rect 40516 29708 40526 29764
rect 41122 29708 41132 29764
rect 41188 29708 42756 29764
rect 45602 29708 45612 29764
rect 45668 29708 46844 29764
rect 46900 29708 46910 29764
rect 21420 29652 21476 29708
rect 19394 29596 19404 29652
rect 19460 29596 21476 29652
rect 33058 29596 33068 29652
rect 33124 29596 33516 29652
rect 33572 29596 33582 29652
rect 36418 29596 36428 29652
rect 36484 29596 37996 29652
rect 38052 29596 40348 29652
rect 40404 29596 40414 29652
rect 25554 29484 25564 29540
rect 25620 29484 27132 29540
rect 27188 29484 27692 29540
rect 27748 29484 27758 29540
rect 30258 29484 30268 29540
rect 30324 29484 34860 29540
rect 34916 29484 34926 29540
rect 40002 29484 40012 29540
rect 40068 29484 40908 29540
rect 40964 29484 40974 29540
rect 47058 29484 47068 29540
rect 47124 29484 48860 29540
rect 48916 29484 49084 29540
rect 49140 29484 49150 29540
rect 4610 29372 4620 29428
rect 4676 29372 5516 29428
rect 5572 29372 5582 29428
rect 6626 29372 6636 29428
rect 6692 29372 7308 29428
rect 7364 29372 7980 29428
rect 8036 29372 8046 29428
rect 24658 29372 24668 29428
rect 24724 29372 25228 29428
rect 25284 29372 25294 29428
rect 31378 29372 31388 29428
rect 31444 29372 32172 29428
rect 32228 29372 33068 29428
rect 33124 29372 33134 29428
rect 33506 29372 33516 29428
rect 33572 29372 33740 29428
rect 33796 29372 35196 29428
rect 35252 29372 35262 29428
rect 37986 29372 37996 29428
rect 38052 29372 42924 29428
rect 42980 29372 44716 29428
rect 44772 29372 44782 29428
rect 12114 29260 12124 29316
rect 12180 29260 14476 29316
rect 14532 29260 14542 29316
rect 14690 29260 14700 29316
rect 14756 29260 15484 29316
rect 15540 29260 15550 29316
rect 33842 29260 33852 29316
rect 33908 29260 35756 29316
rect 35812 29260 35822 29316
rect 39788 29260 40236 29316
rect 40292 29260 41468 29316
rect 41524 29260 41534 29316
rect 41906 29260 41916 29316
rect 41972 29260 42812 29316
rect 42868 29260 42878 29316
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 14476 28980 14532 29260
rect 30706 29148 30716 29204
rect 30772 29148 31052 29204
rect 31108 29148 35588 29204
rect 35970 29148 35980 29204
rect 36036 29148 38668 29204
rect 38724 29148 38734 29204
rect 35532 29092 35588 29148
rect 39788 29092 39844 29260
rect 40002 29148 40012 29204
rect 40068 29148 41804 29204
rect 41860 29148 41870 29204
rect 19842 29036 19852 29092
rect 19908 29036 29148 29092
rect 29204 29036 29214 29092
rect 35532 29036 39844 29092
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 14476 28924 21084 28980
rect 21140 28924 21150 28980
rect 41682 28924 41692 28980
rect 41748 28924 42140 28980
rect 42196 28924 42206 28980
rect 4722 28812 4732 28868
rect 4788 28812 5628 28868
rect 5684 28812 5694 28868
rect 22978 28812 22988 28868
rect 23044 28812 25452 28868
rect 25508 28812 25518 28868
rect 26852 28812 30828 28868
rect 30884 28812 31724 28868
rect 31780 28812 31790 28868
rect 34626 28812 34636 28868
rect 34692 28812 41244 28868
rect 41300 28812 43148 28868
rect 43204 28812 43214 28868
rect 43698 28812 43708 28868
rect 43764 28812 47740 28868
rect 47796 28812 47806 28868
rect 26852 28756 26908 28812
rect 43148 28756 43204 28812
rect 3266 28700 3276 28756
rect 3332 28700 4396 28756
rect 4452 28700 4462 28756
rect 6402 28700 6412 28756
rect 6468 28700 6478 28756
rect 14018 28700 14028 28756
rect 14084 28700 14924 28756
rect 14980 28700 21868 28756
rect 21924 28700 23100 28756
rect 23156 28700 23166 28756
rect 26338 28700 26348 28756
rect 26404 28700 26908 28756
rect 29922 28700 29932 28756
rect 29988 28700 33908 28756
rect 35298 28700 35308 28756
rect 35364 28700 35980 28756
rect 36036 28700 36046 28756
rect 38434 28700 38444 28756
rect 38500 28700 40460 28756
rect 40516 28700 40526 28756
rect 40898 28700 40908 28756
rect 40964 28700 41636 28756
rect 43148 28700 44044 28756
rect 44100 28700 45500 28756
rect 45556 28700 45566 28756
rect 6412 28644 6468 28700
rect 2594 28588 2604 28644
rect 2660 28588 3388 28644
rect 3444 28588 3454 28644
rect 3602 28588 3612 28644
rect 3668 28588 4508 28644
rect 4564 28588 5292 28644
rect 5348 28588 5358 28644
rect 5954 28588 5964 28644
rect 6020 28588 6636 28644
rect 6692 28588 8764 28644
rect 8820 28588 8830 28644
rect 16258 28588 16268 28644
rect 16324 28588 17052 28644
rect 17108 28588 17118 28644
rect 19618 28588 19628 28644
rect 19684 28588 20636 28644
rect 20692 28588 21644 28644
rect 21700 28588 21710 28644
rect 22530 28588 22540 28644
rect 22596 28588 23324 28644
rect 23380 28588 23390 28644
rect 25330 28588 25340 28644
rect 25396 28588 27692 28644
rect 27748 28588 27758 28644
rect 28578 28588 28588 28644
rect 28644 28588 31276 28644
rect 31332 28588 31342 28644
rect 7756 28532 7812 28588
rect 33852 28532 33908 28700
rect 41580 28644 41636 28700
rect 34066 28588 34076 28644
rect 34132 28588 35868 28644
rect 35924 28588 35934 28644
rect 39890 28588 39900 28644
rect 39956 28588 41356 28644
rect 41412 28588 41422 28644
rect 41580 28588 43764 28644
rect 44370 28588 44380 28644
rect 44436 28588 46060 28644
rect 46116 28588 46126 28644
rect 47394 28588 47404 28644
rect 47460 28588 48076 28644
rect 48132 28588 48142 28644
rect 43708 28532 43764 28588
rect 3714 28476 3724 28532
rect 3780 28476 4844 28532
rect 4900 28476 4910 28532
rect 7746 28476 7756 28532
rect 7812 28476 7822 28532
rect 17826 28476 17836 28532
rect 17892 28476 19180 28532
rect 19236 28476 19246 28532
rect 21074 28476 21084 28532
rect 21140 28476 22428 28532
rect 22484 28476 22494 28532
rect 28466 28476 28476 28532
rect 28532 28476 29484 28532
rect 29540 28476 29550 28532
rect 33852 28476 35756 28532
rect 35812 28476 35822 28532
rect 37426 28476 37436 28532
rect 37492 28476 38332 28532
rect 38388 28476 40348 28532
rect 40404 28476 40414 28532
rect 42578 28476 42588 28532
rect 42644 28476 43148 28532
rect 43204 28476 43214 28532
rect 43708 28476 45388 28532
rect 45444 28476 45454 28532
rect 7074 28364 7084 28420
rect 7140 28364 8988 28420
rect 9044 28364 9054 28420
rect 17714 28364 17724 28420
rect 17780 28364 19404 28420
rect 19460 28364 19852 28420
rect 19908 28364 19918 28420
rect 26562 28364 26572 28420
rect 26628 28364 27580 28420
rect 27636 28364 27646 28420
rect 27794 28364 27804 28420
rect 27860 28364 28700 28420
rect 28756 28364 29372 28420
rect 29428 28364 29438 28420
rect 16706 28252 16716 28308
rect 16772 28252 18732 28308
rect 18788 28252 18798 28308
rect 22754 28252 22764 28308
rect 22820 28252 24108 28308
rect 24164 28252 24174 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 23202 28140 23212 28196
rect 23268 28140 38108 28196
rect 38164 28140 38174 28196
rect 12338 28028 12348 28084
rect 12404 28028 13468 28084
rect 13524 28028 13534 28084
rect 16370 28028 16380 28084
rect 16436 28028 19348 28084
rect 20738 28028 20748 28084
rect 20804 28028 21196 28084
rect 21252 28028 21262 28084
rect 26898 28028 26908 28084
rect 26964 28028 27916 28084
rect 27972 28028 27982 28084
rect 32274 28028 32284 28084
rect 32340 28028 33180 28084
rect 33236 28028 33246 28084
rect 19292 27972 19348 28028
rect 13794 27916 13804 27972
rect 13860 27916 14700 27972
rect 14756 27916 15260 27972
rect 15316 27916 16604 27972
rect 16660 27916 16670 27972
rect 19282 27916 19292 27972
rect 19348 27916 21756 27972
rect 21812 27916 27356 27972
rect 27412 27916 27422 27972
rect 33618 27916 33628 27972
rect 33684 27916 35644 27972
rect 35700 27916 35710 27972
rect 36194 27916 36204 27972
rect 36260 27916 36988 27972
rect 37044 27916 37054 27972
rect 4610 27804 4620 27860
rect 4676 27804 5516 27860
rect 5572 27804 5582 27860
rect 5842 27804 5852 27860
rect 5908 27804 7420 27860
rect 7476 27804 7486 27860
rect 15026 27804 15036 27860
rect 15092 27804 15932 27860
rect 15988 27804 16156 27860
rect 16212 27804 16222 27860
rect 16482 27804 16492 27860
rect 16548 27804 17388 27860
rect 17444 27804 17454 27860
rect 18162 27804 18172 27860
rect 18228 27804 19628 27860
rect 19684 27804 20300 27860
rect 20356 27804 20366 27860
rect 24770 27804 24780 27860
rect 24836 27804 27468 27860
rect 27524 27804 27534 27860
rect 31154 27804 31164 27860
rect 31220 27804 32340 27860
rect 32498 27804 32508 27860
rect 32564 27804 34412 27860
rect 34468 27804 34478 27860
rect 44706 27804 44716 27860
rect 44772 27804 45836 27860
rect 45892 27804 45902 27860
rect 32284 27748 32340 27804
rect 6514 27692 6524 27748
rect 6580 27692 7868 27748
rect 7924 27692 8988 27748
rect 9044 27692 9054 27748
rect 11442 27692 11452 27748
rect 11508 27692 12012 27748
rect 12068 27692 12078 27748
rect 12786 27692 12796 27748
rect 12852 27692 13132 27748
rect 13188 27692 13692 27748
rect 13748 27692 13758 27748
rect 23874 27692 23884 27748
rect 23940 27692 25228 27748
rect 25284 27692 25294 27748
rect 25442 27692 25452 27748
rect 25508 27692 30716 27748
rect 30772 27692 32060 27748
rect 32116 27692 32126 27748
rect 32274 27692 32284 27748
rect 32340 27692 34132 27748
rect 36194 27692 36204 27748
rect 36260 27692 37996 27748
rect 38052 27692 38668 27748
rect 38724 27692 38734 27748
rect 39330 27692 39340 27748
rect 39396 27692 39900 27748
rect 39956 27692 44156 27748
rect 44212 27692 45052 27748
rect 45108 27692 45118 27748
rect 46610 27692 46620 27748
rect 46676 27692 48972 27748
rect 49028 27692 49038 27748
rect 34076 27636 34132 27692
rect 50200 27636 51000 27664
rect 6066 27580 6076 27636
rect 6132 27580 8540 27636
rect 8596 27580 8606 27636
rect 17938 27580 17948 27636
rect 18004 27580 18396 27636
rect 18452 27580 19852 27636
rect 19908 27580 19918 27636
rect 20066 27580 20076 27636
rect 20132 27580 24892 27636
rect 24948 27580 26348 27636
rect 26404 27580 26414 27636
rect 33170 27580 33180 27636
rect 33236 27580 33852 27636
rect 33908 27580 33918 27636
rect 34076 27580 37548 27636
rect 37604 27580 37614 27636
rect 46470 27580 46508 27636
rect 46564 27580 46574 27636
rect 48402 27580 48412 27636
rect 48468 27580 48748 27636
rect 48804 27580 48814 27636
rect 49186 27580 49196 27636
rect 49252 27580 51000 27636
rect 50200 27552 51000 27580
rect 18274 27468 18284 27524
rect 18340 27468 19180 27524
rect 19236 27468 19246 27524
rect 33842 27468 33852 27524
rect 33908 27468 34076 27524
rect 34132 27468 34142 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 12562 27356 12572 27412
rect 12628 27356 13300 27412
rect 16818 27356 16828 27412
rect 16884 27356 18620 27412
rect 18676 27356 18686 27412
rect 31490 27356 31500 27412
rect 31556 27356 34860 27412
rect 34916 27356 34926 27412
rect 13244 27300 13300 27356
rect 3266 27244 3276 27300
rect 3332 27244 3836 27300
rect 3892 27244 4508 27300
rect 4564 27244 4574 27300
rect 5058 27244 5068 27300
rect 5124 27244 5964 27300
rect 6020 27244 6030 27300
rect 6402 27244 6412 27300
rect 6468 27244 7084 27300
rect 7140 27244 7150 27300
rect 13234 27244 13244 27300
rect 13300 27244 15260 27300
rect 15316 27244 15820 27300
rect 15876 27244 15886 27300
rect 17378 27244 17388 27300
rect 17444 27244 18284 27300
rect 18340 27244 19740 27300
rect 19796 27244 19806 27300
rect 20412 27244 21980 27300
rect 22036 27244 22046 27300
rect 20412 27188 20468 27244
rect 15260 27132 20412 27188
rect 20468 27132 20478 27188
rect 20738 27132 20748 27188
rect 20804 27132 21420 27188
rect 21476 27132 30156 27188
rect 30212 27132 30222 27188
rect 35746 27132 35756 27188
rect 35812 27132 39116 27188
rect 39172 27132 39182 27188
rect 48066 27132 48076 27188
rect 48132 27132 48860 27188
rect 48916 27132 49196 27188
rect 49252 27132 49262 27188
rect 4834 27020 4844 27076
rect 4900 27020 5292 27076
rect 5348 27020 5358 27076
rect 15260 26964 15316 27132
rect 16594 27020 16604 27076
rect 16660 27020 17164 27076
rect 17220 27020 17230 27076
rect 18050 27020 18060 27076
rect 18116 27020 18508 27076
rect 18564 27020 18574 27076
rect 35634 27020 35644 27076
rect 35700 27020 36988 27076
rect 37044 27020 37054 27076
rect 2482 26908 2492 26964
rect 2548 26908 3612 26964
rect 3668 26908 3678 26964
rect 13916 26908 15316 26964
rect 15474 26908 15484 26964
rect 15540 26908 16380 26964
rect 16436 26908 16446 26964
rect 21410 26908 21420 26964
rect 21476 26908 23436 26964
rect 23492 26908 23502 26964
rect 27570 26908 27580 26964
rect 27636 26908 28476 26964
rect 28532 26908 29372 26964
rect 29428 26908 29438 26964
rect 29586 26908 29596 26964
rect 29652 26908 30380 26964
rect 30436 26908 31724 26964
rect 31780 26908 31790 26964
rect 37958 26908 37996 26964
rect 38052 26908 38062 26964
rect 47058 26908 47068 26964
rect 47124 26908 47516 26964
rect 47572 26908 47582 26964
rect 13916 26852 13972 26908
rect 3938 26796 3948 26852
rect 4004 26796 5068 26852
rect 5124 26796 5134 26852
rect 13906 26796 13916 26852
rect 13972 26796 13982 26852
rect 16706 26796 16716 26852
rect 16772 26796 17388 26852
rect 17444 26796 17454 26852
rect 17826 26796 17836 26852
rect 17892 26796 22988 26852
rect 23044 26796 23054 26852
rect 26786 26796 26796 26852
rect 26852 26796 28252 26852
rect 28308 26796 28318 26852
rect 30594 26796 30604 26852
rect 30660 26796 31612 26852
rect 31668 26796 32060 26852
rect 32116 26796 32508 26852
rect 32564 26796 33292 26852
rect 33348 26796 37660 26852
rect 37716 26796 37726 26852
rect 43026 26796 43036 26852
rect 43092 26796 44044 26852
rect 44100 26796 44110 26852
rect 19292 26628 19348 26796
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 19282 26572 19292 26628
rect 19348 26572 19358 26628
rect 16482 26460 16492 26516
rect 16548 26460 17612 26516
rect 17668 26460 17678 26516
rect 20514 26460 20524 26516
rect 20580 26460 20972 26516
rect 21028 26460 23212 26516
rect 23268 26460 23278 26516
rect 28252 26404 28308 26796
rect 42690 26684 42700 26740
rect 42756 26684 43596 26740
rect 43652 26684 43662 26740
rect 30370 26572 30380 26628
rect 30436 26572 30940 26628
rect 30996 26572 31006 26628
rect 38882 26572 38892 26628
rect 38948 26572 40236 26628
rect 40292 26572 47628 26628
rect 47684 26572 48748 26628
rect 48804 26572 48814 26628
rect 30146 26460 30156 26516
rect 30212 26460 30716 26516
rect 30772 26460 30782 26516
rect 42130 26460 42140 26516
rect 42196 26460 42924 26516
rect 42980 26460 42990 26516
rect 45266 26460 45276 26516
rect 45332 26460 46060 26516
rect 46116 26460 46508 26516
rect 46564 26460 47516 26516
rect 47572 26460 47582 26516
rect 13570 26348 13580 26404
rect 13636 26348 14140 26404
rect 14196 26348 14206 26404
rect 14588 26348 15708 26404
rect 15764 26348 17836 26404
rect 17892 26348 17902 26404
rect 28242 26348 28252 26404
rect 28308 26348 28318 26404
rect 30482 26348 30492 26404
rect 30548 26348 33460 26404
rect 40786 26348 40796 26404
rect 40852 26348 46620 26404
rect 46676 26348 46686 26404
rect 46834 26348 46844 26404
rect 46900 26348 47852 26404
rect 47908 26348 47918 26404
rect 14588 26292 14644 26348
rect 33404 26292 33460 26348
rect 1810 26236 1820 26292
rect 1876 26236 6188 26292
rect 6244 26236 8428 26292
rect 8484 26236 9212 26292
rect 9268 26236 9548 26292
rect 9604 26236 9614 26292
rect 12450 26236 12460 26292
rect 12516 26236 13692 26292
rect 13748 26236 14588 26292
rect 14644 26236 14654 26292
rect 15810 26236 15820 26292
rect 15876 26236 16604 26292
rect 16660 26236 17500 26292
rect 17556 26236 17566 26292
rect 25442 26236 25452 26292
rect 25508 26236 28588 26292
rect 28644 26236 28654 26292
rect 28802 26236 28812 26292
rect 28868 26236 32732 26292
rect 32788 26236 32798 26292
rect 33394 26236 33404 26292
rect 33460 26236 34636 26292
rect 34692 26236 34702 26292
rect 44258 26236 44268 26292
rect 44324 26236 45724 26292
rect 45780 26236 45790 26292
rect 47058 26236 47068 26292
rect 47124 26236 48188 26292
rect 48244 26236 48254 26292
rect 21298 26124 21308 26180
rect 21364 26124 22092 26180
rect 22148 26124 22158 26180
rect 23090 26124 23100 26180
rect 23156 26124 23884 26180
rect 23940 26124 23950 26180
rect 25778 26124 25788 26180
rect 25844 26124 30492 26180
rect 30548 26124 31052 26180
rect 31108 26124 31118 26180
rect 33058 26124 33068 26180
rect 33124 26124 33852 26180
rect 33908 26124 33918 26180
rect 42466 26124 42476 26180
rect 42532 26124 43484 26180
rect 43540 26124 43550 26180
rect 46722 26124 46732 26180
rect 46788 26124 48860 26180
rect 48916 26124 48926 26180
rect 23986 26012 23996 26068
rect 24052 26012 27860 26068
rect 28018 26012 28028 26068
rect 28084 26012 29148 26068
rect 29204 26012 29214 26068
rect 29372 26012 36204 26068
rect 36260 26012 36270 26068
rect 27804 25956 27860 26012
rect 29372 25956 29428 26012
rect 15250 25900 15260 25956
rect 15316 25900 16044 25956
rect 16100 25900 25228 25956
rect 25284 25900 27356 25956
rect 27412 25900 27422 25956
rect 27804 25900 29428 25956
rect 37874 25900 37884 25956
rect 37940 25900 38220 25956
rect 38276 25900 38286 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 4834 25788 4844 25844
rect 4900 25788 6076 25844
rect 6132 25788 6142 25844
rect 22194 25788 22204 25844
rect 22260 25788 25900 25844
rect 25956 25788 25966 25844
rect 28578 25788 28588 25844
rect 28644 25788 29372 25844
rect 29428 25788 33068 25844
rect 33124 25788 33134 25844
rect 36754 25788 36764 25844
rect 36820 25788 37660 25844
rect 37716 25788 37726 25844
rect 37996 25788 41132 25844
rect 41188 25788 41198 25844
rect 4844 25732 4900 25788
rect 37996 25732 38052 25788
rect 4162 25676 4172 25732
rect 4228 25676 4900 25732
rect 5282 25676 5292 25732
rect 5348 25676 7196 25732
rect 7252 25676 7262 25732
rect 14466 25676 14476 25732
rect 14532 25676 16156 25732
rect 16212 25676 16222 25732
rect 24770 25676 24780 25732
rect 24836 25676 28812 25732
rect 28868 25676 28878 25732
rect 29810 25676 29820 25732
rect 29876 25676 31052 25732
rect 31108 25676 32060 25732
rect 32116 25676 32126 25732
rect 32834 25676 32844 25732
rect 32900 25676 37996 25732
rect 38052 25676 38062 25732
rect 38892 25676 39228 25732
rect 39284 25676 40348 25732
rect 40404 25676 42924 25732
rect 42980 25676 42990 25732
rect 46946 25676 46956 25732
rect 47012 25676 48748 25732
rect 48804 25676 48814 25732
rect 38892 25620 38948 25676
rect 3714 25564 3724 25620
rect 3780 25564 6300 25620
rect 6356 25564 6860 25620
rect 6916 25564 7644 25620
rect 7700 25564 7710 25620
rect 16818 25564 16828 25620
rect 16884 25564 17948 25620
rect 18004 25564 18508 25620
rect 18564 25564 21756 25620
rect 21812 25564 23436 25620
rect 23492 25564 23502 25620
rect 27794 25564 27804 25620
rect 27860 25564 28588 25620
rect 28644 25564 28654 25620
rect 33506 25564 33516 25620
rect 33572 25564 35532 25620
rect 35588 25564 35598 25620
rect 38882 25564 38892 25620
rect 38948 25564 38958 25620
rect 39778 25564 39788 25620
rect 39844 25564 39854 25620
rect 40898 25564 40908 25620
rect 40964 25564 44268 25620
rect 44324 25564 44334 25620
rect 48178 25564 48188 25620
rect 48244 25564 49084 25620
rect 49140 25564 49150 25620
rect 7074 25452 7084 25508
rect 7140 25452 8428 25508
rect 8484 25452 8494 25508
rect 9762 25452 9772 25508
rect 9828 25452 10444 25508
rect 10500 25452 10510 25508
rect 10770 25452 10780 25508
rect 10836 25452 12236 25508
rect 12292 25452 12302 25508
rect 12450 25452 12460 25508
rect 12516 25452 14140 25508
rect 14196 25452 14206 25508
rect 16706 25452 16716 25508
rect 16772 25452 17724 25508
rect 17780 25452 17790 25508
rect 18386 25452 18396 25508
rect 18452 25452 19292 25508
rect 19348 25452 19358 25508
rect 19618 25452 19628 25508
rect 19684 25452 20412 25508
rect 20468 25452 20478 25508
rect 20738 25452 20748 25508
rect 20804 25452 21980 25508
rect 22036 25452 22876 25508
rect 22932 25452 23996 25508
rect 24052 25452 25116 25508
rect 25172 25452 25182 25508
rect 28130 25452 28140 25508
rect 28196 25452 29260 25508
rect 29316 25452 29326 25508
rect 33730 25452 33740 25508
rect 33796 25452 34524 25508
rect 34580 25452 34590 25508
rect 34962 25452 34972 25508
rect 35028 25452 35644 25508
rect 35700 25452 36652 25508
rect 36708 25452 37212 25508
rect 37268 25452 37278 25508
rect 37426 25452 37436 25508
rect 37492 25452 37772 25508
rect 37828 25452 37838 25508
rect 38098 25452 38108 25508
rect 38164 25452 39564 25508
rect 39620 25452 39630 25508
rect 6402 25340 6412 25396
rect 6468 25340 8316 25396
rect 8372 25340 8382 25396
rect 16034 25340 16044 25396
rect 16100 25340 21196 25396
rect 21252 25340 22540 25396
rect 22596 25340 22606 25396
rect 22978 25340 22988 25396
rect 23044 25340 23772 25396
rect 23828 25340 23838 25396
rect 26674 25340 26684 25396
rect 26740 25340 27692 25396
rect 27748 25340 27758 25396
rect 30146 25340 30156 25396
rect 30212 25340 30222 25396
rect 33954 25340 33964 25396
rect 34020 25340 34300 25396
rect 34356 25340 34366 25396
rect 36418 25340 36428 25396
rect 36484 25340 38220 25396
rect 38276 25340 38286 25396
rect 38854 25340 38892 25396
rect 38948 25340 38958 25396
rect 30156 25284 30212 25340
rect 39788 25284 39844 25564
rect 40758 25452 40796 25508
rect 40852 25452 40862 25508
rect 41346 25452 41356 25508
rect 41412 25452 41916 25508
rect 41972 25452 43820 25508
rect 43876 25452 43886 25508
rect 40674 25340 40684 25396
rect 40740 25340 42028 25396
rect 42084 25340 43596 25396
rect 43652 25340 43662 25396
rect 47506 25340 47516 25396
rect 47572 25340 48188 25396
rect 48244 25340 48254 25396
rect 14802 25228 14812 25284
rect 14868 25228 16380 25284
rect 16436 25228 16446 25284
rect 17042 25228 17052 25284
rect 17108 25228 18284 25284
rect 18340 25228 18350 25284
rect 19628 25228 20076 25284
rect 20132 25228 20142 25284
rect 20290 25228 20300 25284
rect 20356 25228 22428 25284
rect 22484 25228 22652 25284
rect 22708 25228 23660 25284
rect 23716 25228 24444 25284
rect 24500 25228 24510 25284
rect 26852 25228 27804 25284
rect 27860 25228 30212 25284
rect 31574 25228 31612 25284
rect 31668 25228 31678 25284
rect 36306 25228 36316 25284
rect 36372 25228 36988 25284
rect 37044 25228 37054 25284
rect 37762 25228 37772 25284
rect 37828 25228 38332 25284
rect 38388 25228 39844 25284
rect 41458 25228 41468 25284
rect 41524 25228 42924 25284
rect 42980 25228 43932 25284
rect 43988 25228 43998 25284
rect 45826 25228 45836 25284
rect 45892 25228 45902 25284
rect 46386 25228 46396 25284
rect 46452 25228 46462 25284
rect 3938 25116 3948 25172
rect 4004 25116 5068 25172
rect 5124 25116 5134 25172
rect 16268 24948 16324 25228
rect 19628 25172 19684 25228
rect 26852 25172 26908 25228
rect 45836 25172 45892 25228
rect 46396 25172 46452 25228
rect 17826 25116 17836 25172
rect 17892 25116 19684 25172
rect 21634 25116 21644 25172
rect 21700 25116 26908 25172
rect 29250 25116 29260 25172
rect 29316 25116 30156 25172
rect 30212 25116 32396 25172
rect 32452 25116 33180 25172
rect 33236 25116 35980 25172
rect 36036 25116 36046 25172
rect 41906 25116 41916 25172
rect 41972 25116 42252 25172
rect 42308 25116 44828 25172
rect 44884 25116 44894 25172
rect 45836 25116 47740 25172
rect 47796 25116 47806 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 21084 25004 21420 25060
rect 21476 25004 22428 25060
rect 22484 25004 22494 25060
rect 29558 25004 29596 25060
rect 29652 25004 29662 25060
rect 21084 24948 21140 25004
rect 16268 24892 21140 24948
rect 21298 24892 21308 24948
rect 21364 24892 22764 24948
rect 22820 24892 22830 24948
rect 30818 24892 30828 24948
rect 30884 24892 31612 24948
rect 31668 24892 31678 24948
rect 31826 24892 31836 24948
rect 31892 24892 32956 24948
rect 33012 24892 33022 24948
rect 43698 24892 43708 24948
rect 43764 24892 47180 24948
rect 47236 24892 47246 24948
rect 14578 24780 14588 24836
rect 14644 24780 17836 24836
rect 17892 24780 17902 24836
rect 21186 24780 21196 24836
rect 21252 24780 26908 24836
rect 28578 24780 28588 24836
rect 28644 24780 28812 24836
rect 28868 24780 38668 24836
rect 41570 24780 41580 24836
rect 41636 24780 46284 24836
rect 46340 24780 46350 24836
rect 13010 24668 13020 24724
rect 13076 24668 23884 24724
rect 23940 24668 25228 24724
rect 25284 24668 25294 24724
rect 26852 24612 26908 24780
rect 29474 24668 29484 24724
rect 29540 24668 31388 24724
rect 31444 24668 32060 24724
rect 32116 24668 32126 24724
rect 38612 24612 38668 24780
rect 40002 24668 40012 24724
rect 40068 24668 42588 24724
rect 42644 24668 43484 24724
rect 43540 24668 43550 24724
rect 45826 24668 45836 24724
rect 45892 24668 47852 24724
rect 47908 24668 47918 24724
rect 48038 24668 48076 24724
rect 48132 24668 48142 24724
rect 2482 24556 2492 24612
rect 2548 24556 6188 24612
rect 6244 24556 6254 24612
rect 10770 24556 10780 24612
rect 10836 24556 11900 24612
rect 11956 24556 11966 24612
rect 14690 24556 14700 24612
rect 14756 24556 15260 24612
rect 15316 24556 15326 24612
rect 15586 24556 15596 24612
rect 15652 24556 16156 24612
rect 16212 24556 16222 24612
rect 26852 24556 30044 24612
rect 30100 24556 34188 24612
rect 34244 24556 34254 24612
rect 36418 24556 36428 24612
rect 36484 24556 37100 24612
rect 37156 24556 37166 24612
rect 38612 24556 41468 24612
rect 41524 24556 41534 24612
rect 41794 24556 41804 24612
rect 41860 24556 43372 24612
rect 43428 24556 43932 24612
rect 43988 24556 43998 24612
rect 44370 24556 44380 24612
rect 44436 24556 46172 24612
rect 46228 24556 46238 24612
rect 4610 24444 4620 24500
rect 4676 24444 5180 24500
rect 5236 24444 5246 24500
rect 11666 24444 11676 24500
rect 11732 24444 12012 24500
rect 12068 24444 12572 24500
rect 12628 24444 13916 24500
rect 13972 24444 13982 24500
rect 28550 24444 28588 24500
rect 28644 24444 28654 24500
rect 29810 24444 29820 24500
rect 29876 24444 30716 24500
rect 30772 24444 30782 24500
rect 31574 24444 31612 24500
rect 31668 24444 31678 24500
rect 47058 24444 47068 24500
rect 47124 24444 48748 24500
rect 48804 24444 48814 24500
rect 31686 24332 31724 24388
rect 31780 24332 31790 24388
rect 43026 24332 43036 24388
rect 43092 24332 47628 24388
rect 47684 24332 48300 24388
rect 48356 24332 48366 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 12114 24220 12124 24276
rect 12180 24220 13468 24276
rect 13524 24220 13534 24276
rect 21522 24220 21532 24276
rect 21588 24220 23436 24276
rect 23492 24220 23502 24276
rect 4610 24108 4620 24164
rect 4676 24108 5404 24164
rect 5460 24108 5470 24164
rect 12898 24108 12908 24164
rect 12964 24108 14028 24164
rect 14084 24108 14094 24164
rect 16482 24108 16492 24164
rect 16548 24108 17164 24164
rect 17220 24108 17230 24164
rect 20132 24108 20748 24164
rect 20804 24108 20814 24164
rect 33954 24108 33964 24164
rect 34020 24108 34860 24164
rect 34916 24108 34926 24164
rect 20132 24052 20188 24108
rect 5954 23996 5964 24052
rect 6020 23996 6636 24052
rect 6692 23996 7868 24052
rect 7924 23996 7934 24052
rect 10994 23996 11004 24052
rect 11060 23996 12348 24052
rect 12404 23996 12414 24052
rect 17042 23996 17052 24052
rect 17108 23996 20188 24052
rect 20850 23996 20860 24052
rect 20916 23996 21532 24052
rect 21588 23996 21598 24052
rect 26852 23996 31948 24052
rect 32004 23996 32014 24052
rect 36082 23996 36092 24052
rect 36148 23996 37324 24052
rect 37380 23996 37390 24052
rect 42018 23996 42028 24052
rect 42084 23996 49196 24052
rect 49252 23996 49262 24052
rect 5170 23884 5180 23940
rect 5236 23884 5628 23940
rect 5684 23884 5694 23940
rect 6290 23884 6300 23940
rect 6356 23884 9100 23940
rect 9156 23884 9166 23940
rect 12002 23884 12012 23940
rect 12068 23884 12236 23940
rect 12292 23884 14252 23940
rect 14308 23884 15484 23940
rect 15540 23884 15550 23940
rect 17490 23884 17500 23940
rect 17556 23884 19404 23940
rect 19460 23884 19470 23940
rect 22866 23884 22876 23940
rect 22932 23884 24780 23940
rect 24836 23884 26460 23940
rect 26516 23884 26526 23940
rect 4834 23772 4844 23828
rect 4900 23772 6188 23828
rect 6244 23772 6254 23828
rect 7746 23772 7756 23828
rect 7812 23772 8428 23828
rect 13122 23772 13132 23828
rect 13188 23772 14028 23828
rect 14084 23772 15036 23828
rect 15092 23772 15102 23828
rect 15250 23772 15260 23828
rect 15316 23772 16604 23828
rect 16660 23772 16670 23828
rect 8372 23716 8428 23772
rect 8372 23660 8764 23716
rect 8820 23660 8830 23716
rect 26852 23604 26908 23996
rect 27010 23884 27020 23940
rect 27076 23884 27086 23940
rect 28018 23884 28028 23940
rect 28084 23884 28588 23940
rect 28644 23884 28654 23940
rect 34962 23884 34972 23940
rect 35028 23884 35038 23940
rect 35186 23884 35196 23940
rect 35252 23884 36876 23940
rect 36932 23884 37548 23940
rect 37604 23884 37614 23940
rect 37874 23884 37884 23940
rect 37940 23884 38556 23940
rect 38612 23884 38622 23940
rect 43474 23884 43484 23940
rect 43540 23884 44828 23940
rect 44884 23884 44894 23940
rect 26226 23548 26236 23604
rect 26292 23548 26908 23604
rect 27020 23604 27076 23884
rect 34972 23828 35028 23884
rect 28354 23772 28364 23828
rect 28420 23772 29484 23828
rect 29540 23772 29550 23828
rect 30370 23772 30380 23828
rect 30436 23772 30828 23828
rect 30884 23772 30894 23828
rect 34972 23772 35868 23828
rect 35924 23772 37772 23828
rect 37828 23772 37838 23828
rect 38612 23772 40236 23828
rect 40292 23772 40302 23828
rect 47842 23772 47852 23828
rect 47908 23772 48524 23828
rect 48580 23772 48590 23828
rect 38612 23716 38668 23772
rect 28018 23660 28028 23716
rect 28084 23660 28476 23716
rect 28532 23660 38668 23716
rect 38994 23660 39004 23716
rect 39060 23660 40348 23716
rect 40404 23660 40414 23716
rect 41010 23660 41020 23716
rect 41076 23660 44156 23716
rect 44212 23660 45500 23716
rect 45556 23660 45566 23716
rect 40348 23604 40404 23660
rect 27020 23548 29260 23604
rect 29316 23548 29764 23604
rect 40348 23548 42028 23604
rect 42084 23548 42094 23604
rect 43138 23548 43148 23604
rect 43204 23548 43214 23604
rect 44930 23548 44940 23604
rect 44996 23548 46116 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 15026 23436 15036 23492
rect 15092 23436 15820 23492
rect 15876 23436 15886 23492
rect 28130 23436 28140 23492
rect 28196 23436 28924 23492
rect 28980 23436 28990 23492
rect 29708 23380 29764 23548
rect 43148 23492 43204 23548
rect 46060 23492 46116 23548
rect 29922 23436 29932 23492
rect 29988 23436 31500 23492
rect 31556 23436 33516 23492
rect 33572 23436 33582 23492
rect 33954 23436 33964 23492
rect 34020 23436 34412 23492
rect 34468 23436 34478 23492
rect 37762 23436 37772 23492
rect 37828 23436 39116 23492
rect 39172 23436 39182 23492
rect 41682 23436 41692 23492
rect 41748 23436 43372 23492
rect 43428 23436 43438 23492
rect 46050 23436 46060 23492
rect 46116 23436 46126 23492
rect 50200 23380 51000 23408
rect 2482 23324 2492 23380
rect 2548 23324 4284 23380
rect 4340 23324 4350 23380
rect 29708 23324 30268 23380
rect 30324 23324 31164 23380
rect 31220 23324 31230 23380
rect 33590 23324 33628 23380
rect 33684 23324 33694 23380
rect 34514 23324 34524 23380
rect 34580 23324 35084 23380
rect 35140 23324 35150 23380
rect 38882 23324 38892 23380
rect 38948 23324 41804 23380
rect 41860 23324 41870 23380
rect 48066 23324 48076 23380
rect 48132 23324 51000 23380
rect 50200 23296 51000 23324
rect 3378 23212 3388 23268
rect 3444 23212 4844 23268
rect 4900 23212 4910 23268
rect 12002 23212 12012 23268
rect 12068 23212 13132 23268
rect 13188 23212 13198 23268
rect 27794 23212 27804 23268
rect 27860 23212 28924 23268
rect 28980 23212 28990 23268
rect 30482 23212 30492 23268
rect 30548 23212 31948 23268
rect 32004 23212 38220 23268
rect 38276 23212 38286 23268
rect 4050 23100 4060 23156
rect 4116 23100 5292 23156
rect 5348 23100 5358 23156
rect 19170 23100 19180 23156
rect 19236 23100 21196 23156
rect 21252 23100 21262 23156
rect 35410 23100 35420 23156
rect 35476 23100 35644 23156
rect 35700 23100 35710 23156
rect 38322 23100 38332 23156
rect 38388 23100 39676 23156
rect 39732 23100 39742 23156
rect 2818 22988 2828 23044
rect 2884 22988 3500 23044
rect 3556 22988 3566 23044
rect 14578 22988 14588 23044
rect 14644 22988 15484 23044
rect 15540 22988 16044 23044
rect 16100 22988 16110 23044
rect 18498 22988 18508 23044
rect 18564 22988 20188 23044
rect 20934 22988 20972 23044
rect 21028 22988 21038 23044
rect 33842 22988 33852 23044
rect 33908 22988 33918 23044
rect 34188 22988 34748 23044
rect 34804 22988 35980 23044
rect 36036 22988 36046 23044
rect 42578 22988 42588 23044
rect 42644 22988 42812 23044
rect 42868 22988 43596 23044
rect 43652 22988 43662 23044
rect 20132 22932 20188 22988
rect 17266 22876 17276 22932
rect 17332 22876 19404 22932
rect 19460 22876 19470 22932
rect 20132 22876 33516 22932
rect 33572 22876 33582 22932
rect 33852 22820 33908 22988
rect 34188 22932 34244 22988
rect 34178 22876 34188 22932
rect 34244 22876 34254 22932
rect 34514 22876 34524 22932
rect 34580 22876 37324 22932
rect 37380 22876 37390 22932
rect 34524 22820 34580 22876
rect 22866 22764 22876 22820
rect 22932 22764 30492 22820
rect 30548 22764 30558 22820
rect 33590 22764 33628 22820
rect 33684 22764 33694 22820
rect 33852 22764 34580 22820
rect 35634 22764 35644 22820
rect 35700 22764 36876 22820
rect 36932 22764 39228 22820
rect 39284 22764 39294 22820
rect 43026 22764 43036 22820
rect 43092 22764 43372 22820
rect 43428 22764 43438 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 8978 22652 8988 22708
rect 9044 22652 11004 22708
rect 11060 22652 11070 22708
rect 20178 22652 20188 22708
rect 20244 22652 20282 22708
rect 20598 22652 20636 22708
rect 20692 22652 21644 22708
rect 21700 22652 21710 22708
rect 38612 22652 44604 22708
rect 44660 22652 44670 22708
rect 38612 22596 38668 22652
rect 3602 22540 3612 22596
rect 3668 22540 4620 22596
rect 4676 22540 5404 22596
rect 5460 22540 5470 22596
rect 17042 22540 17052 22596
rect 17108 22540 38668 22596
rect 38882 22540 38892 22596
rect 38948 22540 40908 22596
rect 40964 22540 40974 22596
rect 44146 22540 44156 22596
rect 44212 22540 45388 22596
rect 45444 22540 45454 22596
rect 21746 22428 21756 22484
rect 21812 22428 23772 22484
rect 23828 22428 23838 22484
rect 24210 22428 24220 22484
rect 24276 22428 24668 22484
rect 24724 22428 25340 22484
rect 25396 22428 25676 22484
rect 25732 22428 25742 22484
rect 27346 22428 27356 22484
rect 27412 22428 28476 22484
rect 28532 22428 29260 22484
rect 29316 22428 29326 22484
rect 34626 22428 34636 22484
rect 34692 22428 36764 22484
rect 36820 22428 36830 22484
rect 39218 22428 39228 22484
rect 39284 22428 44940 22484
rect 44996 22428 45006 22484
rect 6626 22316 6636 22372
rect 6692 22316 10332 22372
rect 10388 22316 11340 22372
rect 11396 22316 11406 22372
rect 30902 22316 30940 22372
rect 30996 22316 31006 22372
rect 34178 22316 34188 22372
rect 34244 22316 36204 22372
rect 36260 22316 36270 22372
rect 40226 22316 40236 22372
rect 40292 22316 42140 22372
rect 42196 22316 42206 22372
rect 42578 22316 42588 22372
rect 42644 22316 45948 22372
rect 46004 22316 46014 22372
rect 19058 22204 19068 22260
rect 19124 22204 21084 22260
rect 21140 22204 21150 22260
rect 22754 22204 22764 22260
rect 22820 22204 23884 22260
rect 23940 22204 23950 22260
rect 26002 22204 26012 22260
rect 26068 22204 26460 22260
rect 26516 22204 26526 22260
rect 32162 22204 32172 22260
rect 32228 22204 32620 22260
rect 32676 22204 33068 22260
rect 33124 22204 33134 22260
rect 37090 22204 37100 22260
rect 37156 22204 39228 22260
rect 39284 22204 39294 22260
rect 40674 22204 40684 22260
rect 40740 22204 40908 22260
rect 40964 22204 40974 22260
rect 19506 22092 19516 22148
rect 19572 22092 20076 22148
rect 20132 22092 20142 22148
rect 31826 22092 31836 22148
rect 31892 22092 31902 22148
rect 36418 22092 36428 22148
rect 36484 22092 37212 22148
rect 37268 22092 37278 22148
rect 45490 22092 45500 22148
rect 45556 22092 47292 22148
rect 47348 22092 47358 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 24882 21868 24892 21924
rect 24948 21868 29372 21924
rect 29428 21868 29438 21924
rect 31836 21812 31892 22092
rect 33926 21868 33964 21924
rect 34020 21868 34030 21924
rect 34150 21868 34188 21924
rect 34244 21868 34254 21924
rect 37314 21868 37324 21924
rect 37380 21868 38108 21924
rect 38164 21868 38174 21924
rect 39890 21868 39900 21924
rect 39956 21868 40236 21924
rect 40292 21868 40302 21924
rect 3938 21756 3948 21812
rect 4004 21756 5516 21812
rect 5572 21756 6188 21812
rect 6244 21756 6748 21812
rect 6804 21756 6814 21812
rect 8754 21756 8764 21812
rect 8820 21756 9660 21812
rect 9716 21756 9726 21812
rect 11442 21756 11452 21812
rect 11508 21756 14028 21812
rect 14084 21756 14094 21812
rect 18946 21756 18956 21812
rect 19012 21756 20860 21812
rect 20916 21756 20926 21812
rect 23538 21756 23548 21812
rect 23604 21756 25788 21812
rect 25844 21756 25854 21812
rect 27458 21756 27468 21812
rect 27524 21756 28588 21812
rect 28644 21756 28654 21812
rect 29698 21756 29708 21812
rect 29764 21756 31892 21812
rect 32162 21756 32172 21812
rect 32228 21756 33068 21812
rect 33124 21756 33134 21812
rect 35970 21756 35980 21812
rect 36036 21756 36988 21812
rect 37044 21756 37054 21812
rect 37510 21756 37548 21812
rect 37604 21756 37614 21812
rect 40114 21756 40124 21812
rect 40180 21756 41356 21812
rect 41412 21756 41422 21812
rect 46834 21756 46844 21812
rect 46900 21756 47740 21812
rect 47796 21756 47806 21812
rect 10210 21644 10220 21700
rect 10276 21644 10892 21700
rect 10948 21644 10958 21700
rect 19394 21644 19404 21700
rect 19460 21644 21196 21700
rect 21252 21644 21262 21700
rect 21532 21644 49420 21700
rect 49476 21644 49486 21700
rect 21532 21588 21588 21644
rect 16034 21532 16044 21588
rect 16100 21532 21588 21588
rect 21746 21532 21756 21588
rect 21812 21532 23996 21588
rect 24052 21532 24062 21588
rect 24546 21532 24556 21588
rect 24612 21532 27468 21588
rect 27524 21532 27534 21588
rect 29474 21532 29484 21588
rect 29540 21532 29550 21588
rect 30258 21532 30268 21588
rect 30324 21532 30940 21588
rect 30996 21532 31006 21588
rect 31490 21532 31500 21588
rect 31556 21532 31836 21588
rect 31892 21532 31902 21588
rect 32498 21532 32508 21588
rect 32564 21532 35084 21588
rect 35140 21532 36820 21588
rect 40898 21532 40908 21588
rect 40964 21532 42028 21588
rect 42084 21532 42094 21588
rect 42354 21532 42364 21588
rect 42420 21532 43036 21588
rect 43092 21532 43102 21588
rect 46722 21532 46732 21588
rect 46788 21532 47516 21588
rect 47572 21532 48636 21588
rect 48692 21532 48702 21588
rect 29484 21476 29540 21532
rect 11218 21420 11228 21476
rect 11284 21420 11788 21476
rect 11844 21420 11854 21476
rect 16482 21420 16492 21476
rect 16548 21420 18396 21476
rect 18452 21420 18462 21476
rect 19618 21420 19628 21476
rect 19684 21420 20412 21476
rect 20468 21420 21308 21476
rect 21364 21420 22652 21476
rect 22708 21420 22718 21476
rect 26114 21420 26124 21476
rect 26180 21420 26852 21476
rect 26908 21420 26918 21476
rect 27010 21420 27020 21476
rect 27076 21420 29540 21476
rect 29922 21420 29932 21476
rect 29988 21420 31388 21476
rect 31444 21420 31612 21476
rect 31668 21420 32396 21476
rect 32452 21420 32462 21476
rect 33842 21420 33852 21476
rect 33908 21420 34636 21476
rect 34692 21420 34702 21476
rect 35746 21420 35756 21476
rect 35812 21420 36092 21476
rect 36148 21420 36428 21476
rect 36484 21420 36494 21476
rect 36764 21364 36820 21532
rect 38210 21420 38220 21476
rect 38276 21420 39452 21476
rect 39508 21420 39518 21476
rect 6514 21308 6524 21364
rect 6580 21308 9660 21364
rect 9716 21308 9726 21364
rect 17378 21308 17388 21364
rect 17444 21308 21532 21364
rect 21588 21308 21598 21364
rect 23314 21308 23324 21364
rect 23380 21308 27356 21364
rect 27412 21308 27422 21364
rect 28242 21308 28252 21364
rect 28308 21308 29596 21364
rect 29652 21308 29662 21364
rect 34066 21308 34076 21364
rect 34132 21308 34142 21364
rect 34300 21308 35868 21364
rect 35924 21308 35934 21364
rect 36754 21308 36764 21364
rect 36820 21308 41468 21364
rect 41524 21308 41534 21364
rect 34076 21252 34132 21308
rect 16818 21196 16828 21252
rect 16884 21196 17948 21252
rect 18004 21196 22988 21252
rect 23044 21196 23054 21252
rect 23202 21196 23212 21252
rect 23268 21196 34132 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 34300 21140 34356 21308
rect 37874 21196 37884 21252
rect 37940 21196 39340 21252
rect 39396 21196 40124 21252
rect 40180 21196 40190 21252
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 19170 21084 19180 21140
rect 19236 21084 21756 21140
rect 21812 21084 23436 21140
rect 23492 21084 23502 21140
rect 26898 21084 26908 21140
rect 26964 21084 29708 21140
rect 29764 21084 29774 21140
rect 33954 21084 33964 21140
rect 34020 21084 34188 21140
rect 34244 21084 34356 21140
rect 20132 20972 20636 21028
rect 20692 20972 20702 21028
rect 25778 20972 25788 21028
rect 25844 20972 27356 21028
rect 27412 20972 27422 21028
rect 28690 20972 28700 21028
rect 28756 20972 29820 21028
rect 29876 20972 30156 21028
rect 30212 20972 30222 21028
rect 35522 20972 35532 21028
rect 35588 20972 35980 21028
rect 36036 20972 36046 21028
rect 20132 20916 20188 20972
rect 18162 20860 18172 20916
rect 18228 20860 20188 20916
rect 22306 20860 22316 20916
rect 22372 20860 22876 20916
rect 22932 20860 22942 20916
rect 24546 20860 24556 20916
rect 24612 20860 25900 20916
rect 25956 20860 25966 20916
rect 28018 20860 28028 20916
rect 28084 20860 30268 20916
rect 30324 20860 30334 20916
rect 30706 20860 30716 20916
rect 30772 20860 31276 20916
rect 31332 20860 33068 20916
rect 33124 20860 33134 20916
rect 1810 20748 1820 20804
rect 1876 20748 3948 20804
rect 4004 20748 4014 20804
rect 10098 20748 10108 20804
rect 10164 20748 11116 20804
rect 11172 20748 12684 20804
rect 12740 20748 14140 20804
rect 14196 20748 14206 20804
rect 17042 20748 17052 20804
rect 17108 20748 19740 20804
rect 19796 20748 19806 20804
rect 26114 20748 26124 20804
rect 26180 20748 27244 20804
rect 27300 20748 27310 20804
rect 35186 20748 35196 20804
rect 35252 20748 36988 20804
rect 37044 20748 37054 20804
rect 37314 20748 37324 20804
rect 37380 20748 38332 20804
rect 38388 20748 38398 20804
rect 38658 20748 38668 20804
rect 38724 20748 39676 20804
rect 39732 20748 39742 20804
rect 42018 20748 42028 20804
rect 42084 20748 42588 20804
rect 42644 20748 43148 20804
rect 43204 20748 43214 20804
rect 45714 20748 45724 20804
rect 45780 20748 46844 20804
rect 46900 20748 46910 20804
rect 16594 20636 16604 20692
rect 16660 20636 17388 20692
rect 17444 20636 19628 20692
rect 19684 20636 19694 20692
rect 20738 20636 20748 20692
rect 20804 20636 23212 20692
rect 23268 20636 23278 20692
rect 26852 20636 27580 20692
rect 27636 20636 27916 20692
rect 27972 20636 27982 20692
rect 33618 20636 33628 20692
rect 33684 20636 37548 20692
rect 37604 20636 39564 20692
rect 39620 20636 39630 20692
rect 40422 20636 40460 20692
rect 40516 20636 40526 20692
rect 42354 20636 42364 20692
rect 42420 20636 44044 20692
rect 44100 20636 44110 20692
rect 26852 20580 26908 20636
rect 14914 20524 14924 20580
rect 14980 20524 17836 20580
rect 17892 20524 17902 20580
rect 25218 20524 25228 20580
rect 25284 20524 26124 20580
rect 26180 20524 26908 20580
rect 28354 20524 28364 20580
rect 28420 20524 29708 20580
rect 29764 20524 29774 20580
rect 30034 20524 30044 20580
rect 30100 20524 31612 20580
rect 31668 20524 31678 20580
rect 34290 20524 34300 20580
rect 34356 20524 34748 20580
rect 34804 20524 34814 20580
rect 35746 20524 35756 20580
rect 35812 20524 37548 20580
rect 37604 20524 39228 20580
rect 39284 20524 39294 20580
rect 40674 20524 40684 20580
rect 40740 20524 41356 20580
rect 41412 20524 41422 20580
rect 43362 20524 43372 20580
rect 43428 20524 44828 20580
rect 44884 20524 44894 20580
rect 39452 20412 42812 20468
rect 42868 20412 43260 20468
rect 43316 20412 43326 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 39452 20356 39508 20412
rect 15362 20300 15372 20356
rect 15428 20300 19516 20356
rect 19572 20300 19582 20356
rect 27234 20300 27244 20356
rect 27300 20300 27916 20356
rect 27972 20300 27982 20356
rect 32610 20300 32620 20356
rect 32676 20300 39508 20356
rect 39666 20300 39676 20356
rect 39732 20300 41020 20356
rect 41076 20300 41086 20356
rect 8306 20188 8316 20244
rect 8372 20188 10556 20244
rect 10612 20188 10622 20244
rect 23986 20188 23996 20244
rect 24052 20188 27692 20244
rect 27748 20188 28252 20244
rect 28308 20188 28318 20244
rect 31892 20188 33852 20244
rect 33908 20188 33918 20244
rect 34290 20188 34300 20244
rect 34356 20188 35868 20244
rect 35924 20188 35934 20244
rect 37874 20188 37884 20244
rect 37940 20188 40908 20244
rect 40964 20188 40974 20244
rect 41356 20188 42252 20244
rect 42308 20188 42318 20244
rect 47058 20188 47068 20244
rect 47124 20188 48748 20244
rect 48804 20188 48814 20244
rect 31892 20132 31948 20188
rect 2482 20076 2492 20132
rect 2548 20076 4620 20132
rect 4676 20076 5068 20132
rect 5124 20076 7420 20132
rect 7476 20076 7486 20132
rect 13794 20076 13804 20132
rect 13860 20076 14140 20132
rect 14196 20076 15932 20132
rect 15988 20076 15998 20132
rect 23090 20076 23100 20132
rect 23156 20076 23660 20132
rect 23716 20076 23726 20132
rect 24210 20076 24220 20132
rect 24276 20076 24668 20132
rect 24724 20076 31948 20132
rect 36978 20076 36988 20132
rect 37044 20076 39676 20132
rect 39732 20076 39742 20132
rect 41356 20020 41412 20188
rect 41570 20076 41580 20132
rect 41636 20076 42588 20132
rect 42644 20076 44940 20132
rect 44996 20076 45006 20132
rect 45154 20076 45164 20132
rect 45220 20076 46284 20132
rect 46340 20076 46350 20132
rect 49074 20076 49084 20132
rect 49140 20076 49644 20132
rect 49700 20076 49710 20132
rect 13682 19964 13692 20020
rect 13748 19964 14364 20020
rect 14420 19964 16044 20020
rect 16100 19964 16110 20020
rect 21970 19964 21980 20020
rect 22036 19964 23884 20020
rect 23940 19964 23950 20020
rect 31042 19964 31052 20020
rect 31108 19964 33236 20020
rect 34178 19964 34188 20020
rect 34244 19964 34524 20020
rect 34580 19964 38220 20020
rect 38276 19964 38286 20020
rect 38612 19964 41412 20020
rect 43026 19964 43036 20020
rect 43092 19964 43596 20020
rect 43652 19964 43662 20020
rect 45042 19964 45052 20020
rect 45108 19964 45724 20020
rect 45780 19964 46732 20020
rect 46788 19964 46798 20020
rect 33180 19908 33236 19964
rect 38612 19908 38668 19964
rect 4610 19852 4620 19908
rect 4676 19852 5964 19908
rect 6020 19852 6030 19908
rect 15138 19852 15148 19908
rect 15204 19852 16828 19908
rect 16884 19852 16894 19908
rect 23426 19852 23436 19908
rect 23492 19852 27132 19908
rect 27188 19852 27198 19908
rect 33170 19852 33180 19908
rect 33236 19852 38668 19908
rect 41356 19852 42476 19908
rect 42532 19852 43260 19908
rect 43316 19852 43326 19908
rect 44034 19852 44044 19908
rect 44100 19852 45612 19908
rect 45668 19852 45678 19908
rect 46050 19852 46060 19908
rect 46116 19852 48748 19908
rect 48804 19852 48814 19908
rect 41356 19796 41412 19852
rect 7522 19740 7532 19796
rect 7588 19740 8652 19796
rect 8708 19740 8718 19796
rect 12786 19740 12796 19796
rect 12852 19740 13916 19796
rect 13972 19740 13982 19796
rect 15474 19740 15484 19796
rect 15540 19740 16044 19796
rect 16100 19740 16110 19796
rect 16258 19740 16268 19796
rect 16324 19740 16716 19796
rect 16772 19740 16782 19796
rect 31602 19740 31612 19796
rect 31668 19740 34636 19796
rect 34692 19740 34702 19796
rect 41010 19740 41020 19796
rect 41076 19740 41356 19796
rect 41412 19740 41422 19796
rect 42242 19740 42252 19796
rect 42308 19740 42700 19796
rect 42756 19740 45052 19796
rect 45108 19740 45118 19796
rect 14690 19628 14700 19684
rect 14756 19628 15372 19684
rect 15428 19628 17724 19684
rect 17780 19628 17790 19684
rect 28466 19628 28476 19684
rect 28532 19628 30604 19684
rect 30660 19628 30670 19684
rect 40338 19628 40348 19684
rect 40404 19628 42028 19684
rect 42084 19628 42924 19684
rect 42980 19628 42990 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 22978 19516 22988 19572
rect 23044 19516 23436 19572
rect 23492 19516 23502 19572
rect 26852 19516 29932 19572
rect 29988 19516 29998 19572
rect 37426 19516 37436 19572
rect 37492 19516 37884 19572
rect 37940 19516 37950 19572
rect 38612 19516 44268 19572
rect 44324 19516 44334 19572
rect 26852 19460 26908 19516
rect 38612 19460 38668 19516
rect 19058 19404 19068 19460
rect 19124 19404 22428 19460
rect 22484 19404 22494 19460
rect 24994 19404 25004 19460
rect 25060 19404 26236 19460
rect 26292 19404 26908 19460
rect 28018 19404 28028 19460
rect 28084 19404 29596 19460
rect 29652 19404 29662 19460
rect 30566 19404 30604 19460
rect 30660 19404 30670 19460
rect 33506 19404 33516 19460
rect 33572 19404 38668 19460
rect 41234 19404 41244 19460
rect 41300 19404 41804 19460
rect 41860 19404 41870 19460
rect 5842 19292 5852 19348
rect 5908 19292 8316 19348
rect 8372 19292 8382 19348
rect 18386 19292 18396 19348
rect 18452 19292 20972 19348
rect 21028 19292 21038 19348
rect 21298 19292 21308 19348
rect 21364 19292 21756 19348
rect 21812 19292 24332 19348
rect 24388 19292 24398 19348
rect 25442 19292 25452 19348
rect 25508 19292 25900 19348
rect 25956 19292 25966 19348
rect 28214 19292 28252 19348
rect 28308 19292 28318 19348
rect 28578 19292 28588 19348
rect 28644 19292 29708 19348
rect 29764 19292 29774 19348
rect 30454 19292 30492 19348
rect 30548 19292 30558 19348
rect 31238 19292 31276 19348
rect 31332 19292 31342 19348
rect 32050 19292 32060 19348
rect 32116 19292 43036 19348
rect 43092 19292 43102 19348
rect 47842 19292 47852 19348
rect 47908 19292 49196 19348
rect 49252 19292 49262 19348
rect 6066 19180 6076 19236
rect 6132 19180 7420 19236
rect 7476 19180 7486 19236
rect 8866 19180 8876 19236
rect 8932 19180 9436 19236
rect 9492 19180 9502 19236
rect 14018 19180 14028 19236
rect 14084 19180 14812 19236
rect 14868 19180 14878 19236
rect 18722 19180 18732 19236
rect 18788 19180 20076 19236
rect 20132 19180 21196 19236
rect 21252 19180 21262 19236
rect 21522 19180 21532 19236
rect 21588 19180 22316 19236
rect 22372 19180 22382 19236
rect 26450 19180 26460 19236
rect 26516 19180 26796 19236
rect 26852 19180 26862 19236
rect 27010 19180 27020 19236
rect 27076 19180 27244 19236
rect 27300 19180 29148 19236
rect 29204 19180 29214 19236
rect 29484 19180 32620 19236
rect 32676 19180 32686 19236
rect 34626 19180 34636 19236
rect 34692 19180 35420 19236
rect 35476 19180 35486 19236
rect 43586 19180 43596 19236
rect 43652 19180 45500 19236
rect 45556 19180 45566 19236
rect 29484 19124 29540 19180
rect 50200 19124 51000 19152
rect 6738 19068 6748 19124
rect 6804 19068 9772 19124
rect 9828 19068 9838 19124
rect 13794 19068 13804 19124
rect 13860 19068 16268 19124
rect 16324 19068 16334 19124
rect 22754 19068 22764 19124
rect 22820 19068 23548 19124
rect 23604 19068 23614 19124
rect 25442 19068 25452 19124
rect 25508 19068 26012 19124
rect 26068 19068 26078 19124
rect 29474 19068 29484 19124
rect 29540 19068 29550 19124
rect 30258 19068 30268 19124
rect 30324 19068 31388 19124
rect 31444 19068 31454 19124
rect 37426 19068 37436 19124
rect 37492 19068 37996 19124
rect 38052 19068 38062 19124
rect 38546 19068 38556 19124
rect 38612 19068 39228 19124
rect 39284 19068 39294 19124
rect 44258 19068 44268 19124
rect 44324 19068 51000 19124
rect 29484 19012 29540 19068
rect 50200 19040 51000 19068
rect 12114 18956 12124 19012
rect 12180 18956 14252 19012
rect 14308 18956 14318 19012
rect 20962 18956 20972 19012
rect 21028 18956 24444 19012
rect 24500 18956 25564 19012
rect 25620 18956 25630 19012
rect 25778 18956 25788 19012
rect 25844 18956 28588 19012
rect 28644 18956 28654 19012
rect 28924 18956 29540 19012
rect 29698 18956 29708 19012
rect 29764 18956 30044 19012
rect 30100 18956 30110 19012
rect 30370 18956 30380 19012
rect 30436 18956 30446 19012
rect 30818 18956 30828 19012
rect 30884 18956 31164 19012
rect 31220 18956 31230 19012
rect 32162 18956 32172 19012
rect 32228 18956 33852 19012
rect 33908 18956 33918 19012
rect 34402 18956 34412 19012
rect 34468 18956 38444 19012
rect 38500 18956 38510 19012
rect 42466 18956 42476 19012
rect 42532 18956 42924 19012
rect 42980 18956 42990 19012
rect 46162 18956 46172 19012
rect 46228 18956 47852 19012
rect 47908 18956 47918 19012
rect 28924 18900 28980 18956
rect 24322 18844 24332 18900
rect 24388 18844 28140 18900
rect 28196 18844 28980 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 30380 18788 30436 18956
rect 31266 18844 31276 18900
rect 31332 18844 32844 18900
rect 32900 18844 32910 18900
rect 35858 18844 35868 18900
rect 35924 18844 43932 18900
rect 43988 18844 43998 18900
rect 44146 18844 44156 18900
rect 44212 18844 48748 18900
rect 48804 18844 48814 18900
rect 23650 18732 23660 18788
rect 23716 18732 28700 18788
rect 28756 18732 32060 18788
rect 32116 18732 32126 18788
rect 2594 18620 2604 18676
rect 2660 18620 4620 18676
rect 4676 18620 4686 18676
rect 13570 18620 13580 18676
rect 13636 18620 17276 18676
rect 17332 18620 17612 18676
rect 17668 18620 17678 18676
rect 18722 18620 18732 18676
rect 18788 18620 19404 18676
rect 19460 18620 19470 18676
rect 30604 18620 31612 18676
rect 31668 18620 31948 18676
rect 32004 18620 32014 18676
rect 30604 18564 30660 18620
rect 3042 18508 3052 18564
rect 3108 18508 4284 18564
rect 4340 18508 4350 18564
rect 13906 18508 13916 18564
rect 13972 18508 15148 18564
rect 15204 18508 15708 18564
rect 15764 18508 15774 18564
rect 17490 18508 17500 18564
rect 17556 18508 19180 18564
rect 19236 18508 19246 18564
rect 27570 18508 27580 18564
rect 27636 18508 29372 18564
rect 29428 18508 30604 18564
rect 30660 18508 30670 18564
rect 30818 18508 30828 18564
rect 30884 18508 32508 18564
rect 32564 18508 32574 18564
rect 35980 18508 36876 18564
rect 36932 18508 37548 18564
rect 37604 18508 37614 18564
rect 41906 18508 41916 18564
rect 41972 18508 43036 18564
rect 43092 18508 43102 18564
rect 43474 18508 43484 18564
rect 43540 18508 45780 18564
rect 45938 18508 45948 18564
rect 46004 18508 46508 18564
rect 46564 18508 46574 18564
rect 35980 18452 36036 18508
rect 44268 18452 44324 18508
rect 2258 18396 2268 18452
rect 2324 18396 3724 18452
rect 3780 18396 3790 18452
rect 3938 18396 3948 18452
rect 4004 18396 5516 18452
rect 5572 18396 5582 18452
rect 7746 18396 7756 18452
rect 7812 18396 9548 18452
rect 9604 18396 9614 18452
rect 14802 18396 14812 18452
rect 14868 18396 15260 18452
rect 15316 18396 15326 18452
rect 16482 18396 16492 18452
rect 16548 18396 18060 18452
rect 18116 18396 19740 18452
rect 19796 18396 19806 18452
rect 25330 18396 25340 18452
rect 25396 18396 27692 18452
rect 27748 18396 27758 18452
rect 28914 18396 28924 18452
rect 28980 18396 29260 18452
rect 29316 18396 29326 18452
rect 29810 18396 29820 18452
rect 29876 18396 31052 18452
rect 31108 18396 31118 18452
rect 33170 18396 33180 18452
rect 33236 18396 33964 18452
rect 34020 18396 34030 18452
rect 35970 18396 35980 18452
rect 36036 18396 36046 18452
rect 40226 18396 40236 18452
rect 40292 18396 42028 18452
rect 42084 18396 42094 18452
rect 42354 18396 42364 18452
rect 42420 18396 42812 18452
rect 42868 18396 42878 18452
rect 44258 18396 44268 18452
rect 44324 18396 44334 18452
rect 45724 18340 45780 18508
rect 2706 18284 2716 18340
rect 2772 18284 3612 18340
rect 3668 18284 3678 18340
rect 7858 18284 7868 18340
rect 7924 18284 10220 18340
rect 10276 18284 15036 18340
rect 15092 18284 15102 18340
rect 17826 18284 17836 18340
rect 17892 18284 18620 18340
rect 18676 18284 18686 18340
rect 20402 18284 20412 18340
rect 20468 18284 26572 18340
rect 26628 18284 26638 18340
rect 27804 18284 29036 18340
rect 29092 18284 30604 18340
rect 30660 18284 30670 18340
rect 34514 18284 34524 18340
rect 34580 18284 36092 18340
rect 36148 18284 36158 18340
rect 36316 18284 36988 18340
rect 37044 18284 37054 18340
rect 40450 18284 40460 18340
rect 40516 18284 42140 18340
rect 42196 18284 42206 18340
rect 45714 18284 45724 18340
rect 45780 18284 46620 18340
rect 46676 18284 46686 18340
rect 3154 18172 3164 18228
rect 3220 18172 4508 18228
rect 4564 18172 4574 18228
rect 7522 18172 7532 18228
rect 7588 18172 8316 18228
rect 8372 18172 8382 18228
rect 15810 18172 15820 18228
rect 15876 18172 20076 18228
rect 20132 18172 20142 18228
rect 24210 18172 24220 18228
rect 24276 18172 27020 18228
rect 27076 18172 27356 18228
rect 27412 18172 27422 18228
rect 27804 18116 27860 18284
rect 36316 18228 36372 18284
rect 28018 18172 28028 18228
rect 28084 18172 29708 18228
rect 29764 18172 31052 18228
rect 31108 18172 31836 18228
rect 31892 18172 31902 18228
rect 34972 18172 36372 18228
rect 36530 18172 36540 18228
rect 36596 18172 37324 18228
rect 37380 18172 37390 18228
rect 42550 18172 42588 18228
rect 42644 18172 42654 18228
rect 1698 18060 1708 18116
rect 1764 18060 3500 18116
rect 3556 18060 3948 18116
rect 4004 18060 4014 18116
rect 17826 18060 17836 18116
rect 17892 18060 19068 18116
rect 19124 18060 19134 18116
rect 22306 18060 22316 18116
rect 22372 18060 27860 18116
rect 29260 18060 30380 18116
rect 30436 18060 30446 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 15698 17948 15708 18004
rect 15764 17948 17388 18004
rect 17444 17948 18508 18004
rect 18564 17948 18574 18004
rect 20178 17948 20188 18004
rect 20244 17948 21308 18004
rect 21364 17948 23212 18004
rect 23268 17948 23278 18004
rect 24546 17948 24556 18004
rect 24612 17948 26460 18004
rect 26516 17948 27804 18004
rect 27860 17948 27870 18004
rect 20188 17892 20244 17948
rect 29260 17892 29316 18060
rect 30380 18004 30436 18060
rect 34972 18004 35028 18172
rect 37622 18060 37660 18116
rect 37716 18060 37726 18116
rect 38966 18060 39004 18116
rect 39060 18060 39070 18116
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 30380 17948 35028 18004
rect 35532 17948 36204 18004
rect 36260 17948 38892 18004
rect 38948 17948 43372 18004
rect 43428 17948 43438 18004
rect 35532 17892 35588 17948
rect 16370 17836 16380 17892
rect 16436 17836 20244 17892
rect 23874 17836 23884 17892
rect 23940 17836 29316 17892
rect 29586 17836 29596 17892
rect 29652 17836 31276 17892
rect 31332 17836 31342 17892
rect 34066 17836 34076 17892
rect 34132 17836 35588 17892
rect 36082 17836 36092 17892
rect 36148 17836 39900 17892
rect 39956 17836 41132 17892
rect 41188 17836 41198 17892
rect 47842 17836 47852 17892
rect 47908 17836 48636 17892
rect 48692 17836 49196 17892
rect 49252 17836 49262 17892
rect 2482 17724 2492 17780
rect 2548 17724 4172 17780
rect 4228 17724 4620 17780
rect 4676 17724 4686 17780
rect 9650 17724 9660 17780
rect 9716 17724 10780 17780
rect 10836 17724 10846 17780
rect 11106 17724 11116 17780
rect 11172 17724 12908 17780
rect 12964 17724 13692 17780
rect 13748 17724 13758 17780
rect 16818 17724 16828 17780
rect 16884 17724 19404 17780
rect 19460 17724 19470 17780
rect 22194 17724 22204 17780
rect 22260 17724 23324 17780
rect 23380 17724 23390 17780
rect 24882 17724 24892 17780
rect 24948 17724 28140 17780
rect 28196 17724 28206 17780
rect 28354 17724 28364 17780
rect 28420 17724 28458 17780
rect 28578 17724 28588 17780
rect 28644 17724 30492 17780
rect 30548 17724 30558 17780
rect 31714 17724 31724 17780
rect 31780 17724 32844 17780
rect 32900 17724 32910 17780
rect 33058 17724 33068 17780
rect 33124 17724 33964 17780
rect 34020 17724 34030 17780
rect 6290 17612 6300 17668
rect 6356 17612 7756 17668
rect 7812 17612 7822 17668
rect 15362 17612 15372 17668
rect 15428 17612 16492 17668
rect 16548 17612 16558 17668
rect 20178 17612 20188 17668
rect 20244 17612 21756 17668
rect 21812 17612 22092 17668
rect 22148 17612 22158 17668
rect 24770 17612 24780 17668
rect 24836 17612 25228 17668
rect 25284 17612 25294 17668
rect 28242 17612 28252 17668
rect 28308 17612 29036 17668
rect 29092 17612 29102 17668
rect 32498 17612 32508 17668
rect 32564 17612 33516 17668
rect 33572 17612 35308 17668
rect 37202 17612 37212 17668
rect 37268 17612 38444 17668
rect 38500 17612 38510 17668
rect 38994 17612 39004 17668
rect 39060 17612 39788 17668
rect 39844 17612 39854 17668
rect 44706 17612 44716 17668
rect 44772 17612 46284 17668
rect 46340 17612 46350 17668
rect 21298 17500 21308 17556
rect 21364 17500 23436 17556
rect 23492 17500 23502 17556
rect 26898 17500 26908 17556
rect 26964 17500 27356 17556
rect 27412 17500 29148 17556
rect 29204 17500 29214 17556
rect 32274 17500 32284 17556
rect 32340 17500 33292 17556
rect 33348 17500 34300 17556
rect 34356 17500 34366 17556
rect 35252 17444 35308 17612
rect 35410 17500 35420 17556
rect 35476 17500 36316 17556
rect 36372 17500 36876 17556
rect 36932 17500 36942 17556
rect 38882 17500 38892 17556
rect 38948 17500 40572 17556
rect 40628 17500 40638 17556
rect 6514 17388 6524 17444
rect 6580 17388 8092 17444
rect 8148 17388 8158 17444
rect 9426 17388 9436 17444
rect 9492 17388 11228 17444
rect 11284 17388 11294 17444
rect 12898 17388 12908 17444
rect 12964 17388 14140 17444
rect 14196 17388 14206 17444
rect 18162 17388 18172 17444
rect 18228 17388 21532 17444
rect 21588 17388 21598 17444
rect 27794 17388 27804 17444
rect 27860 17388 28140 17444
rect 28196 17388 29260 17444
rect 29316 17388 29326 17444
rect 33506 17388 33516 17444
rect 33572 17388 34076 17444
rect 34132 17388 34412 17444
rect 34468 17388 34478 17444
rect 35252 17388 35644 17444
rect 35700 17388 35756 17444
rect 35812 17388 36428 17444
rect 36484 17388 36494 17444
rect 30258 17276 30268 17332
rect 30324 17276 35532 17332
rect 35588 17276 35868 17332
rect 35924 17276 35934 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 26226 17164 26236 17220
rect 26292 17164 26908 17220
rect 33394 17164 33404 17220
rect 33460 17164 37660 17220
rect 37716 17164 37996 17220
rect 38052 17164 38062 17220
rect 26852 17108 26908 17164
rect 38892 17108 38948 17500
rect 41234 17388 41244 17444
rect 41300 17388 44156 17444
rect 44212 17388 44222 17444
rect 45798 17388 45836 17444
rect 45892 17388 45902 17444
rect 18946 17052 18956 17108
rect 19012 17052 24444 17108
rect 24500 17052 24510 17108
rect 24658 17052 24668 17108
rect 24724 17052 25676 17108
rect 25732 17052 25742 17108
rect 26852 17052 38948 17108
rect 45826 17052 45836 17108
rect 45892 17052 46396 17108
rect 46452 17052 47964 17108
rect 48020 17052 48030 17108
rect 1810 16940 1820 16996
rect 1876 16940 2828 16996
rect 2884 16940 2894 16996
rect 20178 16940 20188 16996
rect 20244 16940 21700 16996
rect 27682 16940 27692 16996
rect 27748 16940 28364 16996
rect 28420 16940 28430 16996
rect 30258 16940 30268 16996
rect 30324 16940 30604 16996
rect 30660 16940 31332 16996
rect 33954 16940 33964 16996
rect 34020 16940 34188 16996
rect 34244 16940 35756 16996
rect 35812 16940 35822 16996
rect 36530 16940 36540 16996
rect 36596 16940 37548 16996
rect 37604 16940 38892 16996
rect 38948 16940 40908 16996
rect 40964 16940 40974 16996
rect 21644 16884 21700 16940
rect 31276 16884 31332 16940
rect 5842 16828 5852 16884
rect 5908 16828 6524 16884
rect 6580 16828 7196 16884
rect 7252 16828 7262 16884
rect 8530 16828 8540 16884
rect 8596 16828 9884 16884
rect 9940 16828 9950 16884
rect 16818 16828 16828 16884
rect 16884 16828 18172 16884
rect 18228 16828 18238 16884
rect 21634 16828 21644 16884
rect 21700 16828 23492 16884
rect 31266 16828 31276 16884
rect 31332 16828 31342 16884
rect 31490 16828 31500 16884
rect 31556 16828 33180 16884
rect 33236 16828 33246 16884
rect 34514 16828 34524 16884
rect 34580 16828 37884 16884
rect 37940 16828 37950 16884
rect 39442 16828 39452 16884
rect 39508 16828 40348 16884
rect 40404 16828 41468 16884
rect 41524 16828 44716 16884
rect 44772 16828 44782 16884
rect 23436 16772 23492 16828
rect 2594 16716 2604 16772
rect 2660 16716 3052 16772
rect 3108 16716 5964 16772
rect 6020 16716 7084 16772
rect 7140 16716 7150 16772
rect 19954 16716 19964 16772
rect 20020 16716 21532 16772
rect 21588 16716 21598 16772
rect 23436 16716 26684 16772
rect 26740 16716 27244 16772
rect 27300 16716 27310 16772
rect 28130 16716 28140 16772
rect 28196 16716 30156 16772
rect 30212 16716 31724 16772
rect 31780 16716 31790 16772
rect 35186 16716 35196 16772
rect 35252 16716 35262 16772
rect 37426 16716 37436 16772
rect 37492 16716 41020 16772
rect 41076 16716 41086 16772
rect 45938 16716 45948 16772
rect 46004 16716 47516 16772
rect 47572 16716 47582 16772
rect 35196 16660 35252 16716
rect 28018 16604 28028 16660
rect 28084 16604 33404 16660
rect 33460 16604 33470 16660
rect 35196 16604 38668 16660
rect 38770 16604 38780 16660
rect 38836 16604 41916 16660
rect 41972 16604 41982 16660
rect 44594 16604 44604 16660
rect 44660 16604 49084 16660
rect 49140 16604 49150 16660
rect 38612 16548 38668 16604
rect 9538 16492 9548 16548
rect 9604 16492 10108 16548
rect 10164 16492 12348 16548
rect 12404 16492 12796 16548
rect 12852 16492 12862 16548
rect 25778 16492 25788 16548
rect 25844 16492 29596 16548
rect 29652 16492 29662 16548
rect 38612 16492 39116 16548
rect 39172 16492 39182 16548
rect 44482 16492 44492 16548
rect 44548 16492 44940 16548
rect 44996 16492 47068 16548
rect 47124 16492 47134 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 30146 16380 30156 16436
rect 30212 16380 32284 16436
rect 32340 16380 32350 16436
rect 9874 16268 9884 16324
rect 9940 16268 10668 16324
rect 10724 16268 11228 16324
rect 11284 16268 12572 16324
rect 12628 16268 18844 16324
rect 18900 16268 26124 16324
rect 26180 16268 26190 16324
rect 7970 16156 7980 16212
rect 8036 16156 8932 16212
rect 17154 16156 17164 16212
rect 17220 16156 18620 16212
rect 18676 16156 18686 16212
rect 21186 16156 21196 16212
rect 21252 16156 22540 16212
rect 22596 16156 22606 16212
rect 27682 16156 27692 16212
rect 27748 16156 28476 16212
rect 28532 16156 28542 16212
rect 47058 16156 47068 16212
rect 47124 16156 48412 16212
rect 48468 16156 48478 16212
rect 8876 16100 8932 16156
rect 6402 16044 6412 16100
rect 6468 16044 8428 16100
rect 8866 16044 8876 16100
rect 8932 16044 8942 16100
rect 9314 16044 9324 16100
rect 9380 16044 9390 16100
rect 17266 16044 17276 16100
rect 17332 16044 17836 16100
rect 17892 16044 21532 16100
rect 21588 16044 21598 16100
rect 24546 16044 24556 16100
rect 24612 16044 27580 16100
rect 27636 16044 28252 16100
rect 28308 16044 28318 16100
rect 28578 16044 28588 16100
rect 28644 16044 31276 16100
rect 31332 16044 31342 16100
rect 36642 16044 36652 16100
rect 36708 16044 37324 16100
rect 37380 16044 37390 16100
rect 38658 16044 38668 16100
rect 38724 16044 38780 16100
rect 38836 16044 38846 16100
rect 8372 15988 8428 16044
rect 9324 15988 9380 16044
rect 2482 15932 2492 15988
rect 2548 15932 3388 15988
rect 3444 15932 3454 15988
rect 8372 15932 9380 15988
rect 11106 15932 11116 15988
rect 11172 15932 12684 15988
rect 12740 15932 12750 15988
rect 13010 15932 13020 15988
rect 13076 15932 13692 15988
rect 13748 15932 13758 15988
rect 15474 15932 15484 15988
rect 15540 15932 17612 15988
rect 17668 15932 22540 15988
rect 22596 15932 23548 15988
rect 23604 15932 23614 15988
rect 26450 15932 26460 15988
rect 26516 15932 27244 15988
rect 27300 15932 28028 15988
rect 28084 15932 28094 15988
rect 29922 15932 29932 15988
rect 29988 15932 30940 15988
rect 30996 15932 42924 15988
rect 42980 15932 43820 15988
rect 43876 15932 43886 15988
rect 8978 15820 8988 15876
rect 9044 15820 10556 15876
rect 10612 15820 10622 15876
rect 14466 15820 14476 15876
rect 14532 15820 15148 15876
rect 15204 15820 15214 15876
rect 19628 15820 22036 15876
rect 22194 15820 22204 15876
rect 22260 15820 35308 15876
rect 35364 15820 36988 15876
rect 37044 15820 37054 15876
rect 37398 15820 37436 15876
rect 37492 15820 37502 15876
rect 37986 15820 37996 15876
rect 38052 15820 38444 15876
rect 38500 15820 38510 15876
rect 38658 15820 38668 15876
rect 38724 15820 39564 15876
rect 39620 15820 39630 15876
rect 40338 15820 40348 15876
rect 40404 15820 45052 15876
rect 45108 15820 45118 15876
rect 19628 15764 19684 15820
rect 12114 15708 12124 15764
rect 12180 15708 12796 15764
rect 12852 15708 13804 15764
rect 13860 15708 14028 15764
rect 14084 15708 14812 15764
rect 14868 15708 19684 15764
rect 21980 15764 22036 15820
rect 21980 15708 39676 15764
rect 39732 15708 39742 15764
rect 19628 15652 19684 15708
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 19618 15596 19628 15652
rect 19684 15596 19694 15652
rect 36978 15596 36988 15652
rect 37044 15596 37324 15652
rect 37380 15596 38556 15652
rect 38612 15596 38622 15652
rect 2258 15484 2268 15540
rect 2324 15484 4172 15540
rect 4228 15484 4238 15540
rect 5954 15484 5964 15540
rect 6020 15484 6748 15540
rect 6804 15484 8260 15540
rect 8418 15484 8428 15540
rect 8484 15484 9884 15540
rect 9940 15484 9950 15540
rect 15026 15484 15036 15540
rect 15092 15484 17276 15540
rect 17332 15484 18396 15540
rect 18452 15484 19404 15540
rect 19460 15484 20524 15540
rect 20580 15484 20590 15540
rect 26114 15484 26124 15540
rect 26180 15484 26908 15540
rect 29922 15484 29932 15540
rect 29988 15484 30828 15540
rect 30884 15484 30894 15540
rect 32274 15484 32284 15540
rect 32340 15484 33852 15540
rect 33908 15484 33918 15540
rect 38882 15484 38892 15540
rect 38948 15484 39340 15540
rect 39396 15484 39406 15540
rect 8204 15428 8260 15484
rect 26852 15428 26908 15484
rect 2818 15372 2828 15428
rect 2884 15372 4620 15428
rect 4676 15372 5852 15428
rect 5908 15372 6972 15428
rect 7028 15372 7038 15428
rect 8194 15372 8204 15428
rect 8260 15372 8764 15428
rect 8820 15372 10892 15428
rect 10948 15372 10958 15428
rect 13356 15372 14252 15428
rect 14308 15372 14318 15428
rect 26852 15372 30604 15428
rect 30660 15372 30670 15428
rect 32050 15372 32060 15428
rect 32116 15372 32956 15428
rect 33012 15372 33022 15428
rect 38770 15372 38780 15428
rect 38836 15372 39228 15428
rect 39284 15372 39294 15428
rect 39890 15372 39900 15428
rect 39956 15372 41132 15428
rect 41188 15372 41198 15428
rect 13356 15316 13412 15372
rect 38780 15316 38836 15372
rect 3266 15260 3276 15316
rect 3332 15260 6748 15316
rect 6804 15260 6814 15316
rect 8372 15260 13412 15316
rect 13570 15260 13580 15316
rect 13636 15260 14476 15316
rect 14532 15260 14542 15316
rect 16818 15260 16828 15316
rect 16884 15260 18060 15316
rect 18116 15260 18732 15316
rect 18788 15260 18798 15316
rect 22306 15260 22316 15316
rect 22372 15260 27804 15316
rect 27860 15260 27870 15316
rect 29250 15260 29260 15316
rect 29316 15260 30828 15316
rect 30884 15260 30894 15316
rect 32722 15260 32732 15316
rect 32788 15260 33516 15316
rect 33572 15260 33582 15316
rect 38770 15260 38780 15316
rect 38836 15260 38846 15316
rect 39340 15260 39788 15316
rect 39844 15260 39854 15316
rect 40562 15260 40572 15316
rect 40628 15260 48860 15316
rect 48916 15260 48926 15316
rect 8372 15204 8428 15260
rect 39340 15204 39396 15260
rect 3826 15148 3836 15204
rect 3892 15148 4844 15204
rect 4900 15148 6188 15204
rect 6244 15148 6254 15204
rect 6514 15148 6524 15204
rect 6580 15148 8428 15204
rect 8866 15148 8876 15204
rect 8932 15148 10108 15204
rect 10164 15148 10174 15204
rect 14130 15148 14140 15204
rect 14196 15148 15820 15204
rect 15876 15148 15886 15204
rect 17938 15148 17948 15204
rect 18004 15148 22204 15204
rect 22260 15148 22270 15204
rect 30706 15148 30716 15204
rect 30772 15148 33068 15204
rect 33124 15148 33134 15204
rect 33842 15148 33852 15204
rect 33908 15148 34524 15204
rect 34580 15148 34590 15204
rect 39330 15148 39340 15204
rect 39396 15148 39406 15204
rect 17948 15092 18004 15148
rect 42018 15092 42028 15148
rect 42084 15092 42094 15148
rect 6850 15036 6860 15092
rect 6916 15036 8092 15092
rect 8148 15036 8158 15092
rect 11778 15036 11788 15092
rect 11844 15036 18004 15092
rect 20738 15036 20748 15092
rect 20804 15036 21084 15092
rect 21140 15036 21644 15092
rect 21700 15036 21710 15092
rect 31938 15036 31948 15092
rect 32004 15036 34188 15092
rect 34244 15036 34254 15092
rect 37650 15036 37660 15092
rect 37716 15036 39228 15092
rect 39284 15036 39294 15092
rect 41682 15036 41692 15092
rect 41748 15036 42084 15092
rect 9202 14924 9212 14980
rect 9268 14924 18956 14980
rect 19012 14924 19022 14980
rect 20402 14924 20412 14980
rect 20468 14924 31948 14980
rect 32498 14924 32508 14980
rect 32564 14924 33516 14980
rect 33572 14924 33582 14980
rect 38546 14924 38556 14980
rect 38612 14924 40796 14980
rect 40852 14924 40862 14980
rect 44818 14924 44828 14980
rect 44884 14924 46060 14980
rect 46116 14924 46126 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 4834 14812 4844 14868
rect 4900 14812 5740 14868
rect 5796 14812 7084 14868
rect 7140 14812 7150 14868
rect 17938 14812 17948 14868
rect 18004 14812 26348 14868
rect 26404 14812 26414 14868
rect 3602 14700 3612 14756
rect 3668 14700 6860 14756
rect 6916 14700 6926 14756
rect 31892 14644 31948 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 50200 14868 51000 14896
rect 36642 14812 36652 14868
rect 36708 14812 39004 14868
rect 39060 14812 39070 14868
rect 49074 14812 49084 14868
rect 49140 14812 51000 14868
rect 50200 14784 51000 14812
rect 33506 14700 33516 14756
rect 33572 14700 35532 14756
rect 35588 14700 35598 14756
rect 9538 14588 9548 14644
rect 9604 14588 12908 14644
rect 12964 14588 12974 14644
rect 14130 14588 14140 14644
rect 14196 14588 29932 14644
rect 29988 14588 29998 14644
rect 31892 14588 34132 14644
rect 34290 14588 34300 14644
rect 34356 14588 38108 14644
rect 38164 14588 38174 14644
rect 41346 14588 41356 14644
rect 41412 14588 42252 14644
rect 42308 14588 42318 14644
rect 47730 14588 47740 14644
rect 47796 14588 49196 14644
rect 49252 14588 49262 14644
rect 34076 14532 34132 14588
rect 8082 14476 8092 14532
rect 8148 14476 9436 14532
rect 9492 14476 12460 14532
rect 12516 14476 12526 14532
rect 29362 14476 29372 14532
rect 29428 14476 30156 14532
rect 30212 14476 32732 14532
rect 32788 14476 32798 14532
rect 34076 14476 35308 14532
rect 35364 14476 35868 14532
rect 35924 14476 35934 14532
rect 37538 14476 37548 14532
rect 37604 14476 37660 14532
rect 37716 14476 37726 14532
rect 38546 14476 38556 14532
rect 38612 14476 39004 14532
rect 39060 14476 39070 14532
rect 45378 14476 45388 14532
rect 45444 14476 46732 14532
rect 46788 14476 46798 14532
rect 21634 14364 21644 14420
rect 21700 14364 23660 14420
rect 23716 14364 23726 14420
rect 37202 14364 37212 14420
rect 37268 14364 38892 14420
rect 38948 14364 38958 14420
rect 39554 14364 39564 14420
rect 39620 14364 40236 14420
rect 40292 14364 40302 14420
rect 38892 14308 38948 14364
rect 2930 14252 2940 14308
rect 2996 14252 5628 14308
rect 5684 14252 5694 14308
rect 9762 14252 9772 14308
rect 9828 14252 10556 14308
rect 10612 14252 10622 14308
rect 18162 14252 18172 14308
rect 18228 14252 19516 14308
rect 19572 14252 19582 14308
rect 38892 14252 39788 14308
rect 39844 14252 39854 14308
rect 40002 14252 40012 14308
rect 40068 14252 40460 14308
rect 40516 14252 40526 14308
rect 45798 14252 45836 14308
rect 45892 14252 45902 14308
rect 8082 14140 8092 14196
rect 8148 14140 11116 14196
rect 11172 14140 12124 14196
rect 12180 14140 12190 14196
rect 32722 14140 32732 14196
rect 32788 14140 40348 14196
rect 40404 14140 40414 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 5516 14028 6300 14084
rect 6356 14028 7196 14084
rect 7252 14028 7262 14084
rect 8306 14028 8316 14084
rect 8372 14028 8876 14084
rect 8932 14028 11956 14084
rect 31714 14028 31724 14084
rect 31780 14028 34636 14084
rect 34692 14028 34702 14084
rect 5516 13972 5572 14028
rect 11900 13972 11956 14028
rect 3154 13916 3164 13972
rect 3220 13916 5516 13972
rect 5572 13916 5582 13972
rect 5954 13916 5964 13972
rect 6020 13916 6748 13972
rect 6804 13916 9996 13972
rect 10052 13916 10062 13972
rect 11890 13916 11900 13972
rect 11956 13916 12684 13972
rect 12740 13916 12750 13972
rect 22642 13916 22652 13972
rect 22708 13916 23996 13972
rect 24052 13916 24062 13972
rect 24434 13916 24444 13972
rect 24500 13916 26572 13972
rect 26628 13916 26638 13972
rect 32610 13916 32620 13972
rect 32676 13916 34412 13972
rect 34468 13916 34478 13972
rect 40338 13916 40348 13972
rect 40404 13916 41020 13972
rect 41076 13916 41086 13972
rect 41234 13916 41244 13972
rect 41300 13916 42140 13972
rect 42196 13916 42206 13972
rect 42802 13916 42812 13972
rect 42868 13916 46732 13972
rect 46788 13916 46798 13972
rect 2482 13804 2492 13860
rect 2548 13804 4396 13860
rect 4452 13804 4462 13860
rect 10322 13804 10332 13860
rect 10388 13804 11564 13860
rect 11620 13804 11630 13860
rect 31826 13804 31836 13860
rect 31892 13804 33740 13860
rect 33796 13804 33806 13860
rect 39666 13804 39676 13860
rect 39732 13804 41468 13860
rect 41524 13804 41534 13860
rect 42018 13804 42028 13860
rect 42084 13804 42364 13860
rect 42420 13804 42430 13860
rect 44482 13804 44492 13860
rect 44548 13804 48860 13860
rect 48916 13804 48926 13860
rect 3826 13692 3836 13748
rect 3892 13692 4620 13748
rect 4676 13692 4686 13748
rect 7970 13692 7980 13748
rect 8036 13692 10892 13748
rect 10948 13692 10958 13748
rect 16034 13692 16044 13748
rect 16100 13692 17612 13748
rect 17668 13692 18060 13748
rect 18116 13692 18126 13748
rect 19282 13692 19292 13748
rect 19348 13692 22764 13748
rect 22820 13692 22830 13748
rect 23762 13692 23772 13748
rect 23828 13692 27020 13748
rect 27076 13692 27086 13748
rect 27682 13692 27692 13748
rect 27748 13692 28252 13748
rect 28308 13692 28812 13748
rect 28868 13692 31500 13748
rect 31556 13692 32508 13748
rect 32564 13692 32732 13748
rect 32788 13692 32798 13748
rect 33030 13692 33068 13748
rect 33124 13692 33134 13748
rect 40226 13692 40236 13748
rect 40292 13692 41356 13748
rect 41412 13692 41422 13748
rect 46946 13692 46956 13748
rect 47012 13692 48076 13748
rect 48132 13692 48142 13748
rect 23772 13636 23828 13692
rect 3714 13580 3724 13636
rect 3780 13580 6636 13636
rect 6692 13580 6702 13636
rect 16594 13580 16604 13636
rect 16660 13580 17500 13636
rect 17556 13580 17566 13636
rect 18946 13580 18956 13636
rect 19012 13580 19628 13636
rect 19684 13580 19694 13636
rect 20738 13580 20748 13636
rect 20804 13580 21756 13636
rect 21812 13580 23828 13636
rect 26562 13580 26572 13636
rect 26628 13580 27356 13636
rect 27412 13580 27422 13636
rect 29922 13580 29932 13636
rect 29988 13580 34748 13636
rect 34804 13580 34814 13636
rect 43474 13580 43484 13636
rect 43540 13580 44268 13636
rect 44324 13580 44828 13636
rect 44884 13580 44894 13636
rect 15922 13468 15932 13524
rect 15988 13468 16268 13524
rect 16324 13468 17276 13524
rect 17332 13468 18620 13524
rect 18676 13468 18686 13524
rect 31378 13468 31388 13524
rect 31444 13468 33516 13524
rect 33572 13468 33582 13524
rect 41794 13468 41804 13524
rect 41860 13468 42588 13524
rect 42644 13468 42654 13524
rect 42802 13468 42812 13524
rect 42868 13468 42878 13524
rect 44146 13468 44156 13524
rect 44212 13468 44940 13524
rect 44996 13468 45006 13524
rect 47954 13468 47964 13524
rect 48020 13468 48524 13524
rect 48580 13468 48590 13524
rect 42812 13412 42868 13468
rect 6962 13356 6972 13412
rect 7028 13356 7644 13412
rect 7700 13356 12124 13412
rect 12180 13356 12190 13412
rect 12338 13356 12348 13412
rect 12404 13356 14028 13412
rect 14084 13356 26740 13412
rect 27458 13356 27468 13412
rect 27524 13356 29484 13412
rect 29540 13356 29550 13412
rect 31826 13356 31836 13412
rect 31892 13356 34972 13412
rect 35028 13356 35038 13412
rect 36082 13356 36092 13412
rect 36148 13356 37324 13412
rect 37380 13356 37390 13412
rect 42812 13356 43708 13412
rect 43764 13356 43774 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 26684 13300 26740 13356
rect 29484 13300 29540 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 11106 13244 11116 13300
rect 11172 13244 21084 13300
rect 21140 13244 21150 13300
rect 26684 13244 28028 13300
rect 28084 13244 28094 13300
rect 29484 13244 33292 13300
rect 33348 13244 33358 13300
rect 39106 13244 39116 13300
rect 39172 13244 41580 13300
rect 41636 13244 42700 13300
rect 42756 13244 42766 13300
rect 3266 13132 3276 13188
rect 3332 13132 4620 13188
rect 4676 13132 4686 13188
rect 18722 13132 18732 13188
rect 18788 13132 26460 13188
rect 26516 13132 27804 13188
rect 27860 13132 27870 13188
rect 28140 13132 34860 13188
rect 34916 13132 37548 13188
rect 37604 13132 37614 13188
rect 45490 13132 45500 13188
rect 45556 13132 46844 13188
rect 46900 13132 46910 13188
rect 2482 13020 2492 13076
rect 2548 13020 5964 13076
rect 6020 13020 6030 13076
rect 11890 13020 11900 13076
rect 11956 13020 12348 13076
rect 12404 13020 12414 13076
rect 19730 13020 19740 13076
rect 19796 13020 20636 13076
rect 20692 13020 20702 13076
rect 28140 12964 28196 13132
rect 28354 13020 28364 13076
rect 28420 13020 30380 13076
rect 30436 13020 31612 13076
rect 31668 13020 31678 13076
rect 36530 13020 36540 13076
rect 36596 13020 37324 13076
rect 37380 13020 37390 13076
rect 42326 13020 42364 13076
rect 42420 13020 42430 13076
rect 45154 13020 45164 13076
rect 45220 13020 47852 13076
rect 47908 13020 48300 13076
rect 48356 13020 48366 13076
rect 4498 12908 4508 12964
rect 4564 12908 4956 12964
rect 5012 12908 5628 12964
rect 5684 12908 5694 12964
rect 11666 12908 11676 12964
rect 11732 12908 12460 12964
rect 12516 12908 12526 12964
rect 13234 12908 13244 12964
rect 13300 12908 14364 12964
rect 14420 12908 14430 12964
rect 16370 12908 16380 12964
rect 16436 12908 16828 12964
rect 16884 12908 16894 12964
rect 22754 12908 22764 12964
rect 22820 12908 28196 12964
rect 29922 12908 29932 12964
rect 29988 12908 31052 12964
rect 31108 12908 31118 12964
rect 33282 12908 33292 12964
rect 33348 12908 36316 12964
rect 36372 12908 36382 12964
rect 38658 12908 38668 12964
rect 38724 12908 38762 12964
rect 46050 12908 46060 12964
rect 46116 12908 47964 12964
rect 48020 12908 48030 12964
rect 12898 12796 12908 12852
rect 12964 12796 13692 12852
rect 13748 12796 13758 12852
rect 17714 12796 17724 12852
rect 17780 12796 20412 12852
rect 20468 12796 20478 12852
rect 21970 12796 21980 12852
rect 22036 12796 22876 12852
rect 22932 12796 22942 12852
rect 23202 12796 23212 12852
rect 23268 12796 24668 12852
rect 24724 12796 24734 12852
rect 28018 12796 28028 12852
rect 28084 12796 33404 12852
rect 33460 12796 34300 12852
rect 34356 12796 34366 12852
rect 38994 12796 39004 12852
rect 39060 12796 42028 12852
rect 42084 12796 42094 12852
rect 43586 12796 43596 12852
rect 43652 12796 44044 12852
rect 44100 12796 49084 12852
rect 49140 12796 49150 12852
rect 4834 12684 4844 12740
rect 4900 12684 6636 12740
rect 6692 12684 6702 12740
rect 19506 12684 19516 12740
rect 19572 12684 21644 12740
rect 21700 12684 22652 12740
rect 22708 12684 22718 12740
rect 38210 12684 38220 12740
rect 38276 12684 40012 12740
rect 40068 12684 40078 12740
rect 41906 12684 41916 12740
rect 41972 12684 42476 12740
rect 42532 12684 42542 12740
rect 46162 12684 46172 12740
rect 46228 12684 47068 12740
rect 47124 12684 47134 12740
rect 5170 12572 5180 12628
rect 5236 12572 14140 12628
rect 14196 12572 14206 12628
rect 23090 12572 23100 12628
rect 23156 12572 24444 12628
rect 24500 12572 25452 12628
rect 25508 12572 25518 12628
rect 31892 12572 36428 12628
rect 36484 12572 36494 12628
rect 41234 12572 41244 12628
rect 41300 12572 45388 12628
rect 45444 12572 45454 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 31892 12516 31948 12572
rect 21074 12460 21084 12516
rect 21140 12460 31948 12516
rect 45154 12460 45164 12516
rect 45220 12460 46508 12516
rect 46564 12460 49644 12516
rect 49700 12460 49710 12516
rect 3490 12348 3500 12404
rect 3556 12348 5068 12404
rect 5124 12348 5134 12404
rect 7634 12348 7644 12404
rect 7700 12348 9772 12404
rect 9828 12348 9838 12404
rect 16370 12348 16380 12404
rect 16436 12348 39116 12404
rect 39172 12348 42588 12404
rect 42644 12348 42654 12404
rect 42802 12348 42812 12404
rect 42868 12348 43372 12404
rect 43428 12348 43438 12404
rect 46274 12348 46284 12404
rect 46340 12348 47516 12404
rect 47572 12348 48748 12404
rect 48804 12348 48814 12404
rect 24658 12236 24668 12292
rect 24724 12236 26180 12292
rect 26786 12236 26796 12292
rect 26852 12236 27916 12292
rect 27972 12236 30156 12292
rect 30212 12236 30222 12292
rect 31042 12236 31052 12292
rect 31108 12236 32396 12292
rect 32452 12236 32462 12292
rect 42690 12236 42700 12292
rect 42756 12236 43260 12292
rect 43316 12236 43326 12292
rect 47730 12236 47740 12292
rect 47796 12236 49196 12292
rect 49252 12236 49262 12292
rect 26124 12180 26180 12236
rect 14466 12124 14476 12180
rect 14532 12124 16716 12180
rect 16772 12124 17388 12180
rect 17444 12124 17454 12180
rect 26114 12124 26124 12180
rect 26180 12124 26908 12180
rect 26964 12124 26974 12180
rect 29698 12124 29708 12180
rect 29764 12124 31948 12180
rect 32004 12124 32844 12180
rect 32900 12124 35756 12180
rect 35812 12124 35822 12180
rect 37090 12124 37100 12180
rect 37156 12124 38948 12180
rect 39554 12124 39564 12180
rect 39620 12124 41244 12180
rect 41300 12124 41310 12180
rect 41458 12124 41468 12180
rect 41524 12124 43484 12180
rect 43540 12124 43550 12180
rect 45826 12124 45836 12180
rect 45892 12124 49084 12180
rect 49140 12124 49420 12180
rect 49476 12124 49486 12180
rect 2482 12012 2492 12068
rect 2548 12012 4060 12068
rect 4116 12012 4126 12068
rect 14130 12012 14140 12068
rect 14196 12012 14700 12068
rect 14756 12012 14766 12068
rect 18834 12012 18844 12068
rect 18900 12012 22428 12068
rect 22484 12012 22494 12068
rect 24658 12012 24668 12068
rect 24724 12012 25564 12068
rect 25620 12012 25630 12068
rect 38892 11956 38948 12124
rect 39106 12012 39116 12068
rect 39172 12012 41020 12068
rect 41076 12012 42924 12068
rect 42980 12012 42990 12068
rect 45938 12012 45948 12068
rect 46004 12012 47068 12068
rect 47124 12012 47134 12068
rect 5506 11900 5516 11956
rect 5572 11900 7196 11956
rect 7252 11900 7262 11956
rect 18386 11900 18396 11956
rect 18452 11900 19068 11956
rect 19124 11900 19134 11956
rect 38882 11900 38892 11956
rect 38948 11900 38958 11956
rect 42466 11900 42476 11956
rect 42532 11900 43708 11956
rect 43764 11900 44268 11956
rect 44324 11900 44334 11956
rect 20402 11788 20412 11844
rect 20468 11788 22092 11844
rect 22148 11788 22158 11844
rect 30268 11788 31668 11844
rect 31826 11788 31836 11844
rect 31892 11788 32228 11844
rect 37314 11788 37324 11844
rect 37380 11788 37390 11844
rect 39554 11788 39564 11844
rect 39620 11788 39788 11844
rect 39844 11788 41692 11844
rect 41748 11788 43484 11844
rect 43540 11788 43550 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 30268 11732 30324 11788
rect 31612 11732 31668 11788
rect 32172 11732 32228 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 9090 11676 9100 11732
rect 9156 11676 9996 11732
rect 10052 11676 16380 11732
rect 16436 11676 16446 11732
rect 20850 11676 20860 11732
rect 20916 11676 23324 11732
rect 23380 11676 23996 11732
rect 24052 11676 25228 11732
rect 25284 11676 25294 11732
rect 29250 11676 29260 11732
rect 29316 11676 29326 11732
rect 29474 11676 29484 11732
rect 29540 11676 30044 11732
rect 30100 11676 30110 11732
rect 30258 11676 30268 11732
rect 30324 11676 30334 11732
rect 31612 11676 31948 11732
rect 32004 11676 32014 11732
rect 32172 11676 32508 11732
rect 32564 11676 33964 11732
rect 34020 11676 34030 11732
rect 29260 11620 29316 11676
rect 37324 11620 37380 11788
rect 43138 11676 43148 11732
rect 43204 11676 44716 11732
rect 44772 11676 44782 11732
rect 47618 11676 47628 11732
rect 47684 11676 49084 11732
rect 49140 11676 49150 11732
rect 16930 11564 16940 11620
rect 16996 11564 25340 11620
rect 25396 11564 25788 11620
rect 25844 11564 25854 11620
rect 29260 11564 31724 11620
rect 31780 11564 31790 11620
rect 32274 11564 32284 11620
rect 32340 11564 37380 11620
rect 43586 11564 43596 11620
rect 43652 11564 44268 11620
rect 44324 11564 44334 11620
rect 47954 11564 47964 11620
rect 48020 11564 48748 11620
rect 48804 11564 48814 11620
rect 1810 11452 1820 11508
rect 1876 11452 5292 11508
rect 5348 11452 8764 11508
rect 8820 11452 8830 11508
rect 12786 11452 12796 11508
rect 12852 11452 13804 11508
rect 13860 11452 13870 11508
rect 18274 11452 18284 11508
rect 18340 11452 19180 11508
rect 19236 11452 19246 11508
rect 29362 11452 29372 11508
rect 29428 11452 30940 11508
rect 30996 11452 31006 11508
rect 31612 11452 37156 11508
rect 19954 11340 19964 11396
rect 20020 11340 20300 11396
rect 20356 11340 20366 11396
rect 28578 11340 28588 11396
rect 28644 11340 31276 11396
rect 31332 11340 31342 11396
rect 11554 11228 11564 11284
rect 11620 11228 12572 11284
rect 12628 11228 12638 11284
rect 19618 11228 19628 11284
rect 19684 11228 20860 11284
rect 20916 11228 20926 11284
rect 21634 11228 21644 11284
rect 21700 11228 22988 11284
rect 23044 11228 23054 11284
rect 29810 11228 29820 11284
rect 29876 11228 31388 11284
rect 31444 11228 31454 11284
rect 31612 11172 31668 11452
rect 37100 11396 37156 11452
rect 37324 11396 37380 11564
rect 37090 11340 37100 11396
rect 37156 11340 37166 11396
rect 37314 11340 37324 11396
rect 37380 11340 37390 11396
rect 37538 11340 37548 11396
rect 37604 11340 38332 11396
rect 38388 11340 38398 11396
rect 47282 11340 47292 11396
rect 47348 11340 49196 11396
rect 49252 11340 49262 11396
rect 37548 11284 37604 11340
rect 31826 11228 31836 11284
rect 31892 11228 33068 11284
rect 33124 11228 33134 11284
rect 35746 11228 35756 11284
rect 35812 11228 37604 11284
rect 15250 11116 15260 11172
rect 15316 11116 22036 11172
rect 26450 11116 26460 11172
rect 26516 11116 27468 11172
rect 27524 11116 28028 11172
rect 28084 11116 28812 11172
rect 28868 11116 28878 11172
rect 30034 11116 30044 11172
rect 30100 11116 31668 11172
rect 31826 11116 31836 11172
rect 31892 11116 32508 11172
rect 32564 11116 32574 11172
rect 21980 11060 22036 11116
rect 21970 11004 21980 11060
rect 22036 11004 33404 11060
rect 33460 11004 35532 11060
rect 35588 11004 36988 11060
rect 37044 11004 37054 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 38612 10948 38668 11284
rect 38724 11228 38734 11284
rect 43026 11228 43036 11284
rect 43092 11228 43484 11284
rect 43540 11228 43550 11284
rect 43810 11228 43820 11284
rect 43876 11228 45388 11284
rect 45444 11228 45454 11284
rect 10994 10892 11004 10948
rect 11060 10892 14476 10948
rect 14532 10892 14542 10948
rect 25778 10892 25788 10948
rect 25844 10892 31836 10948
rect 31892 10892 31902 10948
rect 36418 10892 36428 10948
rect 36484 10892 37548 10948
rect 37604 10892 38108 10948
rect 38164 10892 38668 10948
rect 4274 10780 4284 10836
rect 4340 10780 5516 10836
rect 5572 10780 5582 10836
rect 5730 10780 5740 10836
rect 5796 10780 6412 10836
rect 6468 10780 6478 10836
rect 15026 10780 15036 10836
rect 15092 10780 16716 10836
rect 16772 10780 16782 10836
rect 20962 10780 20972 10836
rect 21028 10780 25116 10836
rect 25172 10780 25182 10836
rect 28914 10780 28924 10836
rect 28980 10780 31724 10836
rect 31780 10780 31790 10836
rect 31892 10780 48076 10836
rect 48132 10780 48142 10836
rect 31892 10724 31948 10780
rect 29138 10668 29148 10724
rect 29204 10668 30044 10724
rect 30100 10668 30110 10724
rect 30380 10668 31948 10724
rect 34066 10668 34076 10724
rect 34132 10668 34972 10724
rect 35028 10668 36652 10724
rect 36708 10668 36718 10724
rect 41234 10668 41244 10724
rect 41300 10668 42924 10724
rect 42980 10668 44044 10724
rect 44100 10668 44110 10724
rect 44594 10668 44604 10724
rect 44660 10668 46732 10724
rect 46788 10668 46798 10724
rect 10546 10556 10556 10612
rect 10612 10556 11228 10612
rect 11284 10556 13580 10612
rect 13636 10556 13646 10612
rect 13906 10556 13916 10612
rect 13972 10556 15372 10612
rect 15428 10556 16156 10612
rect 16212 10556 16222 10612
rect 17714 10556 17724 10612
rect 17780 10556 21308 10612
rect 21364 10556 23548 10612
rect 23604 10556 23614 10612
rect 28354 10556 28364 10612
rect 28420 10556 29372 10612
rect 29428 10556 29438 10612
rect 9762 10444 9772 10500
rect 9828 10444 13020 10500
rect 13076 10444 13692 10500
rect 13748 10444 13758 10500
rect 14802 10444 14812 10500
rect 14868 10444 15932 10500
rect 15988 10444 16604 10500
rect 16660 10444 16670 10500
rect 26674 10444 26684 10500
rect 26740 10444 27244 10500
rect 27300 10444 28140 10500
rect 28196 10444 28206 10500
rect 9426 10332 9436 10388
rect 9492 10332 11900 10388
rect 11956 10332 11966 10388
rect 25778 10220 25788 10276
rect 25844 10220 27356 10276
rect 27412 10220 27422 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 8194 10108 8204 10164
rect 8260 10108 24668 10164
rect 24724 10108 27804 10164
rect 27860 10108 29148 10164
rect 29204 10108 29214 10164
rect 30380 10052 30436 10668
rect 48076 10612 48132 10780
rect 48962 10668 48972 10724
rect 49028 10668 49644 10724
rect 49700 10668 49710 10724
rect 50200 10612 51000 10640
rect 31378 10556 31388 10612
rect 31444 10556 32172 10612
rect 32228 10556 32238 10612
rect 34402 10556 34412 10612
rect 34468 10556 35084 10612
rect 35140 10556 36316 10612
rect 36372 10556 36382 10612
rect 45378 10556 45388 10612
rect 45444 10556 46060 10612
rect 46116 10556 46126 10612
rect 48076 10556 51000 10612
rect 50200 10528 51000 10556
rect 41906 10444 41916 10500
rect 41972 10444 42588 10500
rect 42644 10444 43708 10500
rect 43764 10444 43774 10500
rect 46946 10444 46956 10500
rect 47012 10444 48524 10500
rect 48580 10444 48590 10500
rect 40338 10332 40348 10388
rect 40404 10332 41468 10388
rect 41524 10332 43372 10388
rect 43428 10332 43438 10388
rect 45266 10332 45276 10388
rect 45332 10332 46844 10388
rect 46900 10332 46910 10388
rect 47068 10332 47628 10388
rect 47684 10332 47694 10388
rect 47068 10276 47124 10332
rect 41234 10220 41244 10276
rect 41300 10220 47124 10276
rect 47282 10220 47292 10276
rect 47348 10220 49532 10276
rect 49588 10220 49598 10276
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 32162 10108 32172 10164
rect 32228 10108 34188 10164
rect 34244 10108 34254 10164
rect 37202 10108 37212 10164
rect 37268 10108 38332 10164
rect 38388 10108 38398 10164
rect 41794 10108 41804 10164
rect 41860 10108 44492 10164
rect 44548 10108 44558 10164
rect 5842 9996 5852 10052
rect 5908 9996 7644 10052
rect 7700 9996 8260 10052
rect 16034 9996 16044 10052
rect 16100 9996 18284 10052
rect 18340 9996 18350 10052
rect 18834 9996 18844 10052
rect 18900 9996 20300 10052
rect 20356 9996 20366 10052
rect 26012 9996 30436 10052
rect 38210 9996 38220 10052
rect 38276 9996 39340 10052
rect 39396 9996 39406 10052
rect 42018 9996 42028 10052
rect 42084 9996 42588 10052
rect 42644 9996 42654 10052
rect 8204 9940 8260 9996
rect 26012 9940 26068 9996
rect 8194 9884 8204 9940
rect 8260 9884 8270 9940
rect 11330 9884 11340 9940
rect 11396 9884 11564 9940
rect 11620 9884 12460 9940
rect 12516 9884 12526 9940
rect 12684 9884 26068 9940
rect 27458 9884 27468 9940
rect 27524 9884 33516 9940
rect 33572 9884 33582 9940
rect 34514 9884 34524 9940
rect 34580 9884 35644 9940
rect 35700 9884 35710 9940
rect 37090 9884 37100 9940
rect 37156 9884 38668 9940
rect 38724 9884 38734 9940
rect 41122 9884 41132 9940
rect 41188 9884 41692 9940
rect 41748 9884 44828 9940
rect 44884 9884 44894 9940
rect 47058 9884 47068 9940
rect 47124 9884 48860 9940
rect 48916 9884 48926 9940
rect 12684 9828 12740 9884
rect 33516 9828 33572 9884
rect 4722 9772 4732 9828
rect 4788 9772 12740 9828
rect 12898 9772 12908 9828
rect 12964 9772 15596 9828
rect 15652 9772 16940 9828
rect 16996 9772 17006 9828
rect 21970 9772 21980 9828
rect 22036 9772 22652 9828
rect 22708 9772 22718 9828
rect 22866 9772 22876 9828
rect 22932 9772 23604 9828
rect 28466 9772 28476 9828
rect 28532 9772 30940 9828
rect 30996 9772 31006 9828
rect 33516 9772 36428 9828
rect 36484 9772 37884 9828
rect 37940 9772 37950 9828
rect 42018 9772 42028 9828
rect 42084 9772 44604 9828
rect 44660 9772 45052 9828
rect 45108 9772 45118 9828
rect 23548 9716 23604 9772
rect 5170 9660 5180 9716
rect 5236 9660 7700 9716
rect 19506 9660 19516 9716
rect 19572 9660 21644 9716
rect 21700 9660 23212 9716
rect 23268 9660 23278 9716
rect 23538 9660 23548 9716
rect 23604 9660 28140 9716
rect 28196 9660 29372 9716
rect 29428 9660 29438 9716
rect 32722 9660 32732 9716
rect 32788 9660 33516 9716
rect 33572 9660 33582 9716
rect 38994 9660 39004 9716
rect 39060 9660 39788 9716
rect 39844 9660 39854 9716
rect 7644 9604 7700 9660
rect 5954 9548 5964 9604
rect 6020 9548 7196 9604
rect 7252 9548 7262 9604
rect 7634 9548 7644 9604
rect 7700 9548 8092 9604
rect 8148 9548 8158 9604
rect 8306 9548 8316 9604
rect 8372 9548 11004 9604
rect 11060 9548 11070 9604
rect 11666 9548 11676 9604
rect 11732 9548 12236 9604
rect 12292 9548 18284 9604
rect 18340 9548 20636 9604
rect 20692 9548 20702 9604
rect 22642 9548 22652 9604
rect 22708 9548 23772 9604
rect 23828 9548 23838 9604
rect 40450 9548 40460 9604
rect 40516 9548 45836 9604
rect 45892 9548 45902 9604
rect 13682 9436 13692 9492
rect 13748 9436 16324 9492
rect 20178 9436 20188 9492
rect 20244 9436 22428 9492
rect 22484 9436 22494 9492
rect 38770 9436 38780 9492
rect 38836 9436 42476 9492
rect 42532 9436 42542 9492
rect 8530 9324 8540 9380
rect 8596 9324 12012 9380
rect 12068 9324 12078 9380
rect 16268 9268 16324 9436
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 22866 9324 22876 9380
rect 22932 9324 24108 9380
rect 24164 9324 29372 9380
rect 29428 9324 41356 9380
rect 41412 9324 42140 9380
rect 42196 9324 42206 9380
rect 47842 9324 47852 9380
rect 47908 9324 49084 9380
rect 49140 9324 49150 9380
rect 8978 9212 8988 9268
rect 9044 9212 10780 9268
rect 10836 9212 14364 9268
rect 14420 9212 16044 9268
rect 16100 9212 16110 9268
rect 16268 9212 21308 9268
rect 21364 9212 22316 9268
rect 22372 9212 22382 9268
rect 24434 9212 24444 9268
rect 24500 9212 25564 9268
rect 25620 9212 25630 9268
rect 27122 9212 27132 9268
rect 27188 9212 31500 9268
rect 31556 9212 31566 9268
rect 42466 9212 42476 9268
rect 42532 9212 46508 9268
rect 46564 9212 46574 9268
rect 14466 9100 14476 9156
rect 14532 9100 17164 9156
rect 17220 9100 17230 9156
rect 20626 9100 20636 9156
rect 20692 9100 23212 9156
rect 23268 9100 23278 9156
rect 25330 9100 25340 9156
rect 25396 9100 25900 9156
rect 25956 9100 25966 9156
rect 31042 9100 31052 9156
rect 31108 9100 31948 9156
rect 33842 9100 33852 9156
rect 33908 9100 34524 9156
rect 34580 9100 34590 9156
rect 46386 9100 46396 9156
rect 46452 9100 48076 9156
rect 48132 9100 48748 9156
rect 48804 9100 48814 9156
rect 31892 9044 31948 9100
rect 22530 8988 22540 9044
rect 22596 8988 24780 9044
rect 24836 8988 24846 9044
rect 28914 8988 28924 9044
rect 28980 8988 29820 9044
rect 29876 8988 29886 9044
rect 30034 8988 30044 9044
rect 30100 8988 30716 9044
rect 30772 8988 30782 9044
rect 31892 8988 41468 9044
rect 41524 8988 41534 9044
rect 47058 8988 47068 9044
rect 47124 8988 47852 9044
rect 47908 8988 49196 9044
rect 49252 8988 49262 9044
rect 10434 8876 10444 8932
rect 10500 8876 15036 8932
rect 15092 8876 15102 8932
rect 20066 8876 20076 8932
rect 20132 8820 20188 8932
rect 20738 8876 20748 8932
rect 20804 8876 23660 8932
rect 23716 8876 23726 8932
rect 38434 8876 38444 8932
rect 38500 8876 38892 8932
rect 38948 8876 38958 8932
rect 42550 8876 42588 8932
rect 42644 8876 42654 8932
rect 45938 8876 45948 8932
rect 46004 8876 48748 8932
rect 48804 8876 48814 8932
rect 9874 8764 9884 8820
rect 9940 8764 11900 8820
rect 11956 8764 11966 8820
rect 20132 8764 22652 8820
rect 22708 8764 23548 8820
rect 23604 8764 23614 8820
rect 24434 8764 24444 8820
rect 24500 8764 24510 8820
rect 28578 8764 28588 8820
rect 28644 8764 29148 8820
rect 29204 8764 30156 8820
rect 30212 8764 30222 8820
rect 31490 8764 31500 8820
rect 31556 8764 32396 8820
rect 32452 8764 32462 8820
rect 45490 8764 45500 8820
rect 45556 8764 46844 8820
rect 46900 8764 47628 8820
rect 47684 8764 47694 8820
rect 24444 8708 24500 8764
rect 6626 8652 6636 8708
rect 6692 8652 6702 8708
rect 21970 8652 21980 8708
rect 22036 8652 23324 8708
rect 23380 8652 23390 8708
rect 23538 8652 23548 8708
rect 23604 8652 24500 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 6636 8596 6692 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 5170 8540 5180 8596
rect 5236 8540 20188 8596
rect 20514 8540 20524 8596
rect 20580 8540 21420 8596
rect 21476 8540 23772 8596
rect 23828 8540 24668 8596
rect 24724 8540 24734 8596
rect 20132 8484 20188 8540
rect 4610 8428 4620 8484
rect 4676 8428 5292 8484
rect 5348 8428 5358 8484
rect 14802 8428 14812 8484
rect 14868 8428 16548 8484
rect 20132 8428 22876 8484
rect 22932 8428 22942 8484
rect 23202 8428 23212 8484
rect 23268 8428 23548 8484
rect 23604 8428 23614 8484
rect 31602 8428 31612 8484
rect 31668 8428 33740 8484
rect 33796 8428 33806 8484
rect 34066 8428 34076 8484
rect 34132 8428 41356 8484
rect 41412 8428 41422 8484
rect 45938 8428 45948 8484
rect 46004 8428 46396 8484
rect 46452 8428 46462 8484
rect 16492 8372 16548 8428
rect 33740 8372 33796 8428
rect 7074 8316 7084 8372
rect 7140 8316 8652 8372
rect 8708 8316 8718 8372
rect 11666 8316 11676 8372
rect 11732 8316 13132 8372
rect 13188 8316 13198 8372
rect 15026 8316 15036 8372
rect 15092 8316 15372 8372
rect 15428 8316 15438 8372
rect 16482 8316 16492 8372
rect 16548 8316 16558 8372
rect 16706 8316 16716 8372
rect 16772 8316 16940 8372
rect 16996 8316 17006 8372
rect 20178 8316 20188 8372
rect 20244 8316 25564 8372
rect 25620 8316 25630 8372
rect 28130 8316 28140 8372
rect 28196 8316 28700 8372
rect 28756 8316 30716 8372
rect 30772 8316 30782 8372
rect 33740 8316 35980 8372
rect 36036 8316 40908 8372
rect 40964 8316 40974 8372
rect 7746 8204 7756 8260
rect 7812 8204 8428 8260
rect 8484 8204 8494 8260
rect 12646 8204 12684 8260
rect 12740 8204 12750 8260
rect 16146 8204 16156 8260
rect 16212 8204 16828 8260
rect 16884 8204 16894 8260
rect 20626 8204 20636 8260
rect 20692 8204 21420 8260
rect 21476 8204 21486 8260
rect 23090 8204 23100 8260
rect 23156 8204 25228 8260
rect 25284 8204 25294 8260
rect 28354 8204 28364 8260
rect 28420 8204 28924 8260
rect 28980 8204 28990 8260
rect 35298 8204 35308 8260
rect 35364 8204 35868 8260
rect 35924 8204 37100 8260
rect 37156 8204 37166 8260
rect 6962 8092 6972 8148
rect 7028 8092 7924 8148
rect 9874 8092 9884 8148
rect 9940 8092 10668 8148
rect 10724 8092 10734 8148
rect 13010 8092 13020 8148
rect 13076 8092 16940 8148
rect 16996 8092 17006 8148
rect 17938 8092 17948 8148
rect 18004 8092 21308 8148
rect 21364 8092 21374 8148
rect 22194 8092 22204 8148
rect 22260 8092 22988 8148
rect 23044 8092 24892 8148
rect 24948 8092 26572 8148
rect 26628 8092 26638 8148
rect 33170 8092 33180 8148
rect 33236 8092 35084 8148
rect 35140 8092 36316 8148
rect 36372 8092 37772 8148
rect 37828 8092 37838 8148
rect 42130 8092 42140 8148
rect 42196 8092 48860 8148
rect 48916 8092 48926 8148
rect 7868 8036 7924 8092
rect 5282 7980 5292 8036
rect 5348 7980 7084 8036
rect 7140 7980 7150 8036
rect 7522 7980 7532 8036
rect 7588 7980 7598 8036
rect 7858 7980 7868 8036
rect 7924 7980 8988 8036
rect 9044 7980 9054 8036
rect 16482 7980 16492 8036
rect 16548 7980 19852 8036
rect 19908 7980 20244 8036
rect 20402 7980 20412 8036
rect 20468 7980 21644 8036
rect 21700 7980 25228 8036
rect 25284 7980 25294 8036
rect 25778 7980 25788 8036
rect 25844 7980 27580 8036
rect 27636 7980 27646 8036
rect 28466 7980 28476 8036
rect 28532 7980 29708 8036
rect 29764 7980 30268 8036
rect 30324 7980 30334 8036
rect 33282 7980 33292 8036
rect 33348 7980 33964 8036
rect 34020 7980 34030 8036
rect 34514 7980 34524 8036
rect 34580 7980 35980 8036
rect 36036 7980 36046 8036
rect 37874 7980 37884 8036
rect 37940 7980 39228 8036
rect 39284 7980 39294 8036
rect 42802 7980 42812 8036
rect 42868 7980 43372 8036
rect 43428 7980 43438 8036
rect 45714 7980 45724 8036
rect 45780 7980 46396 8036
rect 46452 7980 46462 8036
rect 7532 7924 7588 7980
rect 20188 7924 20244 7980
rect 7532 7868 8652 7924
rect 8708 7868 8718 7924
rect 13010 7868 13020 7924
rect 13076 7868 15596 7924
rect 15652 7868 15662 7924
rect 20188 7868 20972 7924
rect 21028 7868 21038 7924
rect 22754 7868 22764 7924
rect 22820 7868 24780 7924
rect 24836 7868 24846 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 12786 7756 12796 7812
rect 12852 7756 12862 7812
rect 22866 7756 22876 7812
rect 22932 7756 24332 7812
rect 24388 7756 25340 7812
rect 25396 7756 26124 7812
rect 26180 7756 26190 7812
rect 34738 7756 34748 7812
rect 34804 7756 40012 7812
rect 40068 7756 42588 7812
rect 42644 7756 42654 7812
rect 12796 7700 12852 7756
rect 9650 7644 9660 7700
rect 9716 7644 13020 7700
rect 13076 7644 13086 7700
rect 15092 7644 22204 7700
rect 22260 7644 22270 7700
rect 23090 7644 23100 7700
rect 23156 7644 23548 7700
rect 23604 7644 23614 7700
rect 31602 7644 31612 7700
rect 31668 7644 36204 7700
rect 36260 7644 36270 7700
rect 40114 7644 40124 7700
rect 40180 7644 41916 7700
rect 41972 7644 41982 7700
rect 45938 7644 45948 7700
rect 46004 7644 46620 7700
rect 46676 7644 49196 7700
rect 49252 7644 49262 7700
rect 15092 7588 15148 7644
rect 6066 7532 6076 7588
rect 6132 7532 12012 7588
rect 12068 7532 15148 7588
rect 21746 7532 21756 7588
rect 21812 7532 23324 7588
rect 23380 7532 23390 7588
rect 32722 7532 32732 7588
rect 32788 7532 33180 7588
rect 33236 7532 33246 7588
rect 33618 7532 33628 7588
rect 33684 7532 34188 7588
rect 34244 7532 34254 7588
rect 37874 7532 37884 7588
rect 37940 7532 45612 7588
rect 45668 7532 45678 7588
rect 46946 7532 46956 7588
rect 47012 7532 48412 7588
rect 48468 7532 48478 7588
rect 6514 7420 6524 7476
rect 6580 7420 8428 7476
rect 8484 7420 8988 7476
rect 9044 7420 14700 7476
rect 14756 7420 14766 7476
rect 19170 7420 19180 7476
rect 19236 7420 22652 7476
rect 22708 7420 22718 7476
rect 24546 7420 24556 7476
rect 24612 7420 26012 7476
rect 26068 7420 26078 7476
rect 27122 7420 27132 7476
rect 27188 7420 28476 7476
rect 28532 7420 29260 7476
rect 29316 7420 29326 7476
rect 29922 7420 29932 7476
rect 29988 7420 30604 7476
rect 30660 7420 31052 7476
rect 31108 7420 31118 7476
rect 31938 7420 31948 7476
rect 32004 7420 32956 7476
rect 33012 7420 33022 7476
rect 34850 7420 34860 7476
rect 34916 7420 37548 7476
rect 37604 7420 37772 7476
rect 37828 7420 37838 7476
rect 39778 7420 39788 7476
rect 39844 7420 41580 7476
rect 41636 7420 41646 7476
rect 47506 7420 47516 7476
rect 47572 7420 48972 7476
rect 49028 7420 49308 7476
rect 49364 7420 49374 7476
rect 12226 7308 12236 7364
rect 12292 7308 12684 7364
rect 12740 7308 13244 7364
rect 13300 7308 13692 7364
rect 13748 7308 13758 7364
rect 16818 7308 16828 7364
rect 16884 7308 17724 7364
rect 17780 7308 17790 7364
rect 24770 7308 24780 7364
rect 24836 7308 25676 7364
rect 25732 7308 26460 7364
rect 26516 7308 26526 7364
rect 31892 7308 38556 7364
rect 38612 7308 38622 7364
rect 39554 7308 39564 7364
rect 39620 7308 41132 7364
rect 41188 7308 41198 7364
rect 7746 7196 7756 7252
rect 7812 7196 8092 7252
rect 8148 7196 8158 7252
rect 12338 7196 12348 7252
rect 12404 7196 13916 7252
rect 13972 7196 13982 7252
rect 15474 7196 15484 7252
rect 15540 7196 30828 7252
rect 30884 7196 30894 7252
rect 12674 7084 12684 7140
rect 12740 7084 13020 7140
rect 13076 7084 13356 7140
rect 13412 7084 13422 7140
rect 14690 7084 14700 7140
rect 14756 7084 15596 7140
rect 15652 7084 15662 7140
rect 16258 7084 16268 7140
rect 16324 7084 17388 7140
rect 17444 7084 17454 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 6626 6972 6636 7028
rect 6692 6972 10892 7028
rect 10948 6972 10958 7028
rect 31892 6916 31948 7308
rect 34290 7196 34300 7252
rect 34356 7196 36876 7252
rect 36932 7196 36942 7252
rect 41234 7196 41244 7252
rect 41300 7196 43036 7252
rect 43092 7196 43102 7252
rect 45378 7196 45388 7252
rect 45444 7196 48748 7252
rect 48804 7196 48814 7252
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 6178 6860 6188 6916
rect 6244 6860 7084 6916
rect 7140 6860 7150 6916
rect 30818 6860 30828 6916
rect 30884 6860 31948 6916
rect 35074 6860 35084 6916
rect 35140 6860 35756 6916
rect 35812 6860 35822 6916
rect 36082 6860 36092 6916
rect 36148 6860 39788 6916
rect 39844 6860 39854 6916
rect 43026 6860 43036 6916
rect 43092 6860 43484 6916
rect 43540 6860 43550 6916
rect 5058 6748 5068 6804
rect 5124 6748 6636 6804
rect 6692 6748 8540 6804
rect 8596 6748 8606 6804
rect 10546 6748 10556 6804
rect 10612 6748 13580 6804
rect 13636 6748 13646 6804
rect 20626 6748 20636 6804
rect 20692 6748 21756 6804
rect 21812 6748 21822 6804
rect 30930 6748 30940 6804
rect 30996 6748 31836 6804
rect 31892 6748 33292 6804
rect 33348 6748 34580 6804
rect 36194 6748 36204 6804
rect 36260 6748 37548 6804
rect 37604 6748 37614 6804
rect 38210 6748 38220 6804
rect 38276 6748 38836 6804
rect 42466 6748 42476 6804
rect 42532 6748 47404 6804
rect 47460 6748 47470 6804
rect 34524 6692 34580 6748
rect 38780 6692 38836 6748
rect 6290 6636 6300 6692
rect 6356 6636 8764 6692
rect 8820 6636 8830 6692
rect 13122 6636 13132 6692
rect 13188 6636 13916 6692
rect 13972 6636 13982 6692
rect 14578 6636 14588 6692
rect 14644 6636 16828 6692
rect 16884 6636 16894 6692
rect 23426 6636 23436 6692
rect 23492 6636 24220 6692
rect 24276 6636 25452 6692
rect 25508 6636 25518 6692
rect 34514 6636 34524 6692
rect 34580 6636 34590 6692
rect 35634 6636 35644 6692
rect 35700 6636 36092 6692
rect 36148 6636 36988 6692
rect 37044 6636 37054 6692
rect 37436 6636 38668 6692
rect 38770 6636 38780 6692
rect 38836 6636 38846 6692
rect 39228 6636 44828 6692
rect 44884 6636 44894 6692
rect 46498 6636 46508 6692
rect 46564 6636 47292 6692
rect 47348 6636 47358 6692
rect 37436 6580 37492 6636
rect 8418 6524 8428 6580
rect 8484 6524 10108 6580
rect 10164 6524 10174 6580
rect 17826 6524 17836 6580
rect 17892 6524 18508 6580
rect 18564 6524 18574 6580
rect 20962 6524 20972 6580
rect 21028 6524 23660 6580
rect 23716 6524 23726 6580
rect 26898 6524 26908 6580
rect 26964 6524 28028 6580
rect 28084 6524 29036 6580
rect 29092 6524 30380 6580
rect 30436 6524 30446 6580
rect 35970 6524 35980 6580
rect 36036 6524 36428 6580
rect 36484 6524 37492 6580
rect 38612 6580 38668 6636
rect 39228 6580 39284 6636
rect 38612 6524 39284 6580
rect 39442 6524 39452 6580
rect 39508 6524 42140 6580
rect 42196 6524 43484 6580
rect 43540 6524 43550 6580
rect 45266 6524 45276 6580
rect 45332 6524 45612 6580
rect 45668 6524 46284 6580
rect 46340 6524 46350 6580
rect 28578 6412 28588 6468
rect 28644 6412 30492 6468
rect 30548 6412 30558 6468
rect 38322 6412 38332 6468
rect 38388 6412 42140 6468
rect 42196 6412 42206 6468
rect 42354 6412 42364 6468
rect 42420 6412 43036 6468
rect 43092 6412 43102 6468
rect 43250 6412 43260 6468
rect 43316 6412 45164 6468
rect 45220 6412 45230 6468
rect 45378 6412 45388 6468
rect 45444 6412 48972 6468
rect 49028 6412 49038 6468
rect 50200 6356 51000 6384
rect 17714 6300 17724 6356
rect 17780 6300 18508 6356
rect 18564 6300 18574 6356
rect 21970 6300 21980 6356
rect 22036 6300 47012 6356
rect 49186 6300 49196 6356
rect 49252 6300 51000 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 46956 6244 47012 6300
rect 50200 6272 51000 6300
rect 31378 6188 31388 6244
rect 31444 6188 36316 6244
rect 36372 6188 36382 6244
rect 36866 6188 36876 6244
rect 36932 6188 43820 6244
rect 43876 6188 43886 6244
rect 44818 6188 44828 6244
rect 44884 6188 45388 6244
rect 45444 6188 45454 6244
rect 46956 6188 47740 6244
rect 47796 6188 48972 6244
rect 49028 6188 49038 6244
rect 15586 6076 15596 6132
rect 15652 6076 17724 6132
rect 17780 6076 31948 6132
rect 32274 6076 32284 6132
rect 32340 6076 34300 6132
rect 34356 6076 34366 6132
rect 38098 6076 38108 6132
rect 38164 6076 38174 6132
rect 31892 6020 31948 6076
rect 38108 6020 38164 6076
rect 16146 5964 16156 6020
rect 16212 5964 18956 6020
rect 19012 5964 19404 6020
rect 19460 5964 20188 6020
rect 20244 5964 21420 6020
rect 21476 5964 21486 6020
rect 22978 5964 22988 6020
rect 23044 5964 24220 6020
rect 24276 5964 24286 6020
rect 31892 5964 38164 6020
rect 38612 5908 38668 6132
rect 38724 6076 38734 6132
rect 42130 6076 42140 6132
rect 42196 6076 44716 6132
rect 44772 6076 45724 6132
rect 45780 6076 49308 6132
rect 49364 6076 49374 6132
rect 39218 5964 39228 6020
rect 39284 5964 44044 6020
rect 44100 5964 44110 6020
rect 44258 5964 44268 6020
rect 44324 5964 45500 6020
rect 45556 5964 45566 6020
rect 46946 5964 46956 6020
rect 47012 5964 48188 6020
rect 48244 5964 48254 6020
rect 6076 5852 10444 5908
rect 10500 5852 10510 5908
rect 16930 5852 16940 5908
rect 16996 5852 18620 5908
rect 18676 5852 18686 5908
rect 20066 5852 20076 5908
rect 20132 5852 23436 5908
rect 23492 5852 23502 5908
rect 27794 5852 27804 5908
rect 27860 5852 31276 5908
rect 31332 5852 32508 5908
rect 32564 5852 32574 5908
rect 38322 5852 38332 5908
rect 38388 5852 38668 5908
rect 38966 5852 39004 5908
rect 39060 5852 39070 5908
rect 45154 5852 45164 5908
rect 45220 5852 46844 5908
rect 46900 5852 46910 5908
rect 6076 5796 6132 5852
rect 5170 5740 5180 5796
rect 5236 5740 6076 5796
rect 6132 5740 6142 5796
rect 8866 5740 8876 5796
rect 8932 5740 9996 5796
rect 10052 5740 10062 5796
rect 12114 5740 12124 5796
rect 12180 5740 13916 5796
rect 13972 5740 13982 5796
rect 17154 5740 17164 5796
rect 17220 5740 23548 5796
rect 23604 5740 23614 5796
rect 38770 5740 38780 5796
rect 38836 5740 40348 5796
rect 40404 5740 41020 5796
rect 41076 5740 41356 5796
rect 41412 5740 42924 5796
rect 42980 5740 42990 5796
rect 22418 5628 22428 5684
rect 22484 5628 23212 5684
rect 23268 5628 23278 5684
rect 26562 5628 26572 5684
rect 26628 5628 27020 5684
rect 27076 5628 27468 5684
rect 27524 5628 27534 5684
rect 32386 5628 32396 5684
rect 32452 5628 34076 5684
rect 34132 5628 34142 5684
rect 36418 5628 36428 5684
rect 36484 5628 39004 5684
rect 39060 5628 39070 5684
rect 45042 5628 45052 5684
rect 45108 5628 47628 5684
rect 47684 5628 47694 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 5170 5404 5180 5460
rect 5236 5404 21980 5460
rect 22036 5404 22046 5460
rect 4834 5292 4844 5348
rect 4900 5292 6524 5348
rect 6580 5292 36148 5348
rect 21522 5180 21532 5236
rect 21588 5180 22316 5236
rect 22372 5180 22382 5236
rect 23762 5180 23772 5236
rect 23828 5180 25228 5236
rect 25284 5180 25294 5236
rect 36092 5124 36148 5292
rect 43138 5180 43148 5236
rect 43204 5180 44044 5236
rect 44100 5180 44110 5236
rect 44370 5180 44380 5236
rect 44436 5180 46060 5236
rect 46116 5180 46126 5236
rect 8418 5068 8428 5124
rect 8484 5068 8988 5124
rect 9044 5068 9054 5124
rect 13346 5068 13356 5124
rect 13412 5068 13692 5124
rect 13748 5068 13758 5124
rect 18610 5068 18620 5124
rect 18676 5068 19740 5124
rect 19796 5068 22428 5124
rect 22484 5068 22494 5124
rect 26450 5068 26460 5124
rect 26516 5068 27580 5124
rect 27636 5068 27646 5124
rect 32946 5068 32956 5124
rect 33012 5068 34188 5124
rect 34244 5068 34254 5124
rect 34738 5068 34748 5124
rect 34804 5068 35420 5124
rect 35476 5068 35486 5124
rect 36092 5068 38220 5124
rect 38276 5068 38286 5124
rect 36092 5012 36148 5068
rect 5058 4956 5068 5012
rect 5124 4956 5516 5012
rect 5572 4956 8876 5012
rect 8932 4956 8942 5012
rect 10770 4956 10780 5012
rect 10836 4956 11788 5012
rect 11844 4956 11854 5012
rect 29586 4956 29596 5012
rect 29652 4956 30268 5012
rect 30324 4956 30334 5012
rect 31266 4956 31276 5012
rect 31332 4956 31612 5012
rect 31668 4956 31678 5012
rect 36082 4956 36092 5012
rect 36148 4956 36158 5012
rect 36316 4956 38668 5012
rect 41010 4956 41020 5012
rect 41076 4956 47516 5012
rect 47572 4956 47582 5012
rect 36316 4900 36372 4956
rect 6850 4844 6860 4900
rect 6916 4844 8540 4900
rect 8596 4844 9660 4900
rect 9716 4844 10444 4900
rect 10500 4844 10510 4900
rect 11218 4844 11228 4900
rect 11284 4844 15596 4900
rect 15652 4844 15662 4900
rect 26338 4844 26348 4900
rect 26404 4844 28140 4900
rect 28196 4844 28206 4900
rect 29698 4844 29708 4900
rect 29764 4844 30716 4900
rect 30772 4844 30782 4900
rect 32274 4844 32284 4900
rect 32340 4844 33852 4900
rect 33908 4844 36372 4900
rect 38612 4788 38668 4956
rect 38770 4844 38780 4900
rect 38836 4844 38874 4900
rect 39778 4844 39788 4900
rect 39844 4844 44156 4900
rect 44212 4844 44222 4900
rect 44930 4844 44940 4900
rect 44996 4844 45948 4900
rect 46004 4844 46014 4900
rect 29810 4732 29820 4788
rect 29876 4732 31276 4788
rect 31332 4732 31342 4788
rect 38612 4732 43260 4788
rect 43316 4732 43326 4788
rect 43474 4732 43484 4788
rect 43540 4732 43932 4788
rect 43988 4732 48748 4788
rect 48804 4732 48814 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 10882 4620 10892 4676
rect 10948 4620 15148 4676
rect 32386 4620 32396 4676
rect 32452 4620 33740 4676
rect 33796 4620 34412 4676
rect 34468 4620 35980 4676
rect 36036 4620 36046 4676
rect 38612 4620 49196 4676
rect 49252 4620 49262 4676
rect 15092 4564 15148 4620
rect 38612 4564 38668 4620
rect 11666 4508 11676 4564
rect 11732 4508 12684 4564
rect 12740 4508 12908 4564
rect 12964 4508 12974 4564
rect 15092 4508 38668 4564
rect 40562 4508 40572 4564
rect 40628 4508 44828 4564
rect 44884 4508 44894 4564
rect 11330 4396 11340 4452
rect 11396 4396 21868 4452
rect 21924 4396 21934 4452
rect 24658 4396 24668 4452
rect 24724 4396 25676 4452
rect 25732 4396 26684 4452
rect 26740 4396 26750 4452
rect 28018 4396 28028 4452
rect 28084 4396 31612 4452
rect 31668 4396 31678 4452
rect 32498 4396 32508 4452
rect 32564 4396 37884 4452
rect 37940 4396 37950 4452
rect 38098 4396 38108 4452
rect 38164 4396 44380 4452
rect 44436 4396 44446 4452
rect 16706 4284 16716 4340
rect 16772 4284 17500 4340
rect 17556 4284 17566 4340
rect 21186 4284 21196 4340
rect 21252 4284 23100 4340
rect 23156 4284 25452 4340
rect 25508 4284 25518 4340
rect 30258 4284 30268 4340
rect 30324 4284 31052 4340
rect 31108 4284 31118 4340
rect 33730 4284 33740 4340
rect 33796 4284 37212 4340
rect 37268 4284 37278 4340
rect 5842 4172 5852 4228
rect 5908 4172 8428 4228
rect 8484 4172 8494 4228
rect 23314 4172 23324 4228
rect 23380 4172 25340 4228
rect 25396 4172 25406 4228
rect 28242 4172 28252 4228
rect 28308 4172 31164 4228
rect 31220 4172 31230 4228
rect 46498 4172 46508 4228
rect 46564 4172 47740 4228
rect 47796 4172 47806 4228
rect 5058 4060 5068 4116
rect 5124 4060 8764 4116
rect 8820 4060 11900 4116
rect 11956 4060 12124 4116
rect 12180 4060 12190 4116
rect 12450 4060 12460 4116
rect 12516 4060 12526 4116
rect 17490 4060 17500 4116
rect 17556 4060 18508 4116
rect 18564 4060 18574 4116
rect 24546 4060 24556 4116
rect 24612 4060 26124 4116
rect 26180 4060 26190 4116
rect 36978 4060 36988 4116
rect 37044 4060 38556 4116
rect 38612 4060 38622 4116
rect 12460 4004 12516 4060
rect 9426 3948 9436 4004
rect 9492 3948 10220 4004
rect 10276 3948 12516 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 9090 3836 9100 3892
rect 9156 3836 9772 3892
rect 9828 3836 11676 3892
rect 11732 3836 11742 3892
rect 44482 3836 44492 3892
rect 44548 3836 48076 3892
rect 48132 3836 48142 3892
rect 8642 3724 8652 3780
rect 8708 3724 10780 3780
rect 10836 3724 10846 3780
rect 12002 3724 12012 3780
rect 12068 3724 13132 3780
rect 13188 3724 13198 3780
rect 35186 3724 35196 3780
rect 35252 3724 39340 3780
rect 39396 3724 39406 3780
rect 43250 3724 43260 3780
rect 43316 3724 47628 3780
rect 47684 3724 48636 3780
rect 48692 3724 48702 3780
rect 10780 3668 10836 3724
rect 10780 3612 13020 3668
rect 13076 3612 13086 3668
rect 30482 3612 30492 3668
rect 30548 3612 31612 3668
rect 31668 3612 31678 3668
rect 33394 3612 33404 3668
rect 33460 3612 40796 3668
rect 40852 3612 40862 3668
rect 42578 3612 42588 3668
rect 42644 3612 48748 3668
rect 48804 3612 48814 3668
rect 8754 3500 8764 3556
rect 8820 3500 13692 3556
rect 13748 3500 13758 3556
rect 16370 3500 16380 3556
rect 16436 3500 21756 3556
rect 21812 3500 21822 3556
rect 35074 3500 35084 3556
rect 35140 3500 39788 3556
rect 39844 3500 39854 3556
rect 44034 3500 44044 3556
rect 44100 3500 44828 3556
rect 44884 3500 44894 3556
rect 8194 3388 8204 3444
rect 8260 3388 11900 3444
rect 11956 3388 11966 3444
rect 29810 3388 29820 3444
rect 29876 3388 33068 3444
rect 33124 3388 33134 3444
rect 42998 3388 43036 3444
rect 43092 3388 43102 3444
rect 4722 3276 4732 3332
rect 4788 3276 5516 3332
rect 5572 3276 5582 3332
rect 7858 3276 7868 3332
rect 7924 3276 10108 3332
rect 10164 3276 10174 3332
rect 24434 3276 24444 3332
rect 24500 3276 28364 3332
rect 28420 3276 28430 3332
rect 31892 3276 32060 3332
rect 32116 3276 32126 3332
rect 42354 3276 42364 3332
rect 42420 3276 48076 3332
rect 48132 3276 48142 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 31892 2996 31948 3276
rect 37426 3164 37436 3220
rect 37492 3164 43932 3220
rect 43988 3164 43998 3220
rect 12226 2940 12236 2996
rect 12292 2940 31948 2996
rect 32162 2828 32172 2884
rect 32228 2828 45612 2884
rect 45668 2828 45678 2884
rect 6962 2716 6972 2772
rect 7028 2716 48972 2772
rect 49028 2716 49038 2772
rect 49186 2268 49196 2324
rect 49252 2268 49262 2324
rect 49196 2212 49252 2268
rect 49196 2156 50036 2212
rect 49980 2100 50036 2156
rect 50200 2100 51000 2128
rect 49980 2044 51000 2100
rect 50200 2016 51000 2044
<< via3 >>
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 32284 46956 32340 47012
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 45836 46172 45892 46228
rect 6076 45612 6132 45668
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 45836 44268 45892 44324
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 6076 43820 6132 43876
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 34972 42812 35028 42868
rect 18284 42476 18340 42532
rect 36428 42476 36484 42532
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 37660 42252 37716 42308
rect 48188 41804 48244 41860
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 17612 41132 17668 41188
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 40908 40236 40964 40292
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 30380 39452 30436 39508
rect 36428 39340 36484 39396
rect 17612 39228 17668 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 46284 39340 46340 39396
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 37660 38332 37716 38388
rect 18284 37996 18340 38052
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 34972 37548 35028 37604
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 40908 36540 40964 36596
rect 30380 36428 30436 36484
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 32284 35308 32340 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 40348 35196 40404 35252
rect 3388 34972 3444 35028
rect 3388 34636 3444 34692
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 30492 34300 30548 34356
rect 46508 34076 46564 34132
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 28588 33292 28644 33348
rect 31164 33068 31220 33124
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 48076 32844 48132 32900
rect 45500 32172 45556 32228
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 31164 32060 31220 32116
rect 40796 31500 40852 31556
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 29596 31276 29652 31332
rect 33852 31276 33908 31332
rect 31948 30828 32004 30884
rect 40460 30828 40516 30884
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 31164 30156 31220 30212
rect 31724 30156 31780 30212
rect 40236 30044 40292 30100
rect 48076 30156 48132 30212
rect 46284 30044 46340 30100
rect 45500 29820 45556 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 37996 29596 38052 29652
rect 40348 29596 40404 29652
rect 40236 29260 40292 29316
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 21196 28028 21252 28084
rect 46508 27580 46564 27636
rect 33852 27468 33908 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 37996 26908 38052 26964
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 30380 26572 30436 26628
rect 40796 26348 40852 26404
rect 30492 26124 30548 26180
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 37996 25676 38052 25732
rect 38892 25564 38948 25620
rect 38892 25340 38948 25396
rect 40796 25452 40852 25508
rect 31612 25228 31668 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 29596 25004 29652 25060
rect 21196 24780 21252 24836
rect 48076 24668 48132 24724
rect 28588 24444 28644 24500
rect 31612 24444 31668 24500
rect 31724 24332 31780 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 31948 23996 32004 24052
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 33628 23324 33684 23380
rect 35644 23100 35700 23156
rect 20972 22988 21028 23044
rect 33628 22764 33684 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 20188 22652 20244 22708
rect 20636 22652 20692 22708
rect 30940 22316 30996 22372
rect 40908 22204 40964 22260
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 33964 21868 34020 21924
rect 34188 21868 34244 21924
rect 37548 21756 37604 21812
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 33964 21084 34020 21140
rect 20636 20972 20692 21028
rect 33068 20860 33124 20916
rect 40460 20636 40516 20692
rect 37548 20524 37604 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 40908 20188 40964 20244
rect 42588 20076 42644 20132
rect 28476 19628 28532 19684
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 30604 19404 30660 19460
rect 20972 19292 21028 19348
rect 28252 19292 28308 19348
rect 30492 19292 30548 19348
rect 31276 19292 31332 19348
rect 21196 19180 21252 19236
rect 37436 19068 37492 19124
rect 20972 18956 21028 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 30604 18508 30660 18564
rect 36988 18284 37044 18340
rect 42588 18172 42644 18228
rect 30380 18060 30436 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 37660 18060 37716 18116
rect 39004 18060 39060 18116
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 38892 17948 38948 18004
rect 28364 17724 28420 17780
rect 30492 17724 30548 17780
rect 35644 17388 35700 17444
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 45836 17388 45892 17444
rect 45836 17052 45892 17108
rect 20188 16940 20244 16996
rect 28364 16940 28420 16996
rect 34188 16940 34244 16996
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 28476 16156 28532 16212
rect 28252 16044 28308 16100
rect 31276 16044 31332 16100
rect 38780 16044 38836 16100
rect 29932 15932 29988 15988
rect 30940 15932 30996 15988
rect 37436 15820 37492 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 19628 15596 19684 15652
rect 36988 15596 37044 15652
rect 38780 15372 38836 15428
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 39004 14812 39060 14868
rect 29932 14588 29988 14644
rect 37660 14476 37716 14532
rect 45836 14252 45892 14308
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 42364 13804 42420 13860
rect 33068 13692 33124 13748
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 42364 13020 42420 13076
rect 38668 12908 38724 12964
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19628 11228 19684 11284
rect 31836 11228 31892 11284
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 38668 11228 38724 11284
rect 43036 11228 43092 11284
rect 31836 10892 31892 10948
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 38780 9436 38836 9492
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 42588 8876 42644 8932
rect 23548 8652 23604 8708
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 23548 8428 23604 8484
rect 12684 8204 12740 8260
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 23548 7644 23604 7700
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 42140 6412 42196 6468
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 42140 6076 42196 6132
rect 39004 5852 39060 5908
rect 39004 5628 39060 5684
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 38780 4844 38836 4900
rect 43260 4732 43316 4788
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 12684 4508 12740 4564
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 43260 3724 43316 3780
rect 42588 3612 42644 3668
rect 43036 3388 43092 3444
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 47852 4768 47884
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 19808 47068 20128 47884
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 35168 47852 35488 47884
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 6076 45668 6132 45678
rect 6076 43876 6132 45612
rect 6076 43810 6132 43820
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 18284 42532 18340 42542
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 17612 41188 17668 41198
rect 17612 39284 17668 41132
rect 17612 39218 17668 39228
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 18284 38052 18340 42476
rect 18284 37986 18340 37996
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 32284 47012 32340 47022
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 3388 35028 3444 35038
rect 3388 34692 3444 34972
rect 3388 34626 3444 34636
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 30380 39508 30436 39518
rect 30380 36484 30436 39452
rect 30380 36418 30436 36428
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 32284 35364 32340 46956
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 45836 46228 45892 46238
rect 45836 44324 45892 46172
rect 45836 44258 45892 44268
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 34972 42868 35028 42878
rect 34972 37604 35028 42812
rect 34972 37538 35028 37548
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 36428 42532 36484 42542
rect 36428 39396 36484 42476
rect 36428 39330 36484 39340
rect 37660 42308 37716 42318
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 32284 35298 32340 35308
rect 35168 36876 35488 38388
rect 37660 38388 37716 42252
rect 48188 41860 48244 41870
rect 37660 38322 37716 38332
rect 40908 40292 40964 40302
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 40908 36596 40964 40236
rect 40908 36530 40964 36540
rect 46284 39396 46340 39406
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 30492 34356 30548 34366
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 28588 33348 28644 33358
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 21196 28084 21252 28094
rect 21196 24836 21252 28028
rect 20972 23044 21028 23054
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 20188 22708 20244 22718
rect 20188 16996 20244 22652
rect 20636 22708 20692 22718
rect 20636 21028 20692 22652
rect 20636 20962 20692 20972
rect 20972 19348 21028 22988
rect 20972 19012 21028 19292
rect 21196 19236 21252 24780
rect 28588 24500 28644 33292
rect 29596 31332 29652 31342
rect 29596 25060 29652 31276
rect 29596 24994 29652 25004
rect 30380 26628 30436 26638
rect 28588 24434 28644 24444
rect 28476 19684 28532 19694
rect 21196 19170 21252 19180
rect 28252 19348 28308 19358
rect 20972 18946 21028 18956
rect 20188 16930 20244 16940
rect 28252 16100 28308 19292
rect 28364 17780 28420 17790
rect 28364 16996 28420 17724
rect 28364 16930 28420 16940
rect 28476 16212 28532 19628
rect 30380 18116 30436 26572
rect 30492 26180 30548 34300
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 31164 33124 31220 33134
rect 31164 32116 31220 33068
rect 31164 30212 31220 32060
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 33852 31332 33908 31342
rect 31948 30884 32004 30894
rect 31164 30146 31220 30156
rect 31724 30212 31780 30222
rect 30492 26114 30548 26124
rect 31612 25284 31668 25294
rect 31612 24500 31668 25228
rect 31612 24434 31668 24444
rect 31724 24388 31780 30156
rect 31724 24322 31780 24332
rect 31948 24052 32004 30828
rect 33852 27524 33908 31276
rect 33852 27458 33908 27468
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 40348 35252 40404 35262
rect 40236 30100 40292 30110
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 31948 23986 32004 23996
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 37996 29652 38052 29662
rect 37996 26964 38052 29596
rect 40236 29316 40292 30044
rect 40348 29652 40404 35196
rect 45500 32228 45556 32238
rect 40796 31556 40852 31566
rect 40348 29586 40404 29596
rect 40460 30884 40516 30894
rect 40236 29250 40292 29260
rect 37996 25732 38052 26908
rect 37996 25666 38052 25676
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 33628 23380 33684 23390
rect 33628 22820 33684 23324
rect 33628 22754 33684 22764
rect 35168 22764 35488 24276
rect 38892 25620 38948 25630
rect 38892 25396 38948 25564
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 30940 22372 30996 22382
rect 30604 19460 30660 19470
rect 30380 18050 30436 18060
rect 30492 19348 30548 19358
rect 30492 17780 30548 19292
rect 30604 18564 30660 19404
rect 30604 18498 30660 18508
rect 30492 17714 30548 17724
rect 28476 16146 28532 16156
rect 28252 16034 28308 16044
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 19628 15652 19684 15662
rect 19628 11284 19684 15596
rect 19628 11218 19684 11228
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 29932 15988 29988 15998
rect 29932 14644 29988 15932
rect 30940 15988 30996 22316
rect 33964 21924 34020 21934
rect 33964 21140 34020 21868
rect 33964 21074 34020 21084
rect 34188 21924 34244 21934
rect 33068 20916 33124 20926
rect 31276 19348 31332 19358
rect 31276 16100 31332 19292
rect 31276 16034 31332 16044
rect 30940 15922 30996 15932
rect 29932 14578 29988 14588
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 33068 13748 33124 20860
rect 34188 16996 34244 21868
rect 34188 16930 34244 16940
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 33068 13682 33124 13692
rect 35168 16492 35488 18004
rect 35644 23156 35700 23166
rect 35644 17444 35700 23100
rect 37548 21812 37604 21822
rect 37548 20580 37604 21756
rect 37548 20514 37604 20524
rect 37436 19124 37492 19134
rect 35644 17378 35700 17388
rect 36988 18340 37044 18350
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 36988 15652 37044 18284
rect 37436 15876 37492 19068
rect 37436 15810 37492 15820
rect 37660 18116 37716 18126
rect 36988 15586 37044 15596
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 19808 11004 20128 12516
rect 35168 13356 35488 14868
rect 37660 14532 37716 18060
rect 38892 18004 38948 25340
rect 40460 20692 40516 30828
rect 40796 26404 40852 31500
rect 45500 29876 45556 32172
rect 46284 30100 46340 39340
rect 46284 30034 46340 30044
rect 46508 34132 46564 34142
rect 45500 29810 45556 29820
rect 46508 27636 46564 34076
rect 48076 32900 48132 32910
rect 48076 30212 48132 32844
rect 48076 30146 48132 30156
rect 46508 27570 46564 27580
rect 48188 26908 48244 41804
rect 40796 25508 40852 26348
rect 40796 25442 40852 25452
rect 48076 26852 48244 26908
rect 48076 24724 48132 26852
rect 48076 24658 48132 24668
rect 40460 20626 40516 20636
rect 40908 22260 40964 22270
rect 40908 20244 40964 22204
rect 40908 20178 40964 20188
rect 42588 20132 42644 20142
rect 42588 18228 42644 20076
rect 42588 18162 42644 18172
rect 38892 17938 38948 17948
rect 39004 18116 39060 18126
rect 38780 16100 38836 16110
rect 38780 15428 38836 16044
rect 38780 15362 38836 15372
rect 39004 14868 39060 18060
rect 39004 14802 39060 14812
rect 45836 17444 45892 17454
rect 45836 17108 45892 17388
rect 37660 14466 37716 14476
rect 45836 14308 45892 17052
rect 45836 14242 45892 14252
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 42364 13860 42420 13870
rect 42364 13076 42420 13804
rect 42364 13010 42420 13020
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 31836 11284 31892 11294
rect 31836 10948 31892 11228
rect 31836 10882 31892 10892
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 12684 8260 12740 8270
rect 12684 4564 12740 8204
rect 12684 4498 12740 4508
rect 19808 7868 20128 9380
rect 35168 10220 35488 11732
rect 38668 12964 38724 12974
rect 38668 11284 38724 12908
rect 38668 11218 38724 11228
rect 43036 11284 43092 11294
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 23548 8708 23604 8718
rect 23548 8484 23604 8652
rect 23548 7700 23604 8428
rect 23548 7634 23604 7644
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 38780 9492 38836 9502
rect 38780 4900 38836 9436
rect 42588 8932 42644 8942
rect 42140 6468 42196 6478
rect 42140 6132 42196 6412
rect 42140 6066 42196 6076
rect 39004 5908 39060 5918
rect 39004 5684 39060 5852
rect 39004 5618 39060 5628
rect 38780 4834 38836 4844
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 42588 3668 42644 8876
rect 42588 3602 42644 3612
rect 43036 3444 43092 11228
rect 43260 4788 43316 4798
rect 43260 3780 43316 4732
rect 43260 3714 43316 3724
rect 43036 3378 43092 3388
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1190_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1191_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20160 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1192_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24080 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1193_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22848 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1194_
timestamp 1698431365
transform -1 0 17696 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1195_
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1196_
timestamp 1698431365
transform 1 0 18816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1197_
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1198_
timestamp 1698431365
transform -1 0 20720 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1199_
timestamp 1698431365
transform 1 0 19264 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1200_
timestamp 1698431365
transform -1 0 32704 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1201_
timestamp 1698431365
transform 1 0 30016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1202_
timestamp 1698431365
transform -1 0 35280 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1203_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32256 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1204_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46704 0 1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1205_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31024 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1206_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1207_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1208_
timestamp 1698431365
transform -1 0 33376 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1209_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1210_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1211_
timestamp 1698431365
transform -1 0 19152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1212_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1213_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26656 0 1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1214_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27216 0 -1 15680
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1215_
timestamp 1698431365
transform -1 0 29904 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1216_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28336 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1217_
timestamp 1698431365
transform 1 0 30912 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1218_
timestamp 1698431365
transform -1 0 28560 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1219_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1220_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1221_
timestamp 1698431365
transform -1 0 30352 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1222_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30576 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1223_
timestamp 1698431365
transform 1 0 5600 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1224_
timestamp 1698431365
transform -1 0 7504 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1225_
timestamp 1698431365
transform -1 0 10080 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1226_
timestamp 1698431365
transform 1 0 5600 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1227_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7840 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1228_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1229_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8064 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1230_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7952 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1231_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4928 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1232_
timestamp 1698431365
transform 1 0 5712 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1233_
timestamp 1698431365
transform -1 0 6832 0 -1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1234_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1235_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5936 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1236_
timestamp 1698431365
transform -1 0 7952 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1237_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6160 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1238_
timestamp 1698431365
transform 1 0 7168 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1239_
timestamp 1698431365
transform -1 0 8848 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1240_
timestamp 1698431365
transform -1 0 8624 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1241_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7952 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1242_
timestamp 1698431365
transform -1 0 7056 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1243_
timestamp 1698431365
transform -1 0 6160 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1244_
timestamp 1698431365
transform -1 0 5152 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1245_
timestamp 1698431365
transform -1 0 6608 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1246_
timestamp 1698431365
transform -1 0 7504 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1247_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5152 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1248_
timestamp 1698431365
transform 1 0 7280 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1249_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1250_
timestamp 1698431365
transform 1 0 6608 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1251_
timestamp 1698431365
transform -1 0 3696 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1252_
timestamp 1698431365
transform -1 0 10864 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1253_
timestamp 1698431365
transform -1 0 10080 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1254_
timestamp 1698431365
transform 1 0 8624 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1255_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11424 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1256_
timestamp 1698431365
transform -1 0 8400 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1257_
timestamp 1698431365
transform -1 0 13104 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1258_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10864 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1259_
timestamp 1698431365
transform -1 0 12544 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1260_
timestamp 1698431365
transform -1 0 6832 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1261_
timestamp 1698431365
transform -1 0 6160 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1262_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11088 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1263_
timestamp 1698431365
transform -1 0 8624 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1264_
timestamp 1698431365
transform -1 0 5488 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1265_
timestamp 1698431365
transform -1 0 4592 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1266_
timestamp 1698431365
transform -1 0 5040 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1267_
timestamp 1698431365
transform -1 0 3136 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1268_
timestamp 1698431365
transform 1 0 5936 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1269_
timestamp 1698431365
transform 1 0 5936 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1270_
timestamp 1698431365
transform 1 0 6272 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1271_
timestamp 1698431365
transform 1 0 7504 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1272_
timestamp 1698431365
transform 1 0 5040 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1273_
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1274_
timestamp 1698431365
transform -1 0 6496 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1275_
timestamp 1698431365
transform -1 0 3136 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1276_
timestamp 1698431365
transform -1 0 8288 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1277_
timestamp 1698431365
transform 1 0 8064 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1278_
timestamp 1698431365
transform 1 0 8176 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1279_
timestamp 1698431365
transform 1 0 8400 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1280_
timestamp 1698431365
transform -1 0 8064 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1281_
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1282_
timestamp 1698431365
transform -1 0 7056 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1283_
timestamp 1698431365
transform 1 0 7056 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1284_
timestamp 1698431365
transform 1 0 7952 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1285_
timestamp 1698431365
transform 1 0 9744 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1286_
timestamp 1698431365
transform -1 0 11088 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1287_
timestamp 1698431365
transform 1 0 7840 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1288_
timestamp 1698431365
transform 1 0 11200 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1289_
timestamp 1698431365
transform -1 0 9184 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1290_
timestamp 1698431365
transform -1 0 9632 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1291_
timestamp 1698431365
transform -1 0 11312 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1292_
timestamp 1698431365
transform -1 0 12320 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1293_
timestamp 1698431365
transform 1 0 8736 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1294_
timestamp 1698431365
transform 1 0 7280 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1295_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6832 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1296_
timestamp 1698431365
transform -1 0 7168 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1297_
timestamp 1698431365
transform -1 0 11200 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1298_
timestamp 1698431365
transform -1 0 10640 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1299_
timestamp 1698431365
transform 1 0 9408 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1300_
timestamp 1698431365
transform -1 0 6832 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1301_
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1302_
timestamp 1698431365
transform -1 0 8960 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1303_
timestamp 1698431365
transform -1 0 8176 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1304_
timestamp 1698431365
transform -1 0 4368 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1305_
timestamp 1698431365
transform -1 0 5264 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1306_
timestamp 1698431365
transform -1 0 5040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1307_
timestamp 1698431365
transform 1 0 5040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1308_
timestamp 1698431365
transform 1 0 3248 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1309_
timestamp 1698431365
transform -1 0 3024 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1310_
timestamp 1698431365
transform -1 0 6384 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1311_
timestamp 1698431365
transform 1 0 5712 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1312_
timestamp 1698431365
transform -1 0 6944 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1313_
timestamp 1698431365
transform 1 0 8176 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1314_
timestamp 1698431365
transform -1 0 8064 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1315_
timestamp 1698431365
transform -1 0 7504 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1316_
timestamp 1698431365
transform -1 0 5488 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1317_
timestamp 1698431365
transform -1 0 5264 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1318_
timestamp 1698431365
transform -1 0 3472 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1319_
timestamp 1698431365
transform -1 0 4368 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1320_
timestamp 1698431365
transform -1 0 5824 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1321_
timestamp 1698431365
transform 1 0 4032 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1322_
timestamp 1698431365
transform 1 0 3136 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1323_
timestamp 1698431365
transform -1 0 2800 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1324_
timestamp 1698431365
transform -1 0 8400 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1325_
timestamp 1698431365
transform 1 0 3024 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1326_
timestamp 1698431365
transform -1 0 5040 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1327_
timestamp 1698431365
transform -1 0 3696 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1328_
timestamp 1698431365
transform -1 0 2800 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1329_
timestamp 1698431365
transform -1 0 5152 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1330_
timestamp 1698431365
transform -1 0 2464 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1331_
timestamp 1698431365
transform 1 0 1680 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1332_
timestamp 1698431365
transform -1 0 2464 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1333_
timestamp 1698431365
transform 1 0 3360 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1334_
timestamp 1698431365
transform -1 0 3360 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1335_
timestamp 1698431365
transform -1 0 2912 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1336_
timestamp 1698431365
transform -1 0 6160 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1337_
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1338_
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1339_
timestamp 1698431365
transform -1 0 3472 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1340_
timestamp 1698431365
transform -1 0 5264 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1341_
timestamp 1698431365
transform 1 0 2912 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1342_
timestamp 1698431365
transform -1 0 5264 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1343_
timestamp 1698431365
transform 1 0 3920 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1344_
timestamp 1698431365
transform 1 0 6160 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1345_
timestamp 1698431365
transform -1 0 40544 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1346_
timestamp 1698431365
transform -1 0 39760 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1347_
timestamp 1698431365
transform -1 0 35728 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1348_
timestamp 1698431365
transform -1 0 35616 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1349_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41216 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1350_
timestamp 1698431365
transform -1 0 42336 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1351_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1352_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35728 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1353_
timestamp 1698431365
transform 1 0 35840 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1354_
timestamp 1698431365
transform 1 0 34272 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1355_
timestamp 1698431365
transform 1 0 34272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1356_
timestamp 1698431365
transform 1 0 35056 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1357_
timestamp 1698431365
transform 1 0 37520 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1358_
timestamp 1698431365
transform -1 0 36848 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1359_
timestamp 1698431365
transform 1 0 33600 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1360_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35392 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1361_
timestamp 1698431365
transform -1 0 33936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1362_
timestamp 1698431365
transform 1 0 26656 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1363_
timestamp 1698431365
transform -1 0 35504 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1364_
timestamp 1698431365
transform 1 0 33152 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1365_
timestamp 1698431365
transform -1 0 32704 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1366_
timestamp 1698431365
transform -1 0 34944 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1367_
timestamp 1698431365
transform 1 0 33040 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1368_
timestamp 1698431365
transform -1 0 39648 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1369_
timestamp 1698431365
transform -1 0 38976 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1370_
timestamp 1698431365
transform -1 0 41216 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1371_
timestamp 1698431365
transform -1 0 40096 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1372_
timestamp 1698431365
transform -1 0 37968 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1373_
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1374_
timestamp 1698431365
transform -1 0 36624 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1375_
timestamp 1698431365
transform -1 0 27664 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1376_
timestamp 1698431365
transform 1 0 36288 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1377_
timestamp 1698431365
transform 1 0 36848 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1378_
timestamp 1698431365
transform -1 0 34384 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1379_
timestamp 1698431365
transform -1 0 20944 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1380_
timestamp 1698431365
transform 1 0 20272 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1381_
timestamp 1698431365
transform 1 0 23520 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1382_
timestamp 1698431365
transform -1 0 21392 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1383_
timestamp 1698431365
transform -1 0 23520 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1384_
timestamp 1698431365
transform -1 0 21952 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1385_
timestamp 1698431365
transform 1 0 19824 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1386_
timestamp 1698431365
transform 1 0 26320 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1387_
timestamp 1698431365
transform -1 0 19824 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1388_
timestamp 1698431365
transform -1 0 21504 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1389_
timestamp 1698431365
transform -1 0 30912 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1390_
timestamp 1698431365
transform 1 0 26768 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1391_
timestamp 1698431365
transform 1 0 27776 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1392_
timestamp 1698431365
transform 1 0 27104 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1393_
timestamp 1698431365
transform 1 0 22512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1394_
timestamp 1698431365
transform -1 0 38528 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1395_
timestamp 1698431365
transform 1 0 23408 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1396_
timestamp 1698431365
transform 1 0 22512 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1397_
timestamp 1698431365
transform -1 0 21952 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1398_
timestamp 1698431365
transform 1 0 22176 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1399_
timestamp 1698431365
transform -1 0 30016 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1400_
timestamp 1698431365
transform -1 0 31472 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1401_
timestamp 1698431365
transform 1 0 34944 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1402_
timestamp 1698431365
transform 1 0 35616 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1403_
timestamp 1698431365
transform -1 0 39088 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1404_
timestamp 1698431365
transform -1 0 30688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1405_
timestamp 1698431365
transform -1 0 28784 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1406_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28560 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1407_
timestamp 1698431365
transform 1 0 29904 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1408_
timestamp 1698431365
transform -1 0 30240 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1409_
timestamp 1698431365
transform 1 0 30240 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1410_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1411_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27328 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1412_
timestamp 1698431365
transform 1 0 27328 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1413_
timestamp 1698431365
transform -1 0 27104 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1414_
timestamp 1698431365
transform -1 0 27216 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1415_
timestamp 1698431365
transform -1 0 24864 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1416_
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1417_
timestamp 1698431365
transform -1 0 27888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1418_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29904 0 -1 7840
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1419_
timestamp 1698431365
transform 1 0 25648 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1420_
timestamp 1698431365
transform 1 0 25312 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1421_
timestamp 1698431365
transform -1 0 26656 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1422_
timestamp 1698431365
transform -1 0 24752 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1423_
timestamp 1698431365
transform 1 0 22624 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1424_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1425_
timestamp 1698431365
transform -1 0 24640 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1426_
timestamp 1698431365
transform 1 0 19936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1427_
timestamp 1698431365
transform -1 0 25984 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1428_
timestamp 1698431365
transform -1 0 21952 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1429_
timestamp 1698431365
transform 1 0 24192 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1430_
timestamp 1698431365
transform -1 0 23968 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1431_
timestamp 1698431365
transform -1 0 20944 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1432_
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1433_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1434_
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1435_
timestamp 1698431365
transform 1 0 20384 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1436_
timestamp 1698431365
transform -1 0 22512 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1437_
timestamp 1698431365
transform -1 0 18144 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1438_
timestamp 1698431365
transform 1 0 22848 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1439_
timestamp 1698431365
transform -1 0 24752 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1440_
timestamp 1698431365
transform 1 0 34384 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1441_
timestamp 1698431365
transform -1 0 35616 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1442_
timestamp 1698431365
transform -1 0 37296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1443_
timestamp 1698431365
transform 1 0 35504 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1444_
timestamp 1698431365
transform 1 0 35616 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1445_
timestamp 1698431365
transform 1 0 44016 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1446_
timestamp 1698431365
transform -1 0 41888 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1447_
timestamp 1698431365
transform 1 0 34272 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1448_
timestamp 1698431365
transform -1 0 34272 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1449_
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1450_
timestamp 1698431365
transform 1 0 33488 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1451_
timestamp 1698431365
transform 1 0 26992 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1452_
timestamp 1698431365
transform 1 0 37632 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1453_
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1454_
timestamp 1698431365
transform -1 0 40208 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1455_
timestamp 1698431365
transform -1 0 31808 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1456_
timestamp 1698431365
transform 1 0 22400 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1457_
timestamp 1698431365
transform -1 0 49280 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1458_
timestamp 1698431365
transform 1 0 37408 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1459_
timestamp 1698431365
transform -1 0 49280 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1460_
timestamp 1698431365
transform 1 0 41776 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1461_
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1462_
timestamp 1698431365
transform -1 0 44352 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1463_
timestamp 1698431365
transform -1 0 34496 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1464_
timestamp 1698431365
transform -1 0 43904 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1465_
timestamp 1698431365
transform -1 0 43232 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1466_
timestamp 1698431365
transform -1 0 49280 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1467_
timestamp 1698431365
transform 1 0 44800 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1468_
timestamp 1698431365
transform 1 0 45136 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1469_
timestamp 1698431365
transform -1 0 32704 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1470_
timestamp 1698431365
transform -1 0 48048 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1471_
timestamp 1698431365
transform 1 0 46368 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1472_
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1473_
timestamp 1698431365
transform 1 0 47264 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1474_
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1475_
timestamp 1698431365
transform -1 0 47264 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1476_
timestamp 1698431365
transform -1 0 46256 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1477_
timestamp 1698431365
transform -1 0 46144 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1478_
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1479_
timestamp 1698431365
transform -1 0 26880 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1480_
timestamp 1698431365
transform -1 0 27664 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1481_
timestamp 1698431365
transform -1 0 25984 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1482_
timestamp 1698431365
transform -1 0 26208 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1483_
timestamp 1698431365
transform 1 0 25312 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1484_
timestamp 1698431365
transform -1 0 24864 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1485_
timestamp 1698431365
transform -1 0 23520 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1486_
timestamp 1698431365
transform 1 0 22624 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1487_
timestamp 1698431365
transform -1 0 22176 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1488_
timestamp 1698431365
transform -1 0 20272 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1489_
timestamp 1698431365
transform 1 0 18032 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1490_
timestamp 1698431365
transform -1 0 22624 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1491_
timestamp 1698431365
transform 1 0 19376 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1492_
timestamp 1698431365
transform -1 0 19040 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1493_
timestamp 1698431365
transform 1 0 13440 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1494_
timestamp 1698431365
transform -1 0 16128 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1495_
timestamp 1698431365
transform -1 0 16128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1496_
timestamp 1698431365
transform 1 0 38528 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1497_
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1498_
timestamp 1698431365
transform -1 0 18368 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1499_
timestamp 1698431365
transform -1 0 17024 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1500_
timestamp 1698431365
transform -1 0 17024 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1501_
timestamp 1698431365
transform 1 0 14336 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1502_
timestamp 1698431365
transform -1 0 33824 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1503_
timestamp 1698431365
transform 1 0 15344 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1504_
timestamp 1698431365
transform 1 0 16240 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1505_
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1506_
timestamp 1698431365
transform -1 0 34944 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1507_
timestamp 1698431365
transform -1 0 27888 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1508_
timestamp 1698431365
transform -1 0 24192 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1509_
timestamp 1698431365
transform 1 0 24192 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1510_
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1511_
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1512_
timestamp 1698431365
transform 1 0 26096 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1513_
timestamp 1698431365
transform 1 0 26432 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1514_
timestamp 1698431365
transform 1 0 26208 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1515_
timestamp 1698431365
transform 1 0 26544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1516_
timestamp 1698431365
transform 1 0 25312 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1517_
timestamp 1698431365
transform 1 0 24304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1518_
timestamp 1698431365
transform -1 0 24192 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1519_
timestamp 1698431365
transform -1 0 23520 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1520_
timestamp 1698431365
transform 1 0 22512 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1521_
timestamp 1698431365
transform 1 0 22400 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1522_
timestamp 1698431365
transform 1 0 35616 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1523_
timestamp 1698431365
transform 1 0 22736 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1524_
timestamp 1698431365
transform 1 0 22848 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1525_
timestamp 1698431365
transform -1 0 39088 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1526_
timestamp 1698431365
transform 1 0 21840 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1527_
timestamp 1698431365
transform 1 0 20160 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1528_
timestamp 1698431365
transform -1 0 39872 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1529_
timestamp 1698431365
transform 1 0 21728 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1530_
timestamp 1698431365
transform -1 0 20272 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1531_
timestamp 1698431365
transform 1 0 35952 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1532_
timestamp 1698431365
transform -1 0 36400 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1533_
timestamp 1698431365
transform -1 0 38416 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1534_
timestamp 1698431365
transform -1 0 34048 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1535_
timestamp 1698431365
transform -1 0 31696 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1536_
timestamp 1698431365
transform -1 0 30128 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1537_
timestamp 1698431365
transform -1 0 28448 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1538_
timestamp 1698431365
transform 1 0 26768 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1539_
timestamp 1698431365
transform -1 0 29568 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1540_
timestamp 1698431365
transform 1 0 26208 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1541_
timestamp 1698431365
transform 1 0 30128 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1542_
timestamp 1698431365
transform -1 0 31472 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1543_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1544_
timestamp 1698431365
transform -1 0 32256 0 -1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1545_
timestamp 1698431365
transform 1 0 30128 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1546_
timestamp 1698431365
transform -1 0 34384 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1547_
timestamp 1698431365
transform -1 0 41216 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1548_
timestamp 1698431365
transform 1 0 30128 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1549_
timestamp 1698431365
transform 1 0 31584 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1550_
timestamp 1698431365
transform 1 0 35056 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1551_
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1552_
timestamp 1698431365
transform -1 0 36400 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1553_
timestamp 1698431365
transform -1 0 32704 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1554_
timestamp 1698431365
transform 1 0 34944 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1555_
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1556_
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1557_
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1558_
timestamp 1698431365
transform -1 0 29008 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1559_
timestamp 1698431365
transform -1 0 31584 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1560_
timestamp 1698431365
transform -1 0 30800 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1561_
timestamp 1698431365
transform -1 0 30352 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1562_
timestamp 1698431365
transform -1 0 30240 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1563_
timestamp 1698431365
transform 1 0 28336 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1564_
timestamp 1698431365
transform 1 0 27104 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1565_
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1566_
timestamp 1698431365
transform 1 0 27104 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1567_
timestamp 1698431365
transform -1 0 26544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1568_
timestamp 1698431365
transform 1 0 34496 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1569_
timestamp 1698431365
transform -1 0 31808 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1570_
timestamp 1698431365
transform 1 0 32144 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1571_
timestamp 1698431365
transform 1 0 34608 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1572_
timestamp 1698431365
transform -1 0 36624 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1573_
timestamp 1698431365
transform 1 0 34832 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1574_
timestamp 1698431365
transform -1 0 36848 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1575_
timestamp 1698431365
transform 1 0 33936 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1576_
timestamp 1698431365
transform -1 0 34384 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1577_
timestamp 1698431365
transform 1 0 31808 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1578_
timestamp 1698431365
transform 1 0 31248 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1579_
timestamp 1698431365
transform 1 0 33936 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1580_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1581_
timestamp 1698431365
transform -1 0 32704 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1582_
timestamp 1698431365
transform -1 0 23968 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1583_
timestamp 1698431365
transform -1 0 23072 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1584_
timestamp 1698431365
transform -1 0 22176 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1585_
timestamp 1698431365
transform -1 0 20496 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1586_
timestamp 1698431365
transform 1 0 19600 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1587_
timestamp 1698431365
transform -1 0 19600 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1588_
timestamp 1698431365
transform 1 0 19936 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1589_
timestamp 1698431365
transform 1 0 18704 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1590_
timestamp 1698431365
transform -1 0 18704 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1591_
timestamp 1698431365
transform -1 0 12656 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1592_
timestamp 1698431365
transform -1 0 11424 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1593_
timestamp 1698431365
transform -1 0 11872 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1594_
timestamp 1698431365
transform 1 0 11424 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1595_
timestamp 1698431365
transform 1 0 10976 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1596_
timestamp 1698431365
transform -1 0 13440 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1597_
timestamp 1698431365
transform -1 0 10976 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1598_
timestamp 1698431365
transform -1 0 10080 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1599_
timestamp 1698431365
transform 1 0 12880 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1600_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1601_
timestamp 1698431365
transform 1 0 13440 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1602_
timestamp 1698431365
transform 1 0 13664 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1603_
timestamp 1698431365
transform 1 0 15008 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1604_
timestamp 1698431365
transform 1 0 11872 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1605_
timestamp 1698431365
transform -1 0 15792 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1606_
timestamp 1698431365
transform 1 0 7840 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1607_
timestamp 1698431365
transform 1 0 7504 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1608_
timestamp 1698431365
transform -1 0 7504 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1609_
timestamp 1698431365
transform 1 0 8288 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1610_
timestamp 1698431365
transform 1 0 7392 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1611_
timestamp 1698431365
transform -1 0 7392 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1612_
timestamp 1698431365
transform -1 0 8512 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1613_
timestamp 1698431365
transform -1 0 10752 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1614_
timestamp 1698431365
transform 1 0 7616 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1615_
timestamp 1698431365
transform -1 0 7616 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1616_
timestamp 1698431365
transform -1 0 7616 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1617_
timestamp 1698431365
transform 1 0 7616 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1618_
timestamp 1698431365
transform 1 0 8176 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1619_
timestamp 1698431365
transform 1 0 10080 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1620_
timestamp 1698431365
transform 1 0 8512 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1621_
timestamp 1698431365
transform -1 0 9856 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1622_
timestamp 1698431365
transform 1 0 9408 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1623_
timestamp 1698431365
transform 1 0 12768 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1624_
timestamp 1698431365
transform 1 0 11536 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1625_
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1626_
timestamp 1698431365
transform 1 0 13440 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1627_
timestamp 1698431365
transform 1 0 14784 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1628_
timestamp 1698431365
transform 1 0 11872 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1629_
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1630_
timestamp 1698431365
transform -1 0 40208 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1631_
timestamp 1698431365
transform -1 0 39200 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1632_
timestamp 1698431365
transform -1 0 33712 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1633_
timestamp 1698431365
transform 1 0 27104 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1634_
timestamp 1698431365
transform 1 0 26320 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1635_
timestamp 1698431365
transform 1 0 43568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1636_
timestamp 1698431365
transform -1 0 30464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1637_
timestamp 1698431365
transform 1 0 27888 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1638_
timestamp 1698431365
transform 1 0 27664 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1639_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1640_
timestamp 1698431365
transform 1 0 38528 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1641_
timestamp 1698431365
transform -1 0 40544 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1642_
timestamp 1698431365
transform 1 0 37856 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1643_
timestamp 1698431365
transform -1 0 40432 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1644_
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1645_
timestamp 1698431365
transform 1 0 38080 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1646_
timestamp 1698431365
transform -1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1647_
timestamp 1698431365
transform -1 0 39648 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1648_
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1649_
timestamp 1698431365
transform -1 0 41776 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1650_
timestamp 1698431365
transform 1 0 39648 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1651_
timestamp 1698431365
transform -1 0 39088 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1652_
timestamp 1698431365
transform -1 0 38192 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1653_
timestamp 1698431365
transform -1 0 37296 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1654_
timestamp 1698431365
transform 1 0 36960 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1655_
timestamp 1698431365
transform -1 0 40096 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1656_
timestamp 1698431365
transform 1 0 37744 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1657_
timestamp 1698431365
transform -1 0 41664 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1658_
timestamp 1698431365
transform 1 0 38192 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1659_
timestamp 1698431365
transform -1 0 39088 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1660_
timestamp 1698431365
transform -1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1661_
timestamp 1698431365
transform 1 0 41888 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1662_
timestamp 1698431365
transform -1 0 34048 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1663_
timestamp 1698431365
transform -1 0 29680 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1664_
timestamp 1698431365
transform -1 0 33264 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1665_
timestamp 1698431365
transform -1 0 29008 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1666_
timestamp 1698431365
transform 1 0 26208 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1667_
timestamp 1698431365
transform 1 0 26656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1668_
timestamp 1698431365
transform 1 0 42000 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1669_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1670_
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1671_
timestamp 1698431365
transform 1 0 41104 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1672_
timestamp 1698431365
transform 1 0 27216 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1673_
timestamp 1698431365
transform -1 0 25536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1674_
timestamp 1698431365
transform 1 0 41216 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1675_
timestamp 1698431365
transform 1 0 27216 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1676_
timestamp 1698431365
transform 1 0 26544 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1677_
timestamp 1698431365
transform -1 0 25648 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1678_
timestamp 1698431365
transform -1 0 24976 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1679_
timestamp 1698431365
transform 1 0 22288 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1680_
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1681_
timestamp 1698431365
transform 1 0 23296 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1682_
timestamp 1698431365
transform 1 0 22848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1683_
timestamp 1698431365
transform 1 0 19936 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1684_
timestamp 1698431365
transform 1 0 19488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1685_
timestamp 1698431365
transform -1 0 22848 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1686_
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1687_
timestamp 1698431365
transform -1 0 37744 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1688_
timestamp 1698431365
transform -1 0 33376 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1689_
timestamp 1698431365
transform -1 0 44352 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1690_
timestamp 1698431365
transform 1 0 35952 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1691_
timestamp 1698431365
transform -1 0 39648 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1692_
timestamp 1698431365
transform 1 0 35280 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1693_
timestamp 1698431365
transform -1 0 14224 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1694_
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1695_
timestamp 1698431365
transform -1 0 34608 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1696_
timestamp 1698431365
transform -1 0 32368 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1697_
timestamp 1698431365
transform 1 0 33040 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1698_
timestamp 1698431365
transform -1 0 32592 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1699_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1700_
timestamp 1698431365
transform -1 0 25984 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1701_
timestamp 1698431365
transform -1 0 31920 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1702_
timestamp 1698431365
transform -1 0 31360 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1703_
timestamp 1698431365
transform -1 0 31024 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1704_
timestamp 1698431365
transform -1 0 28672 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1705_
timestamp 1698431365
transform 1 0 27216 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1706_
timestamp 1698431365
transform -1 0 25536 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1707_
timestamp 1698431365
transform -1 0 32256 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1708_
timestamp 1698431365
transform -1 0 31136 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1709_
timestamp 1698431365
transform -1 0 34720 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1710_
timestamp 1698431365
transform 1 0 32928 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1711_
timestamp 1698431365
transform 1 0 36960 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1712_
timestamp 1698431365
transform 1 0 40432 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1713_
timestamp 1698431365
transform 1 0 44800 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1714_
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1715_
timestamp 1698431365
transform 1 0 46480 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1716_
timestamp 1698431365
transform -1 0 49056 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1717_
timestamp 1698431365
transform -1 0 49280 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1718_
timestamp 1698431365
transform 1 0 44800 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1719_
timestamp 1698431365
transform 1 0 45360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1720_
timestamp 1698431365
transform 1 0 43904 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1721_
timestamp 1698431365
transform -1 0 48048 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1722_
timestamp 1698431365
transform -1 0 45584 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1723_
timestamp 1698431365
transform 1 0 45584 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1724_
timestamp 1698431365
transform 1 0 44800 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1725_
timestamp 1698431365
transform 1 0 47936 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1726_
timestamp 1698431365
transform 1 0 47824 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1727_
timestamp 1698431365
transform -1 0 46480 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1728_
timestamp 1698431365
transform 1 0 46928 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1729_
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1730_
timestamp 1698431365
transform 1 0 48832 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1731_
timestamp 1698431365
transform -1 0 47824 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1732_
timestamp 1698431365
transform -1 0 46928 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1733_
timestamp 1698431365
transform 1 0 47152 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1734_
timestamp 1698431365
transform 1 0 48048 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1735_
timestamp 1698431365
transform -1 0 48384 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1736_
timestamp 1698431365
transform -1 0 49280 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1737_
timestamp 1698431365
transform -1 0 49056 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1738_
timestamp 1698431365
transform -1 0 49056 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1739_
timestamp 1698431365
transform 1 0 47376 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1740_
timestamp 1698431365
transform -1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1741_
timestamp 1698431365
transform -1 0 47936 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1742_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1743_
timestamp 1698431365
transform -1 0 47152 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1744_
timestamp 1698431365
transform -1 0 45696 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1745_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1746_
timestamp 1698431365
transform 1 0 40768 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1747_
timestamp 1698431365
transform -1 0 43120 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1748_
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1749_
timestamp 1698431365
transform 1 0 45360 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1750_
timestamp 1698431365
transform -1 0 41888 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1751_
timestamp 1698431365
transform 1 0 42224 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1752_
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1753_
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1754_
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1755_
timestamp 1698431365
transform 1 0 46256 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1756_
timestamp 1698431365
transform 1 0 46816 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1757_
timestamp 1698431365
transform -1 0 49280 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1758_
timestamp 1698431365
transform -1 0 48384 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1759_
timestamp 1698431365
transform -1 0 49056 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1760_
timestamp 1698431365
transform 1 0 46928 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1761_
timestamp 1698431365
transform 1 0 42672 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1762_
timestamp 1698431365
transform -1 0 45808 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1763_
timestamp 1698431365
transform -1 0 44464 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1764_
timestamp 1698431365
transform -1 0 48384 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1765_
timestamp 1698431365
transform -1 0 45248 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1766_
timestamp 1698431365
transform -1 0 44800 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1767_
timestamp 1698431365
transform -1 0 49280 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1768_
timestamp 1698431365
transform 1 0 41664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1769_
timestamp 1698431365
transform 1 0 43344 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1770_
timestamp 1698431365
transform -1 0 49280 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1771_
timestamp 1698431365
transform -1 0 43904 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1772_
timestamp 1698431365
transform 1 0 43456 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1773_
timestamp 1698431365
transform 1 0 41104 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1774_
timestamp 1698431365
transform -1 0 45136 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1775_
timestamp 1698431365
transform -1 0 43792 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1776_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45696 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1777_
timestamp 1698431365
transform -1 0 44352 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1778_
timestamp 1698431365
transform 1 0 43232 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1779_
timestamp 1698431365
transform 1 0 42000 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1780_
timestamp 1698431365
transform -1 0 43456 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1781_
timestamp 1698431365
transform -1 0 48048 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1782_
timestamp 1698431365
transform 1 0 41552 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1783_
timestamp 1698431365
transform 1 0 44688 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1784_
timestamp 1698431365
transform 1 0 43792 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1785_
timestamp 1698431365
transform 1 0 44016 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1786_
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1787_
timestamp 1698431365
transform 1 0 44800 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1788_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45136 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1789_
timestamp 1698431365
transform -1 0 45136 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1790_
timestamp 1698431365
transform -1 0 42784 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1791_
timestamp 1698431365
transform 1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1792_
timestamp 1698431365
transform -1 0 48384 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1793_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45920 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1794_
timestamp 1698431365
transform 1 0 42000 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1795_
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1796_
timestamp 1698431365
transform -1 0 43792 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1797_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46704 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1798_
timestamp 1698431365
transform -1 0 48496 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1799_
timestamp 1698431365
transform -1 0 44464 0 1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1800_
timestamp 1698431365
transform 1 0 46032 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1801_
timestamp 1698431365
transform -1 0 46256 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1802_
timestamp 1698431365
transform 1 0 43120 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1803_
timestamp 1698431365
transform -1 0 49392 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1804_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41776 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1805_
timestamp 1698431365
transform 1 0 41104 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1806_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42560 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1807_
timestamp 1698431365
transform 1 0 42896 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1808_
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1809_
timestamp 1698431365
transform -1 0 47152 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1810_
timestamp 1698431365
transform 1 0 47152 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1811_
timestamp 1698431365
transform -1 0 47264 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1812_
timestamp 1698431365
transform -1 0 43344 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1813_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42896 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1814_
timestamp 1698431365
transform -1 0 42336 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1815_
timestamp 1698431365
transform 1 0 30688 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1816_
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1817_
timestamp 1698431365
transform -1 0 32256 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1818_
timestamp 1698431365
transform -1 0 39872 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1819_
timestamp 1698431365
transform 1 0 37184 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1820_
timestamp 1698431365
transform -1 0 41888 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1821_
timestamp 1698431365
transform -1 0 44912 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1822_
timestamp 1698431365
transform -1 0 40768 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1823_
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1824_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32480 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1825_
timestamp 1698431365
transform -1 0 40544 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1826_
timestamp 1698431365
transform 1 0 40208 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1827_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1828_
timestamp 1698431365
transform 1 0 39200 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1829_
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1830_
timestamp 1698431365
transform -1 0 49280 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1831_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45360 0 -1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1832_
timestamp 1698431365
transform 1 0 41776 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1833_
timestamp 1698431365
transform 1 0 43568 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1834_
timestamp 1698431365
transform 1 0 47488 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1835_
timestamp 1698431365
transform 1 0 47824 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1836_
timestamp 1698431365
transform 1 0 43904 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1837_
timestamp 1698431365
transform 1 0 44576 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1838_
timestamp 1698431365
transform 1 0 46928 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1839_
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1840_
timestamp 1698431365
transform -1 0 49280 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1841_
timestamp 1698431365
transform -1 0 46928 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1842_
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1843_
timestamp 1698431365
transform -1 0 49280 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1844_
timestamp 1698431365
transform 1 0 45136 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1845_
timestamp 1698431365
transform -1 0 49280 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1846_
timestamp 1698431365
transform 1 0 45808 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1847_
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1848_
timestamp 1698431365
transform 1 0 43344 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1849_
timestamp 1698431365
transform 1 0 47936 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1850_
timestamp 1698431365
transform -1 0 49280 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1851_
timestamp 1698431365
transform 1 0 45024 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1852_
timestamp 1698431365
transform 1 0 45248 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1853_
timestamp 1698431365
transform 1 0 44912 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1854_
timestamp 1698431365
transform -1 0 46480 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1855_
timestamp 1698431365
transform 1 0 46480 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1856_
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1857_
timestamp 1698431365
transform 1 0 47488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1858_
timestamp 1698431365
transform -1 0 47488 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1859_
timestamp 1698431365
transform 1 0 46928 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1860_
timestamp 1698431365
transform -1 0 42784 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1861_
timestamp 1698431365
transform -1 0 46928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1862_
timestamp 1698431365
transform 1 0 46928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1863_
timestamp 1698431365
transform -1 0 46704 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1864_
timestamp 1698431365
transform -1 0 41776 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1865_
timestamp 1698431365
transform 1 0 47040 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1866_
timestamp 1698431365
transform -1 0 48832 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1867_
timestamp 1698431365
transform 1 0 45248 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1868_
timestamp 1698431365
transform -1 0 47040 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1869_
timestamp 1698431365
transform -1 0 46032 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1870_
timestamp 1698431365
transform -1 0 44464 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1871_
timestamp 1698431365
transform -1 0 42000 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1872_
timestamp 1698431365
transform 1 0 41776 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1873_
timestamp 1698431365
transform 1 0 41552 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1874_
timestamp 1698431365
transform 1 0 42336 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1875_
timestamp 1698431365
transform 1 0 44800 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1876_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46480 0 -1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1877_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46368 0 -1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1878_
timestamp 1698431365
transform -1 0 46144 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1879_
timestamp 1698431365
transform 1 0 45248 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1880_
timestamp 1698431365
transform 1 0 45136 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1881_
timestamp 1698431365
transform -1 0 13104 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1882_
timestamp 1698431365
transform -1 0 12096 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1883_
timestamp 1698431365
transform 1 0 11424 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1884_
timestamp 1698431365
transform 1 0 12544 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1885_
timestamp 1698431365
transform -1 0 12656 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1886_
timestamp 1698431365
transform -1 0 7840 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1887_
timestamp 1698431365
transform 1 0 7616 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1888_
timestamp 1698431365
transform 1 0 12320 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1889_
timestamp 1698431365
transform -1 0 15680 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1890_
timestamp 1698431365
transform 1 0 14336 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1891_
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1892_
timestamp 1698431365
transform 1 0 10976 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1893_
timestamp 1698431365
transform -1 0 12096 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1894_
timestamp 1698431365
transform 1 0 11424 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1895_
timestamp 1698431365
transform -1 0 8512 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1896_
timestamp 1698431365
transform 1 0 9296 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1897_
timestamp 1698431365
transform 1 0 10528 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1898_
timestamp 1698431365
transform -1 0 10528 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1899_
timestamp 1698431365
transform 1 0 7280 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1900_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1901_
timestamp 1698431365
transform -1 0 7056 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1902_
timestamp 1698431365
transform 1 0 7056 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1903_
timestamp 1698431365
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1904_
timestamp 1698431365
transform -1 0 9632 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1905_
timestamp 1698431365
transform -1 0 7168 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1906_
timestamp 1698431365
transform -1 0 9968 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1907_
timestamp 1698431365
transform -1 0 9072 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1908_
timestamp 1698431365
transform -1 0 9072 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1909_
timestamp 1698431365
transform -1 0 9968 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1910_
timestamp 1698431365
transform -1 0 9072 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1911_
timestamp 1698431365
transform -1 0 7952 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1912_
timestamp 1698431365
transform -1 0 9968 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1913_
timestamp 1698431365
transform -1 0 6608 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1914_
timestamp 1698431365
transform -1 0 6160 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1915_
timestamp 1698431365
transform 1 0 4816 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1916_
timestamp 1698431365
transform -1 0 6944 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1917_
timestamp 1698431365
transform -1 0 6048 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1918_
timestamp 1698431365
transform -1 0 6384 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1919_
timestamp 1698431365
transform -1 0 4816 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1920_
timestamp 1698431365
transform -1 0 6496 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1921_
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1922_
timestamp 1698431365
transform 1 0 2800 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1923_
timestamp 1698431365
transform -1 0 2800 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1924_
timestamp 1698431365
transform 1 0 2800 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1925_
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1926_
timestamp 1698431365
transform -1 0 3136 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1927_
timestamp 1698431365
transform -1 0 2576 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1928_
timestamp 1698431365
transform -1 0 2464 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1929_
timestamp 1698431365
transform -1 0 6832 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1930_
timestamp 1698431365
transform -1 0 7392 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1931_
timestamp 1698431365
transform -1 0 7280 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1932_
timestamp 1698431365
transform -1 0 6720 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1933_
timestamp 1698431365
transform 1 0 3136 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1934_
timestamp 1698431365
transform 1 0 3024 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1935_
timestamp 1698431365
transform -1 0 7168 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1936_
timestamp 1698431365
transform 1 0 3584 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1937_
timestamp 1698431365
transform 1 0 4144 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1939_
timestamp 1698431365
transform -1 0 6944 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1940_
timestamp 1698431365
transform -1 0 6384 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1941_
timestamp 1698431365
transform -1 0 6048 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1942_
timestamp 1698431365
transform 1 0 3248 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1943_
timestamp 1698431365
transform 1 0 3808 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1944_
timestamp 1698431365
transform 1 0 6944 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1945_
timestamp 1698431365
transform 1 0 6384 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1946_
timestamp 1698431365
transform 1 0 6944 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1947_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1948_
timestamp 1698431365
transform 1 0 4032 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1949_
timestamp 1698431365
transform 1 0 4704 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1950_
timestamp 1698431365
transform 1 0 5936 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1951_
timestamp 1698431365
transform 1 0 9184 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1952_
timestamp 1698431365
transform 1 0 10304 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1953_
timestamp 1698431365
transform 1 0 8288 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1954_
timestamp 1698431365
transform -1 0 8848 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1955_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1956_
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1957_
timestamp 1698431365
transform -1 0 36624 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1958_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1959_
timestamp 1698431365
transform 1 0 33600 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1960_
timestamp 1698431365
transform 1 0 35616 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1961_
timestamp 1698431365
transform 1 0 33376 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1962_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1963_
timestamp 1698431365
transform 1 0 35504 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1964_
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1965_
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1966_
timestamp 1698431365
transform 1 0 37072 0 -1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1967_
timestamp 1698431365
transform -1 0 38752 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1968_
timestamp 1698431365
transform -1 0 40544 0 -1 28224
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1969_
timestamp 1698431365
transform 1 0 33824 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1970_
timestamp 1698431365
transform 1 0 35168 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1971_
timestamp 1698431365
transform -1 0 35616 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1972_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1973_
timestamp 1698431365
transform -1 0 37856 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1974_
timestamp 1698431365
transform 1 0 34160 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1975_
timestamp 1698431365
transform 1 0 25984 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1976_
timestamp 1698431365
transform 1 0 33264 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1977_
timestamp 1698431365
transform 1 0 35280 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1978_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1979_
timestamp 1698431365
transform -1 0 36848 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1980_
timestamp 1698431365
transform -1 0 35616 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1981_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1982_
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1983_
timestamp 1698431365
transform 1 0 36736 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1984_
timestamp 1698431365
transform 1 0 37744 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1985_
timestamp 1698431365
transform -1 0 49280 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1986_
timestamp 1698431365
transform -1 0 24640 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1987_
timestamp 1698431365
transform -1 0 31808 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1988_
timestamp 1698431365
transform -1 0 24192 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1989_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1990_
timestamp 1698431365
transform 1 0 20496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1991_
timestamp 1698431365
transform -1 0 20944 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1992_
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1993_
timestamp 1698431365
transform 1 0 19040 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1994_
timestamp 1698431365
transform 1 0 18928 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1995_
timestamp 1698431365
transform 1 0 15456 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1996_
timestamp 1698431365
transform 1 0 17920 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1997_
timestamp 1698431365
transform -1 0 19040 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1998_
timestamp 1698431365
transform -1 0 19488 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1999_
timestamp 1698431365
transform 1 0 14896 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2000_
timestamp 1698431365
transform 1 0 17920 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2001_
timestamp 1698431365
transform -1 0 20608 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2002_
timestamp 1698431365
transform 1 0 19152 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2003_
timestamp 1698431365
transform -1 0 18928 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2004_
timestamp 1698431365
transform -1 0 20832 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2005_
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2006_
timestamp 1698431365
transform -1 0 21840 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2007_
timestamp 1698431365
transform -1 0 24304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2008_
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2009_
timestamp 1698431365
transform -1 0 20832 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2010_
timestamp 1698431365
transform -1 0 19488 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2011_
timestamp 1698431365
transform 1 0 18368 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2012_
timestamp 1698431365
transform 1 0 19376 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2013_
timestamp 1698431365
transform -1 0 22288 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2014_
timestamp 1698431365
transform -1 0 20272 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2015_
timestamp 1698431365
transform 1 0 19488 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2016_
timestamp 1698431365
transform 1 0 20384 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2017_
timestamp 1698431365
transform -1 0 21392 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2018_
timestamp 1698431365
transform -1 0 19376 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2019_
timestamp 1698431365
transform -1 0 18592 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2020_
timestamp 1698431365
transform -1 0 16128 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2021_
timestamp 1698431365
transform 1 0 16800 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2022_
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2023_
timestamp 1698431365
transform 1 0 17696 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2024_
timestamp 1698431365
transform 1 0 17808 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2025_
timestamp 1698431365
transform -1 0 22848 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2026_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 1 36064
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2027_
timestamp 1698431365
transform -1 0 20944 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2028_
timestamp 1698431365
transform 1 0 18928 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2029_
timestamp 1698431365
transform -1 0 22064 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2030_
timestamp 1698431365
transform 1 0 21392 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2031_
timestamp 1698431365
transform -1 0 21392 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2032_
timestamp 1698431365
transform -1 0 20384 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2033_
timestamp 1698431365
transform 1 0 18592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2034_
timestamp 1698431365
transform -1 0 19376 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2035_
timestamp 1698431365
transform -1 0 20384 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2036_
timestamp 1698431365
transform 1 0 18704 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2037_
timestamp 1698431365
transform 1 0 19152 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2038_
timestamp 1698431365
transform 1 0 20048 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2039_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24192 0 -1 37632
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2040_
timestamp 1698431365
transform 1 0 31136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2041_
timestamp 1698431365
transform 1 0 21616 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2042_
timestamp 1698431365
transform 1 0 22288 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2043_
timestamp 1698431365
transform -1 0 21392 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2044_
timestamp 1698431365
transform -1 0 26656 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2045_
timestamp 1698431365
transform 1 0 22288 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2046_
timestamp 1698431365
transform 1 0 21168 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2047_
timestamp 1698431365
transform -1 0 23856 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2048_
timestamp 1698431365
transform 1 0 17136 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2049_
timestamp 1698431365
transform 1 0 17472 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2050_
timestamp 1698431365
transform -1 0 19152 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2051_
timestamp 1698431365
transform -1 0 17920 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2052_
timestamp 1698431365
transform 1 0 15680 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2053_
timestamp 1698431365
transform -1 0 17248 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2054_
timestamp 1698431365
transform -1 0 15344 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2055_
timestamp 1698431365
transform 1 0 17696 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2056_
timestamp 1698431365
transform 1 0 16576 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2057_
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2058_
timestamp 1698431365
transform -1 0 17920 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2059_
timestamp 1698431365
transform -1 0 14784 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2060_
timestamp 1698431365
transform -1 0 17024 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2061_
timestamp 1698431365
transform -1 0 19152 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2062_
timestamp 1698431365
transform 1 0 14784 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2063_
timestamp 1698431365
transform -1 0 14448 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2064_
timestamp 1698431365
transform 1 0 13328 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2065_
timestamp 1698431365
transform -1 0 16912 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2066_
timestamp 1698431365
transform -1 0 14336 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2067_
timestamp 1698431365
transform 1 0 12432 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2068_
timestamp 1698431365
transform 1 0 15568 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2069_
timestamp 1698431365
transform 1 0 14672 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2070_
timestamp 1698431365
transform 1 0 16016 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2071_
timestamp 1698431365
transform 1 0 14560 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2072_
timestamp 1698431365
transform -1 0 16128 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2073_
timestamp 1698431365
transform -1 0 16464 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2074_
timestamp 1698431365
transform -1 0 14560 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2075_
timestamp 1698431365
transform 1 0 12432 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2076_
timestamp 1698431365
transform 1 0 15792 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2077_
timestamp 1698431365
transform -1 0 17584 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2078_
timestamp 1698431365
transform -1 0 18592 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2079_
timestamp 1698431365
transform -1 0 16688 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2080_
timestamp 1698431365
transform -1 0 14000 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2081_
timestamp 1698431365
transform -1 0 17808 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2082_
timestamp 1698431365
transform -1 0 18032 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2083_
timestamp 1698431365
transform -1 0 17024 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2084_
timestamp 1698431365
transform 1 0 13664 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2085_
timestamp 1698431365
transform 1 0 24864 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2086_
timestamp 1698431365
transform -1 0 19040 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2087_
timestamp 1698431365
transform 1 0 28112 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2088_
timestamp 1698431365
transform -1 0 30128 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2089_
timestamp 1698431365
transform 1 0 29344 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _2090_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34944 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2091_
timestamp 1698431365
transform -1 0 32704 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2092_
timestamp 1698431365
transform -1 0 30464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2093_
timestamp 1698431365
transform -1 0 30240 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2094_
timestamp 1698431365
transform -1 0 31136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2095_
timestamp 1698431365
transform -1 0 28224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2096_
timestamp 1698431365
transform 1 0 29232 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2097_
timestamp 1698431365
transform 1 0 29120 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2098_
timestamp 1698431365
transform 1 0 29120 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2099_
timestamp 1698431365
transform -1 0 30016 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2100_
timestamp 1698431365
transform -1 0 30016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2101_
timestamp 1698431365
transform -1 0 29568 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2102_
timestamp 1698431365
transform -1 0 28560 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2103_
timestamp 1698431365
transform 1 0 28112 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2104_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2105_
timestamp 1698431365
transform 1 0 29680 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2106_
timestamp 1698431365
transform -1 0 36288 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2107_
timestamp 1698431365
transform -1 0 34944 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2108_
timestamp 1698431365
transform -1 0 36064 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2109_
timestamp 1698431365
transform -1 0 34048 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2110_
timestamp 1698431365
transform -1 0 36288 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2111_
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2112_
timestamp 1698431365
transform 1 0 30912 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2113_
timestamp 1698431365
transform -1 0 34496 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2114_
timestamp 1698431365
transform -1 0 32704 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2115_
timestamp 1698431365
transform -1 0 32368 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2116_
timestamp 1698431365
transform 1 0 33376 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2117_
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2118_
timestamp 1698431365
transform -1 0 34160 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2119_
timestamp 1698431365
transform -1 0 32704 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2120_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2121_
timestamp 1698431365
transform 1 0 27104 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2122_
timestamp 1698431365
transform -1 0 29456 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2123_
timestamp 1698431365
transform 1 0 27776 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2124_
timestamp 1698431365
transform 1 0 27552 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2125_
timestamp 1698431365
transform 1 0 28112 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2126_
timestamp 1698431365
transform 1 0 29008 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2127_
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2128_
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _2129_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39648 0 -1 39200
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2130_
timestamp 1698431365
transform -1 0 32480 0 -1 40768
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2131_
timestamp 1698431365
transform 1 0 32032 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2132_
timestamp 1698431365
transform -1 0 36512 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2133_
timestamp 1698431365
transform 1 0 34048 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2134_
timestamp 1698431365
transform -1 0 33824 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2135_
timestamp 1698431365
transform -1 0 33376 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2136_
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2137_
timestamp 1698431365
transform -1 0 32032 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2138_
timestamp 1698431365
transform 1 0 30688 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2139_
timestamp 1698431365
transform 1 0 29568 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2140_
timestamp 1698431365
transform 1 0 30240 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2141_
timestamp 1698431365
transform 1 0 30016 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2142_
timestamp 1698431365
transform -1 0 34944 0 1 40768
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2143_
timestamp 1698431365
transform -1 0 32144 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2144_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2145_
timestamp 1698431365
transform 1 0 31472 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2146_
timestamp 1698431365
transform 1 0 31584 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2147_
timestamp 1698431365
transform -1 0 38192 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2148_
timestamp 1698431365
transform 1 0 32480 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2149_
timestamp 1698431365
transform -1 0 35392 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2150_
timestamp 1698431365
transform 1 0 32032 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2151_
timestamp 1698431365
transform 1 0 34496 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2152_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2153_
timestamp 1698431365
transform 1 0 35728 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2154_
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2155_
timestamp 1698431365
transform 1 0 34384 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2156_
timestamp 1698431365
transform 1 0 35728 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2157_
timestamp 1698431365
transform -1 0 36512 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2158_
timestamp 1698431365
transform 1 0 34160 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2159_
timestamp 1698431365
transform -1 0 32704 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2160_
timestamp 1698431365
transform -1 0 31024 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2161_
timestamp 1698431365
transform 1 0 31920 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2162_
timestamp 1698431365
transform 1 0 27328 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2163_
timestamp 1698431365
transform 1 0 30464 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2164_
timestamp 1698431365
transform -1 0 34160 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2165_
timestamp 1698431365
transform 1 0 29792 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2166_
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2167_
timestamp 1698431365
transform -1 0 29904 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2168_
timestamp 1698431365
transform 1 0 26656 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2169_
timestamp 1698431365
transform -1 0 27776 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2170_
timestamp 1698431365
transform -1 0 25760 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2171_
timestamp 1698431365
transform -1 0 29120 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2172_
timestamp 1698431365
transform 1 0 27776 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2173_
timestamp 1698431365
transform -1 0 26880 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2174_
timestamp 1698431365
transform -1 0 27776 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2175_
timestamp 1698431365
transform -1 0 26768 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2176_
timestamp 1698431365
transform -1 0 29120 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2177_
timestamp 1698431365
transform 1 0 27888 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2178_
timestamp 1698431365
transform 1 0 29008 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2179_
timestamp 1698431365
transform -1 0 27776 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2180_
timestamp 1698431365
transform -1 0 27888 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2181_
timestamp 1698431365
transform -1 0 28896 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2182_
timestamp 1698431365
transform -1 0 27776 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2183_
timestamp 1698431365
transform 1 0 25312 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2184_
timestamp 1698431365
transform -1 0 28000 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2185_
timestamp 1698431365
transform -1 0 28560 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2186_
timestamp 1698431365
transform -1 0 27440 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2187_
timestamp 1698431365
transform -1 0 26096 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2188_
timestamp 1698431365
transform -1 0 28784 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2189_
timestamp 1698431365
transform -1 0 32368 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2190_
timestamp 1698431365
transform 1 0 31024 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2191_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2192_
timestamp 1698431365
transform -1 0 23184 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2193_
timestamp 1698431365
transform -1 0 24528 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2194_
timestamp 1698431365
transform 1 0 13328 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2195_
timestamp 1698431365
transform -1 0 19936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2196_
timestamp 1698431365
transform -1 0 19824 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2197_
timestamp 1698431365
transform -1 0 17024 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2198_
timestamp 1698431365
transform 1 0 16016 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2199_
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2200_
timestamp 1698431365
transform 1 0 16464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2201_
timestamp 1698431365
transform -1 0 17696 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2202_
timestamp 1698431365
transform -1 0 20384 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2203_
timestamp 1698431365
transform -1 0 17024 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2204_
timestamp 1698431365
transform -1 0 16352 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2205_
timestamp 1698431365
transform 1 0 15008 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2206_
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2207_
timestamp 1698431365
transform -1 0 18256 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2208_
timestamp 1698431365
transform 1 0 15680 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2209_
timestamp 1698431365
transform -1 0 16912 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2210_
timestamp 1698431365
transform -1 0 16800 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2211_
timestamp 1698431365
transform 1 0 16912 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2212_
timestamp 1698431365
transform -1 0 24192 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2213_
timestamp 1698431365
transform 1 0 19040 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2214_
timestamp 1698431365
transform 1 0 15568 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2215_
timestamp 1698431365
transform -1 0 15456 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2216_
timestamp 1698431365
transform 1 0 14224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2217_
timestamp 1698431365
transform 1 0 16016 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2218_
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2219_
timestamp 1698431365
transform 1 0 14672 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2220_
timestamp 1698431365
transform 1 0 14672 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2221_
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2222_
timestamp 1698431365
transform 1 0 17024 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2223_
timestamp 1698431365
transform -1 0 16240 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2224_
timestamp 1698431365
transform 1 0 14448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2225_
timestamp 1698431365
transform -1 0 16352 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2226_
timestamp 1698431365
transform 1 0 14896 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2227_
timestamp 1698431365
transform 1 0 14448 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2228_
timestamp 1698431365
transform 1 0 15344 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2229_
timestamp 1698431365
transform 1 0 15904 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2230_
timestamp 1698431365
transform -1 0 19600 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2231_
timestamp 1698431365
transform 1 0 18144 0 1 28224
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2232_
timestamp 1698431365
transform 1 0 17136 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2233_
timestamp 1698431365
transform -1 0 18704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2234_
timestamp 1698431365
transform 1 0 17584 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2235_
timestamp 1698431365
transform 1 0 18144 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2236_
timestamp 1698431365
transform -1 0 17024 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2237_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2238_
timestamp 1698431365
transform -1 0 16800 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2239_
timestamp 1698431365
transform -1 0 17136 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2240_
timestamp 1698431365
transform -1 0 17696 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2241_
timestamp 1698431365
transform 1 0 17584 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2242_
timestamp 1698431365
transform 1 0 19040 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2243_
timestamp 1698431365
transform 1 0 18592 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _2244_
timestamp 1698431365
transform 1 0 17472 0 -1 25088
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2245_
timestamp 1698431365
transform 1 0 30016 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2246_
timestamp 1698431365
transform -1 0 21616 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2247_
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2248_
timestamp 1698431365
transform -1 0 20944 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _2249_
timestamp 1698431365
transform -1 0 26656 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2250_
timestamp 1698431365
transform -1 0 22064 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2251_
timestamp 1698431365
transform -1 0 22288 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2252_
timestamp 1698431365
transform 1 0 19824 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2253_
timestamp 1698431365
transform 1 0 14000 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2254_
timestamp 1698431365
transform 1 0 14336 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2255_
timestamp 1698431365
transform -1 0 16016 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2256_
timestamp 1698431365
transform -1 0 14224 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2257_
timestamp 1698431365
transform -1 0 13216 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2258_
timestamp 1698431365
transform -1 0 11872 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2259_
timestamp 1698431365
transform -1 0 11200 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2260_
timestamp 1698431365
transform 1 0 14224 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2261_
timestamp 1698431365
transform -1 0 14672 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2262_
timestamp 1698431365
transform 1 0 11984 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2263_
timestamp 1698431365
transform -1 0 12992 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2264_
timestamp 1698431365
transform -1 0 14560 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2265_
timestamp 1698431365
transform 1 0 13888 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2266_
timestamp 1698431365
transform -1 0 13888 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2267_
timestamp 1698431365
transform 1 0 11984 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2268_
timestamp 1698431365
transform -1 0 11200 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2269_
timestamp 1698431365
transform 1 0 9632 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2270_
timestamp 1698431365
transform -1 0 13664 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2271_
timestamp 1698431365
transform 1 0 12208 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2272_
timestamp 1698431365
transform -1 0 14336 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2273_
timestamp 1698431365
transform -1 0 14448 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2274_
timestamp 1698431365
transform 1 0 11536 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2275_
timestamp 1698431365
transform 1 0 11648 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2276_
timestamp 1698431365
transform -1 0 11200 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2277_
timestamp 1698431365
transform -1 0 10528 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2278_
timestamp 1698431365
transform -1 0 12992 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2279_
timestamp 1698431365
transform -1 0 11648 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2280_
timestamp 1698431365
transform 1 0 10080 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2281_
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2282_
timestamp 1698431365
transform -1 0 15008 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2283_
timestamp 1698431365
transform -1 0 16576 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2284_
timestamp 1698431365
transform -1 0 14896 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2285_
timestamp 1698431365
transform 1 0 12432 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2286_
timestamp 1698431365
transform 1 0 13552 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2287_
timestamp 1698431365
transform -1 0 16016 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2288_
timestamp 1698431365
transform -1 0 15232 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2289_
timestamp 1698431365
transform -1 0 12320 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2290_
timestamp 1698431365
transform 1 0 17360 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2291_
timestamp 1698431365
transform -1 0 27776 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2292_
timestamp 1698431365
transform -1 0 26656 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2293_
timestamp 1698431365
transform -1 0 26208 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2294_
timestamp 1698431365
transform -1 0 41664 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2295_
timestamp 1698431365
transform 1 0 39536 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2296_
timestamp 1698431365
transform 1 0 38864 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2297_
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2298_
timestamp 1698431365
transform -1 0 41664 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2299_
timestamp 1698431365
transform 1 0 39536 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2300_
timestamp 1698431365
transform 1 0 41664 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2301_
timestamp 1698431365
transform 1 0 41664 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2302_
timestamp 1698431365
transform 1 0 42112 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2303_
timestamp 1698431365
transform 1 0 43904 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2304_
timestamp 1698431365
transform -1 0 42784 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2305_
timestamp 1698431365
transform 1 0 46368 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2306_
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2307_
timestamp 1698431365
transform -1 0 46368 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2308_
timestamp 1698431365
transform -1 0 42224 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2309_
timestamp 1698431365
transform -1 0 40320 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2310_
timestamp 1698431365
transform 1 0 42560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2311_
timestamp 1698431365
transform 1 0 39424 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2312_
timestamp 1698431365
transform 1 0 39088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2313_
timestamp 1698431365
transform 1 0 41216 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2314_
timestamp 1698431365
transform 1 0 43344 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2315_
timestamp 1698431365
transform -1 0 43904 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2316_
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2317_
timestamp 1698431365
transform 1 0 40096 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2318_
timestamp 1698431365
transform 1 0 34944 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2319_
timestamp 1698431365
transform 1 0 38416 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2320_
timestamp 1698431365
transform -1 0 39536 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2321_
timestamp 1698431365
transform -1 0 37744 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2322_
timestamp 1698431365
transform -1 0 38080 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2323_
timestamp 1698431365
transform 1 0 38752 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2324_
timestamp 1698431365
transform 1 0 37856 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2325_
timestamp 1698431365
transform 1 0 39648 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2326_
timestamp 1698431365
transform 1 0 38416 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2327_
timestamp 1698431365
transform 1 0 36400 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2328_
timestamp 1698431365
transform 1 0 35616 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2329_
timestamp 1698431365
transform -1 0 39312 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2330_
timestamp 1698431365
transform 1 0 39200 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2331_
timestamp 1698431365
transform 1 0 7056 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2332_
timestamp 1698431365
transform -1 0 8176 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2333_
timestamp 1698431365
transform -1 0 34384 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2334_
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2335_
timestamp 1698431365
transform -1 0 22848 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2336_
timestamp 1698431365
transform -1 0 24192 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2337_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2338_
timestamp 1698431365
transform 1 0 21280 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2339_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2340_
timestamp 1698431365
transform 1 0 20048 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2341_
timestamp 1698431365
transform -1 0 23632 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2342_
timestamp 1698431365
transform 1 0 21952 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2343_
timestamp 1698431365
transform -1 0 22848 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2344_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2345_
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2346_
timestamp 1698431365
transform -1 0 44464 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2347_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2348_
timestamp 1698431365
transform -1 0 44464 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2349_
timestamp 1698431365
transform 1 0 43344 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2350_
timestamp 1698431365
transform 1 0 43904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2351_
timestamp 1698431365
transform 1 0 42336 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2352_
timestamp 1698431365
transform -1 0 42112 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2353_
timestamp 1698431365
transform -1 0 43792 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2354_
timestamp 1698431365
transform -1 0 43568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2355_
timestamp 1698431365
transform -1 0 42112 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2356_
timestamp 1698431365
transform -1 0 46480 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2357_
timestamp 1698431365
transform 1 0 45584 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2358_
timestamp 1698431365
transform 1 0 45360 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2359_
timestamp 1698431365
transform -1 0 46032 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2360_
timestamp 1698431365
transform -1 0 46928 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2361_
timestamp 1698431365
transform -1 0 48944 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2362_
timestamp 1698431365
transform -1 0 49056 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2363_
timestamp 1698431365
transform -1 0 48272 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2364_
timestamp 1698431365
transform -1 0 47824 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2365_
timestamp 1698431365
transform -1 0 47264 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2366_
timestamp 1698431365
transform -1 0 49056 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2367_
timestamp 1698431365
transform -1 0 34272 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2368_
timestamp 1698431365
transform -1 0 32704 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2369_
timestamp 1698431365
transform -1 0 30128 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2370_
timestamp 1698431365
transform 1 0 31024 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2371_
timestamp 1698431365
transform -1 0 34832 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2372_
timestamp 1698431365
transform 1 0 32144 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2373_
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2374_
timestamp 1698431365
transform 1 0 32704 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2375_
timestamp 1698431365
transform 1 0 31696 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2376_
timestamp 1698431365
transform 1 0 34048 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2377_
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2378_
timestamp 1698431365
transform -1 0 43904 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2379_
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2380_
timestamp 1698431365
transform -1 0 42896 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2381_
timestamp 1698431365
transform 1 0 43904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2382_
timestamp 1698431365
transform -1 0 43680 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2383_
timestamp 1698431365
transform -1 0 42784 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2384_
timestamp 1698431365
transform -1 0 41776 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2385_
timestamp 1698431365
transform -1 0 41216 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2386_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2387_
timestamp 1698431365
transform -1 0 6496 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2388_
timestamp 1698431365
transform 1 0 2128 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2389_
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2390_
timestamp 1698431365
transform 1 0 7504 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2391_
timestamp 1698431365
transform 1 0 6832 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2392_
timestamp 1698431365
transform 1 0 9744 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2393_
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2394_
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2395_
timestamp 1698431365
transform 1 0 2016 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2396_
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2397_
timestamp 1698431365
transform -1 0 12656 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2398_
timestamp 1698431365
transform -1 0 12432 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2399_
timestamp 1698431365
transform -1 0 9408 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2400_
timestamp 1698431365
transform -1 0 12768 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2401_
timestamp 1698431365
transform 1 0 9632 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2402_
timestamp 1698431365
transform 1 0 9632 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2403_
timestamp 1698431365
transform 1 0 5712 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2404_
timestamp 1698431365
transform -1 0 12320 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2405_
timestamp 1698431365
transform -1 0 9520 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2406_
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2407_
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2408_
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2409_
timestamp 1698431365
transform 1 0 5936 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2410_
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2411_
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2412_
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2413_
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2414_
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2415_
timestamp 1698431365
transform 1 0 2016 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2416_
timestamp 1698431365
transform 1 0 3136 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2417_
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2418_
timestamp 1698431365
transform 1 0 32144 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2419_
timestamp 1698431365
transform -1 0 36176 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2420_
timestamp 1698431365
transform 1 0 33376 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2421_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2422_
timestamp 1698431365
transform -1 0 40096 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2423_
timestamp 1698431365
transform -1 0 20496 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2424_
timestamp 1698431365
transform -1 0 20384 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2425_
timestamp 1698431365
transform 1 0 21504 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2426_
timestamp 1698431365
transform -1 0 24864 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2427_
timestamp 1698431365
transform 1 0 27328 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2428_
timestamp 1698431365
transform 1 0 27664 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2429_
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2430_
timestamp 1698431365
transform 1 0 24080 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2431_
timestamp 1698431365
transform 1 0 23184 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2432_
timestamp 1698431365
transform 1 0 19824 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2433_
timestamp 1698431365
transform -1 0 24304 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2434_
timestamp 1698431365
transform 1 0 17584 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2435_
timestamp 1698431365
transform -1 0 23968 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2436_
timestamp 1698431365
transform -1 0 38416 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2437_
timestamp 1698431365
transform 1 0 38528 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2438_
timestamp 1698431365
transform 1 0 40096 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2439_
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2440_
timestamp 1698431365
transform 1 0 43792 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2441_
timestamp 1698431365
transform 1 0 44688 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2442_
timestamp 1698431365
transform 1 0 45136 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2443_
timestamp 1698431365
transform 1 0 46144 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2444_
timestamp 1698431365
transform 1 0 46144 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2445_
timestamp 1698431365
transform 1 0 41216 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2446_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2447_
timestamp 1698431365
transform 1 0 23520 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2448_
timestamp 1698431365
transform 1 0 20272 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2449_
timestamp 1698431365
transform 1 0 17584 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2450_
timestamp 1698431365
transform 1 0 12992 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2451_
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2452_
timestamp 1698431365
transform 1 0 12880 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2453_
timestamp 1698431365
transform 1 0 16016 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2454_
timestamp 1698431365
transform -1 0 26432 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2455_
timestamp 1698431365
transform -1 0 27776 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2456_
timestamp 1698431365
transform -1 0 28784 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2457_
timestamp 1698431365
transform -1 0 25536 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2458_
timestamp 1698431365
transform -1 0 24416 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2459_
timestamp 1698431365
transform -1 0 24640 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2460_
timestamp 1698431365
transform -1 0 21952 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2461_
timestamp 1698431365
transform 1 0 18144 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2462_
timestamp 1698431365
transform 1 0 25536 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2463_
timestamp 1698431365
transform 1 0 25088 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2464_
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2465_
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2466_
timestamp 1698431365
transform 1 0 36176 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2467_
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2468_
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2469_
timestamp 1698431365
transform -1 0 38304 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2470_
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2471_
timestamp 1698431365
transform 1 0 29008 0 -1 39200
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2472_
timestamp 1698431365
transform 1 0 23856 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2473_
timestamp 1698431365
transform 1 0 24640 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2474_
timestamp 1698431365
transform 1 0 34160 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2475_
timestamp 1698431365
transform -1 0 37632 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2476_
timestamp 1698431365
transform 1 0 32592 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2477_
timestamp 1698431365
transform -1 0 33936 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2478_
timestamp 1698431365
transform 1 0 31136 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2479_
timestamp 1698431365
transform 1 0 21168 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2480_
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2481_
timestamp 1698431365
transform 1 0 16688 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2482_
timestamp 1698431365
transform 1 0 8512 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2483_
timestamp 1698431365
transform 1 0 8624 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2484_
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2485_
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2486_
timestamp 1698431365
transform 1 0 14336 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2487_
timestamp 1698431365
transform 1 0 5040 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2488_
timestamp 1698431365
transform 1 0 4368 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2489_
timestamp 1698431365
transform 1 0 5264 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2490_
timestamp 1698431365
transform 1 0 4928 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2491_
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2492_
timestamp 1698431365
transform 1 0 9856 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2493_
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2494_
timestamp 1698431365
transform -1 0 18704 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2495_
timestamp 1698431365
transform 1 0 23520 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2496_
timestamp 1698431365
transform 1 0 21392 0 -1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2497_
timestamp 1698431365
transform 1 0 40656 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2498_
timestamp 1698431365
transform -1 0 40656 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2499_
timestamp 1698431365
transform 1 0 39648 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2500_
timestamp 1698431365
transform 1 0 39088 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2501_
timestamp 1698431365
transform 1 0 37408 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2502_
timestamp 1698431365
transform 1 0 37184 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2503_
timestamp 1698431365
transform 1 0 37520 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2504_
timestamp 1698431365
transform 1 0 37296 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2505_
timestamp 1698431365
transform -1 0 28000 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2506_
timestamp 1698431365
transform -1 0 32256 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2507_
timestamp 1698431365
transform -1 0 24864 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2508_
timestamp 1698431365
transform -1 0 28336 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2509_
timestamp 1698431365
transform -1 0 24416 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2510_
timestamp 1698431365
transform -1 0 24864 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2511_
timestamp 1698431365
transform -1 0 20944 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2512_
timestamp 1698431365
transform -1 0 24416 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2513_
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2514_
timestamp 1698431365
transform -1 0 40096 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2515_
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2516_
timestamp 1698431365
transform 1 0 10640 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2517_
timestamp 1698431365
transform 1 0 23744 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2518_
timestamp 1698431365
transform 1 0 29792 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2519_
timestamp 1698431365
transform 1 0 26768 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2520_
timestamp 1698431365
transform 1 0 23856 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2521_
timestamp 1698431365
transform 1 0 29120 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2522_
timestamp 1698431365
transform 1 0 33040 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2523_
timestamp 1698431365
transform 1 0 42336 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2524_
timestamp 1698431365
transform 1 0 43232 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2525_
timestamp 1698431365
transform 1 0 46144 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2526_
timestamp 1698431365
transform 1 0 46144 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2527_
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2528_
timestamp 1698431365
transform 1 0 46144 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2529_
timestamp 1698431365
transform 1 0 46144 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2530_
timestamp 1698431365
transform -1 0 40432 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2531_
timestamp 1698431365
transform -1 0 43568 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2532_
timestamp 1698431365
transform 1 0 40768 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2533_
timestamp 1698431365
transform 1 0 41216 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2534_
timestamp 1698431365
transform -1 0 47936 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2535_
timestamp 1698431365
transform 1 0 46144 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2536_
timestamp 1698431365
transform 1 0 46144 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2537_
timestamp 1698431365
transform 1 0 46144 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2538_
timestamp 1698431365
transform 1 0 41776 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2539_
timestamp 1698431365
transform 1 0 46144 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2540_
timestamp 1698431365
transform 1 0 46144 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2541_
timestamp 1698431365
transform 1 0 46144 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2542_
timestamp 1698431365
transform -1 0 49392 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2543_
timestamp 1698431365
transform 1 0 44128 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2544_
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2545_
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2546_
timestamp 1698431365
transform 1 0 44464 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2547_
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2548_
timestamp 1698431365
transform -1 0 13216 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2549_
timestamp 1698431365
transform 1 0 9856 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2550_
timestamp 1698431365
transform -1 0 9072 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2551_
timestamp 1698431365
transform 1 0 7728 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2552_
timestamp 1698431365
transform 1 0 6608 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2553_
timestamp 1698431365
transform 1 0 5264 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2554_
timestamp 1698431365
transform 1 0 3696 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2555_
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2556_
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2557_
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2558_
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2559_
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2560_
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2561_
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2562_
timestamp 1698431365
transform -1 0 9072 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2563_
timestamp 1698431365
transform -1 0 10752 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2564_
timestamp 1698431365
transform -1 0 36624 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2565_
timestamp 1698431365
transform 1 0 32256 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2566_
timestamp 1698431365
transform -1 0 36176 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2567_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2568_
timestamp 1698431365
transform -1 0 40208 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2569_
timestamp 1698431365
transform -1 0 39424 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2570_
timestamp 1698431365
transform 1 0 46144 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2571_
timestamp 1698431365
transform 1 0 21392 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2572_
timestamp 1698431365
transform 1 0 20720 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2573_
timestamp 1698431365
transform 1 0 17472 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2574_
timestamp 1698431365
transform 1 0 13776 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2575_
timestamp 1698431365
transform 1 0 16240 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2576_
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2577_
timestamp 1698431365
transform 1 0 12320 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2578_
timestamp 1698431365
transform 1 0 12768 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2579_
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2580_
timestamp 1698431365
transform 1 0 12208 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2581_
timestamp 1698431365
transform 1 0 13328 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2582_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2583_
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2584_
timestamp 1698431365
transform 1 0 31696 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2585_
timestamp 1698431365
transform 1 0 33376 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2586_
timestamp 1698431365
transform -1 0 38416 0 -1 42336
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2587_
timestamp 1698431365
transform 1 0 34272 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2588_
timestamp 1698431365
transform 1 0 32032 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2589_
timestamp 1698431365
transform 1 0 28672 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2590_
timestamp 1698431365
transform 1 0 23632 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2591_
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2592_
timestamp 1698431365
transform -1 0 32256 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2593_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2594_
timestamp 1698431365
transform 1 0 24416 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2595_
timestamp 1698431365
transform 1 0 27216 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2596_
timestamp 1698431365
transform -1 0 33824 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2597_
timestamp 1698431365
transform 1 0 21168 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2598_
timestamp 1698431365
transform 1 0 20496 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2599_
timestamp 1698431365
transform 1 0 13776 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2600_
timestamp 1698431365
transform 1 0 9520 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2601_
timestamp 1698431365
transform -1 0 13328 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2602_
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2603_
timestamp 1698431365
transform 1 0 12432 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2604_
timestamp 1698431365
transform 1 0 8960 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2605_
timestamp 1698431365
transform 1 0 9856 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2606_
timestamp 1698431365
transform 1 0 13216 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2607_
timestamp 1698431365
transform 1 0 10864 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2608_
timestamp 1698431365
transform 1 0 14000 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2609_
timestamp 1698431365
transform 1 0 23632 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2610_
timestamp 1698431365
transform 1 0 39312 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2611_
timestamp 1698431365
transform 1 0 38528 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2612_
timestamp 1698431365
transform -1 0 44464 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2613_
timestamp 1698431365
transform -1 0 46032 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2614_
timestamp 1698431365
transform 1 0 38080 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2615_
timestamp 1698431365
transform 1 0 37296 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2616_
timestamp 1698431365
transform -1 0 45696 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2617_
timestamp 1698431365
transform 1 0 35616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2618_
timestamp 1698431365
transform 1 0 33376 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2619_
timestamp 1698431365
transform -1 0 40544 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2620_
timestamp 1698431365
transform 1 0 33376 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2621_
timestamp 1698431365
transform 1 0 37296 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2622_
timestamp 1698431365
transform 1 0 5936 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2623_
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2624_
timestamp 1698431365
transform -1 0 21280 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2625_
timestamp 1698431365
transform -1 0 24416 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2626_
timestamp 1698431365
transform -1 0 22176 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2627_
timestamp 1698431365
transform -1 0 45584 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2628_
timestamp 1698431365
transform 1 0 39088 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2629_
timestamp 1698431365
transform -1 0 43792 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2630_
timestamp 1698431365
transform -1 0 45360 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2631_
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2632_
timestamp 1698431365
transform 1 0 46144 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2633_
timestamp 1698431365
transform 1 0 46144 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2634_
timestamp 1698431365
transform 1 0 46032 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2635_
timestamp 1698431365
transform 1 0 30016 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2636_
timestamp 1698431365
transform -1 0 29904 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2637_
timestamp 1698431365
transform 1 0 32480 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2638_
timestamp 1698431365
transform 1 0 29008 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2639_
timestamp 1698431365
transform -1 0 46368 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2640_
timestamp 1698431365
transform -1 0 45360 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2641_
timestamp 1698431365
transform 1 0 41216 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2642_
timestamp 1698431365
transform 1 0 39424 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1191__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14896 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__A1
timestamp 1698431365
transform 1 0 14448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__A2
timestamp 1698431365
transform 1 0 20944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1203__B2
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__A2
timestamp 1698431365
transform 1 0 28784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__A1
timestamp 1698431365
transform 1 0 28336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__B1
timestamp 1698431365
transform -1 0 27328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__I
timestamp 1698431365
transform 1 0 18032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1214__A1
timestamp 1698431365
transform 1 0 26096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1214__B1
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A3
timestamp 1698431365
transform 1 0 37072 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__A2
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__I
timestamp 1698431365
transform 1 0 9072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1294__B
timestamp 1698431365
transform 1 0 8400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1307__B
timestamp 1698431365
transform 1 0 6608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__I
timestamp 1698431365
transform 1 0 49168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1350__I
timestamp 1698431365
transform 1 0 29120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A3
timestamp 1698431365
transform -1 0 36176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A4
timestamp 1698431365
transform -1 0 35616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1355__I
timestamp 1698431365
transform 1 0 34608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__I
timestamp 1698431365
transform 1 0 39200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__A1
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1360__A1
timestamp 1698431365
transform 1 0 38416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__I
timestamp 1698431365
transform -1 0 28672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A1
timestamp 1698431365
transform 1 0 30240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1365__I
timestamp 1698431365
transform -1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__A1
timestamp 1698431365
transform 1 0 33152 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__I
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1369__A1
timestamp 1698431365
transform 1 0 41664 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__A1
timestamp 1698431365
transform 1 0 38864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1374__I
timestamp 1698431365
transform 1 0 21056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1380__I
timestamp 1698431365
transform 1 0 20048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1384__A1
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__I
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1387__A1
timestamp 1698431365
transform -1 0 19040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__I
timestamp 1698431365
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1391__I
timestamp 1698431365
transform -1 0 31024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A2
timestamp 1698431365
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__I
timestamp 1698431365
transform 1 0 39648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1396__A1
timestamp 1698431365
transform 1 0 22288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__B
timestamp 1698431365
transform -1 0 21728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__I
timestamp 1698431365
transform 1 0 36400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A1
timestamp 1698431365
transform -1 0 15120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1413__I
timestamp 1698431365
transform 1 0 27104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A1
timestamp 1698431365
transform -1 0 18928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1419__A1
timestamp 1698431365
transform 1 0 23296 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1424__A1
timestamp 1698431365
transform 1 0 23968 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1432__B
timestamp 1698431365
transform -1 0 23072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__A1
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A1
timestamp 1698431365
transform 1 0 22400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1445__A1
timestamp 1698431365
transform -1 0 6608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1455__I
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__I
timestamp 1698431365
transform 1 0 23520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__I
timestamp 1698431365
transform -1 0 4368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1459__I
timestamp 1698431365
transform -1 0 4928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__A1
timestamp 1698431365
transform -1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__A1
timestamp 1698431365
transform 1 0 12544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1465__A1
timestamp 1698431365
transform 1 0 9856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__I
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A1
timestamp 1698431365
transform 1 0 8736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1470__I
timestamp 1698431365
transform -1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__B1
timestamp 1698431365
transform -1 0 4816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1499__A1
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A1
timestamp 1698431365
transform 1 0 12880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__I
timestamp 1698431365
transform 1 0 27888 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A1
timestamp 1698431365
transform 1 0 25760 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1698431365
transform 1 0 25312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1510__A1
timestamp 1698431365
transform 1 0 28224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__A1
timestamp 1698431365
transform 1 0 27104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__A1
timestamp 1698431365
transform 1 0 28112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A1
timestamp 1698431365
transform 1 0 28112 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1518__I
timestamp 1698431365
transform -1 0 24416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A1
timestamp 1698431365
transform 1 0 23520 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__I
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__A1
timestamp 1698431365
transform -1 0 21728 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A1
timestamp 1698431365
transform 1 0 21616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A1
timestamp 1698431365
transform -1 0 22400 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__I
timestamp 1698431365
transform -1 0 31472 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1545__A1
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__I
timestamp 1698431365
transform 1 0 41440 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__A1
timestamp 1698431365
transform 1 0 29904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__A2
timestamp 1698431365
transform 1 0 30576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1550__A1
timestamp 1698431365
transform -1 0 36512 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A1
timestamp 1698431365
transform -1 0 34384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1554__A1
timestamp 1698431365
transform 1 0 32928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A1
timestamp 1698431365
transform -1 0 37184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__I
timestamp 1698431365
transform 1 0 28560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1560__A1
timestamp 1698431365
transform 1 0 30800 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A1
timestamp 1698431365
transform 1 0 28784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__A1
timestamp 1698431365
transform 1 0 25872 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A1
timestamp 1698431365
transform 1 0 26880 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1569__A1
timestamp 1698431365
transform -1 0 26768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A1
timestamp 1698431365
transform -1 0 10528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1604__A1
timestamp 1698431365
transform -1 0 6048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A2
timestamp 1698431365
transform 1 0 5264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__A2
timestamp 1698431365
transform -1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A1
timestamp 1698431365
transform 1 0 6048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A1
timestamp 1698431365
transform 1 0 6048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__I
timestamp 1698431365
transform -1 0 30688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1640__I
timestamp 1698431365
transform 1 0 38864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__A1
timestamp 1698431365
transform 1 0 42896 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__A2
timestamp 1698431365
transform 1 0 40992 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__A1
timestamp 1698431365
transform 1 0 45920 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A1
timestamp 1698431365
transform 1 0 42000 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__A1
timestamp 1698431365
transform 1 0 39312 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A1
timestamp 1698431365
transform 1 0 46704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I
timestamp 1698431365
transform -1 0 38416 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A1
timestamp 1698431365
transform -1 0 37520 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__A1
timestamp 1698431365
transform 1 0 39760 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__A1
timestamp 1698431365
transform -1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A1
timestamp 1698431365
transform -1 0 39312 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__I
timestamp 1698431365
transform 1 0 42560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A1
timestamp 1698431365
transform -1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1698431365
transform 1 0 28224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__I
timestamp 1698431365
transform 1 0 45808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A1
timestamp 1698431365
transform -1 0 30464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__I
timestamp 1698431365
transform -1 0 41328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__A1
timestamp 1698431365
transform -1 0 29456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__I
timestamp 1698431365
transform -1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__A1
timestamp 1698431365
transform -1 0 28672 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A1
timestamp 1698431365
transform 1 0 24640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A1
timestamp 1698431365
transform -1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A1
timestamp 1698431365
transform 1 0 20944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A1
timestamp 1698431365
transform 1 0 25872 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A1
timestamp 1698431365
transform -1 0 15344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A2
timestamp 1698431365
transform 1 0 6496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__C
timestamp 1698431365
transform -1 0 5264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__A1
timestamp 1698431365
transform 1 0 12208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__A2
timestamp 1698431365
transform -1 0 12880 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__A1
timestamp 1698431365
transform -1 0 30240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A1
timestamp 1698431365
transform 1 0 32592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__A1
timestamp 1698431365
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__A1
timestamp 1698431365
transform 1 0 32032 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__A1
timestamp 1698431365
transform 1 0 29232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A1
timestamp 1698431365
transform 1 0 35504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A1
timestamp 1698431365
transform -1 0 36176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A1
timestamp 1698431365
transform -1 0 32928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__I
timestamp 1698431365
transform -1 0 16128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__B1
timestamp 1698431365
transform -1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__A1
timestamp 1698431365
transform 1 0 30688 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__A1
timestamp 1698431365
transform -1 0 31808 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__A2
timestamp 1698431365
transform 1 0 30688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A2
timestamp 1698431365
transform 1 0 39424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__A1
timestamp 1698431365
transform 1 0 42448 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__A2
timestamp 1698431365
transform 1 0 45360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A1
timestamp 1698431365
transform 1 0 37744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__A1
timestamp 1698431365
transform -1 0 34272 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__A1
timestamp 1698431365
transform 1 0 39984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__A1
timestamp 1698431365
transform -1 0 12320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__A1
timestamp 1698431365
transform 1 0 11312 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__A1
timestamp 1698431365
transform -1 0 9856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__I
timestamp 1698431365
transform -1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__B
timestamp 1698431365
transform 1 0 13552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__B
timestamp 1698431365
transform -1 0 12768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__B
timestamp 1698431365
transform -1 0 8176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__B
timestamp 1698431365
transform -1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__C
timestamp 1698431365
transform 1 0 10640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__A2
timestamp 1698431365
transform -1 0 10080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__A1
timestamp 1698431365
transform -1 0 28112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__A2
timestamp 1698431365
transform -1 0 22624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A1
timestamp 1698431365
transform 1 0 21952 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A1
timestamp 1698431365
transform 1 0 30688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A2
timestamp 1698431365
transform 1 0 31136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A2
timestamp 1698431365
transform -1 0 19376 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__I
timestamp 1698431365
transform 1 0 27104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A2
timestamp 1698431365
transform -1 0 21616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__B1
timestamp 1698431365
transform -1 0 20496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__I
timestamp 1698431365
transform -1 0 18704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__A2
timestamp 1698431365
transform 1 0 30912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__B
timestamp 1698431365
transform -1 0 31360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2044__A3
timestamp 1698431365
transform -1 0 26880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2044__A4
timestamp 1698431365
transform 1 0 28448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A2
timestamp 1698431365
transform 1 0 24528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__I
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2086__A1
timestamp 1698431365
transform 1 0 19264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2086__A2
timestamp 1698431365
transform 1 0 19712 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2086__C
timestamp 1698431365
transform 1 0 19824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__A1
timestamp 1698431365
transform 1 0 29232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__A2
timestamp 1698431365
transform 1 0 30352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__A3
timestamp 1698431365
transform 1 0 29792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2089__B
timestamp 1698431365
transform 1 0 31584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__A2
timestamp 1698431365
transform 1 0 31136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2143__A2
timestamp 1698431365
transform 1 0 30464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2143__B
timestamp 1698431365
transform -1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__A3
timestamp 1698431365
transform 1 0 33936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__A4
timestamp 1698431365
transform 1 0 42112 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2148__A2
timestamp 1698431365
transform -1 0 33824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__A1
timestamp 1698431365
transform -1 0 28224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__A2
timestamp 1698431365
transform 1 0 29680 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__C
timestamp 1698431365
transform -1 0 27776 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__A2
timestamp 1698431365
transform 1 0 32592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__A2
timestamp 1698431365
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__A3
timestamp 1698431365
transform 1 0 33040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__B
timestamp 1698431365
transform 1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A2
timestamp 1698431365
transform -1 0 22512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2245__A2
timestamp 1698431365
transform 1 0 30688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2245__B
timestamp 1698431365
transform 1 0 32032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__A3
timestamp 1698431365
transform 1 0 26656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__A4
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2250__A2
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A1
timestamp 1698431365
transform -1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A2
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__C
timestamp 1698431365
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A2
timestamp 1698431365
transform 1 0 25312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__A2
timestamp 1698431365
transform -1 0 25088 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__A3
timestamp 1698431365
transform -1 0 25536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2293__B
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2295__A2
timestamp 1698431365
transform -1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2302__A1
timestamp 1698431365
transform -1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2304__B
timestamp 1698431365
transform -1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__B
timestamp 1698431365
transform 1 0 6608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A1
timestamp 1698431365
transform -1 0 10080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2316__A4
timestamp 1698431365
transform 1 0 43344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2317__A1
timestamp 1698431365
transform 1 0 26544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2317__A2
timestamp 1698431365
transform 1 0 40768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__A1
timestamp 1698431365
transform -1 0 18032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__A2
timestamp 1698431365
transform -1 0 23968 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__B
timestamp 1698431365
transform 1 0 14112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__A1
timestamp 1698431365
transform -1 0 11200 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2325__A1
timestamp 1698431365
transform -1 0 9296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2327__A1
timestamp 1698431365
transform 1 0 35056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__A1
timestamp 1698431365
transform -1 0 26320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2331__A1
timestamp 1698431365
transform -1 0 8848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2331__A2
timestamp 1698431365
transform 1 0 8400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2344__A1
timestamp 1698431365
transform -1 0 21168 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__A1
timestamp 1698431365
transform -1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__A1
timestamp 1698431365
transform 1 0 47152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__A1
timestamp 1698431365
transform 1 0 45920 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A1
timestamp 1698431365
transform 1 0 42896 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2355__A1
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2359__A1
timestamp 1698431365
transform -1 0 26544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2361__A1
timestamp 1698431365
transform -1 0 29792 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__A1
timestamp 1698431365
transform -1 0 24416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A1
timestamp 1698431365
transform -1 0 25872 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__A1
timestamp 1698431365
transform -1 0 23520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2384__A1
timestamp 1698431365
transform -1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 23856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 18704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 20720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 34720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 34608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 19376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_1_wb_clk_i_I
timestamp 1698431365
transform 1 0 20944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_2_wb_clk_i_I
timestamp 1698431365
transform 1 0 18032 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_3_wb_clk_i_I
timestamp 1698431365
transform -1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_4_wb_clk_i_I
timestamp 1698431365
transform 1 0 9184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_5_wb_clk_i_I
timestamp 1698431365
transform 1 0 16688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_6_wb_clk_i_I
timestamp 1698431365
transform 1 0 8624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_7_wb_clk_i_I
timestamp 1698431365
transform 1 0 12656 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_8_wb_clk_i_I
timestamp 1698431365
transform 1 0 17472 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_9_wb_clk_i_I
timestamp 1698431365
transform -1 0 18816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_10_wb_clk_i_I
timestamp 1698431365
transform 1 0 23072 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_11_wb_clk_i_I
timestamp 1698431365
transform 1 0 20944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_12_wb_clk_i_I
timestamp 1698431365
transform 1 0 24640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_13_wb_clk_i_I
timestamp 1698431365
transform 1 0 40320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_14_wb_clk_i_I
timestamp 1698431365
transform 1 0 34832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_15_wb_clk_i_I
timestamp 1698431365
transform -1 0 36960 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_16_wb_clk_i_I
timestamp 1698431365
transform 1 0 48048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_17_wb_clk_i_I
timestamp 1698431365
transform -1 0 41104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_18_wb_clk_i_I
timestamp 1698431365
transform 1 0 45808 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_19_wb_clk_i_I
timestamp 1698431365
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_20_wb_clk_i_I
timestamp 1698431365
transform -1 0 41888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_21_wb_clk_i_I
timestamp 1698431365
transform 1 0 45808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_22_wb_clk_i_I
timestamp 1698431365
transform 1 0 41440 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_23_wb_clk_i_I
timestamp 1698431365
transform -1 0 38976 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_24_wb_clk_i_I
timestamp 1698431365
transform 1 0 22176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_25_wb_clk_i_I
timestamp 1698431365
transform 1 0 40992 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_26_wb_clk_i_I
timestamp 1698431365
transform -1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_27_wb_clk_i_I
timestamp 1698431365
transform 1 0 5040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_28_wb_clk_i_I
timestamp 1698431365
transform -1 0 4816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_29_wb_clk_i_I
timestamp 1698431365
transform 1 0 8512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_30_wb_clk_i_I
timestamp 1698431365
transform 1 0 6720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_31_wb_clk_i_I
timestamp 1698431365
transform 1 0 11760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_32_wb_clk_i_I
timestamp 1698431365
transform 1 0 38752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_33_wb_clk_i_I
timestamp 1698431365
transform 1 0 24416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_34_wb_clk_i_I
timestamp 1698431365
transform 1 0 20496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_35_wb_clk_i_I
timestamp 1698431365
transform 1 0 16016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_36_wb_clk_i_I
timestamp 1698431365
transform 1 0 10752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_37_wb_clk_i_I
timestamp 1698431365
transform 1 0 19152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_38_wb_clk_i_I
timestamp 1698431365
transform 1 0 6272 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_39_wb_clk_i_I
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_40_wb_clk_i_I
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_41_wb_clk_i_I
timestamp 1698431365
transform 1 0 10192 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_42_wb_clk_i_I
timestamp 1698431365
transform 1 0 11312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 49280 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 38864 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 33824 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 6720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 6384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 4816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 17136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 18592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 48272 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 46368 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 41552 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 30912 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 40656 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 19152 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1698431365
transform -1 0 20832 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1698431365
transform -1 0 20832 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1698431365
transform 1 0 34944 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 34944 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1698431365
transform -1 0 26768 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1698431365
transform 1 0 13440 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1698431365
transform -1 0 12432 0 1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1698431365
transform -1 0 9072 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1698431365
transform -1 0 15008 0 -1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1698431365
transform -1 0 7504 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1698431365
transform -1 0 12432 0 1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1698431365
transform -1 0 17024 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1698431365
transform -1 0 24416 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1698431365
transform 1 0 21392 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1698431365
transform -1 0 38528 0 -1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1698431365
transform -1 0 34608 0 1 39200
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1698431365
transform -1 0 36624 0 1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1698431365
transform -1 0 43792 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1698431365
transform -1 0 48384 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1698431365
transform -1 0 47488 0 -1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_21_wb_clk_i
timestamp 1698431365
transform -1 0 46368 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_22_wb_clk_i
timestamp 1698431365
transform -1 0 40544 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_23_wb_clk_i
timestamp 1698431365
transform -1 0 36512 0 1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_24_wb_clk_i
timestamp 1698431365
transform -1 0 42448 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_25_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_26_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_27_wb_clk_i
timestamp 1698431365
transform 1 0 42784 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_28_wb_clk_i
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_29_wb_clk_i
timestamp 1698431365
transform -1 0 43344 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_30_wb_clk_i
timestamp 1698431365
transform -1 0 38528 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_31_wb_clk_i
timestamp 1698431365
transform -1 0 38528 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_32_wb_clk_i
timestamp 1698431365
transform -1 0 36624 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_33_wb_clk_i
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_34_wb_clk_i
timestamp 1698431365
transform -1 0 26768 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_35_wb_clk_i
timestamp 1698431365
transform 1 0 23184 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_36_wb_clk_i
timestamp 1698431365
transform -1 0 22848 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_37_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_38_wb_clk_i
timestamp 1698431365
transform -1 0 15008 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_39_wb_clk_i
timestamp 1698431365
transform -1 0 11088 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_40_wb_clk_i
timestamp 1698431365
transform -1 0 15232 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_41_wb_clk_i
timestamp 1698431365
transform -1 0 8064 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_42_wb_clk_i
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_6 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_14 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2912 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_19
timestamp 1698431365
transform 1 0 3472 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_27 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_31
timestamp 1698431365
transform 1 0 4816 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_40
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_44
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_51
timestamp 1698431365
transform 1 0 7056 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_86
timestamp 1698431365
transform 1 0 10976 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_99
timestamp 1698431365
transform 1 0 12432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_109
timestamp 1698431365
transform 1 0 13552 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698431365
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_235
timestamp 1698431365
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_244
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_337
timestamp 1698431365
transform 1 0 39088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_378
timestamp 1698431365
transform 1 0 43680 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_420
timestamp 1698431365
transform 1 0 48384 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_18
timestamp 1698431365
transform 1 0 3360 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_26
timestamp 1698431365
transform 1 0 4256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_67
timestamp 1698431365
transform 1 0 8848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_101
timestamp 1698431365
transform 1 0 12656 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_110
timestamp 1698431365
transform 1 0 13664 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_173
timestamp 1698431365
transform 1 0 20720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_175
timestamp 1698431365
transform 1 0 20944 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_231
timestamp 1698431365
transform 1 0 27216 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_273
timestamp 1698431365
transform 1 0 31920 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_286
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_348
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_428
timestamp 1698431365
transform 1 0 49280 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_18
timestamp 1698431365
transform 1 0 3360 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_26
timestamp 1698431365
transform 1 0 4256 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_30
timestamp 1698431365
transform 1 0 4704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_32
timestamp 1698431365
transform 1 0 4928 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_41
timestamp 1698431365
transform 1 0 5936 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_44
timestamp 1698431365
transform 1 0 6272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_64
timestamp 1698431365
transform 1 0 8512 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_155
timestamp 1698431365
transform 1 0 18704 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_242
timestamp 1698431365
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_256
timestamp 1698431365
transform 1 0 30016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_384
timestamp 1698431365
transform 1 0 44352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_420
timestamp 1698431365
transform 1 0 48384 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_18
timestamp 1698431365
transform 1 0 3360 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_22
timestamp 1698431365
transform 1 0 3808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_24
timestamp 1698431365
transform 1 0 4032 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_27
timestamp 1698431365
transform 1 0 4368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_31
timestamp 1698431365
transform 1 0 4816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_122
timestamp 1698431365
transform 1 0 15008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_124
timestamp 1698431365
transform 1 0 15232 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_222
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_232
timestamp 1698431365
transform 1 0 27328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_234
timestamp 1698431365
transform 1 0 27552 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_264
timestamp 1698431365
transform 1 0 30912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_266
timestamp 1698431365
transform 1 0 31136 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_348
timestamp 1698431365
transform 1 0 40320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_417
timestamp 1698431365
transform 1 0 48048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_419
timestamp 1698431365
transform 1 0 48272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_428
timestamp 1698431365
transform 1 0 49280 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_18
timestamp 1698431365
transform 1 0 3360 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_26
timestamp 1698431365
transform 1 0 4256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_28
timestamp 1698431365
transform 1 0 4480 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_31
timestamp 1698431365
transform 1 0 4816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_39
timestamp 1698431365
transform 1 0 5712 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_42
timestamp 1698431365
transform 1 0 6048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_46
timestamp 1698431365
transform 1 0 6496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_64
timestamp 1698431365
transform 1 0 8512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_115
timestamp 1698431365
transform 1 0 14224 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_192
timestamp 1698431365
transform 1 0 22848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_194
timestamp 1698431365
transform 1 0 23072 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_303
timestamp 1698431365
transform 1 0 35280 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_321
timestamp 1698431365
transform 1 0 37296 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_370
timestamp 1698431365
transform 1 0 42784 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_384
timestamp 1698431365
transform 1 0 44352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_18
timestamp 1698431365
transform 1 0 3360 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_26
timestamp 1698431365
transform 1 0 4256 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_64
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_220
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_272
timestamp 1698431365
transform 1 0 31808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_347
timestamp 1698431365
transform 1 0 40208 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_349
timestamp 1698431365
transform 1 0 40432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_428
timestamp 1698431365
transform 1 0 49280 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_18
timestamp 1698431365
transform 1 0 3360 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_26
timestamp 1698431365
transform 1 0 4256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_30
timestamp 1698431365
transform 1 0 4704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_41
timestamp 1698431365
transform 1 0 5936 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_44
timestamp 1698431365
transform 1 0 6272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_70
timestamp 1698431365
transform 1 0 9184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_109
timestamp 1698431365
transform 1 0 13552 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_128
timestamp 1698431365
transform 1 0 15680 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_130
timestamp 1698431365
transform 1 0 15904 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_168
timestamp 1698431365
transform 1 0 20160 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_189
timestamp 1698431365
transform 1 0 22512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_230
timestamp 1698431365
transform 1 0 27104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_232
timestamp 1698431365
transform 1 0 27328 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_273
timestamp 1698431365
transform 1 0 31920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_286
timestamp 1698431365
transform 1 0 33376 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_288
timestamp 1698431365
transform 1 0 33600 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_328
timestamp 1698431365
transform 1 0 38080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_18
timestamp 1698431365
transform 1 0 3360 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_26
timestamp 1698431365
transform 1 0 4256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_30
timestamp 1698431365
transform 1 0 4704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_32
timestamp 1698431365
transform 1 0 4928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_62
timestamp 1698431365
transform 1 0 8288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_78
timestamp 1698431365
transform 1 0 10080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_82
timestamp 1698431365
transform 1 0 10528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_94
timestamp 1698431365
transform 1 0 11872 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_98
timestamp 1698431365
transform 1 0 12320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_113
timestamp 1698431365
transform 1 0 14000 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_119
timestamp 1698431365
transform 1 0 14672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_129
timestamp 1698431365
transform 1 0 15792 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_148
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_163
timestamp 1698431365
transform 1 0 19600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_165
timestamp 1698431365
transform 1 0 19824 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_175
timestamp 1698431365
transform 1 0 20944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_177
timestamp 1698431365
transform 1 0 21168 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_184
timestamp 1698431365
transform 1 0 21952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_226
timestamp 1698431365
transform 1 0 26656 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_232
timestamp 1698431365
transform 1 0 27328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_234
timestamp 1698431365
transform 1 0 27552 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_259
timestamp 1698431365
transform 1 0 30352 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_284
timestamp 1698431365
transform 1 0 33152 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_332
timestamp 1698431365
transform 1 0 38528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_336
timestamp 1698431365
transform 1 0 38976 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_345
timestamp 1698431365
transform 1 0 39984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_347
timestamp 1698431365
transform 1 0 40208 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_354
timestamp 1698431365
transform 1 0 40992 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_365
timestamp 1698431365
transform 1 0 42224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_367
timestamp 1698431365
transform 1 0 42448 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_399
timestamp 1698431365
transform 1 0 46032 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_419
timestamp 1698431365
transform 1 0 48272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_428
timestamp 1698431365
transform 1 0 49280 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_18
timestamp 1698431365
transform 1 0 3360 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_26
timestamp 1698431365
transform 1 0 4256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_28
timestamp 1698431365
transform 1 0 4480 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_31
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_41
timestamp 1698431365
transform 1 0 5936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_63
timestamp 1698431365
transform 1 0 8400 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_114
timestamp 1698431365
transform 1 0 14112 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_118
timestamp 1698431365
transform 1 0 14560 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_121
timestamp 1698431365
transform 1 0 14896 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_135
timestamp 1698431365
transform 1 0 16464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_179
timestamp 1698431365
transform 1 0 21392 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_212
timestamp 1698431365
transform 1 0 25088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_228
timestamp 1698431365
transform 1 0 26880 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_308
timestamp 1698431365
transform 1 0 35840 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_327
timestamp 1698431365
transform 1 0 37968 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_383
timestamp 1698431365
transform 1 0 44240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_395
timestamp 1698431365
transform 1 0 45584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_399
timestamp 1698431365
transform 1 0 46032 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_42
timestamp 1698431365
transform 1 0 6048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_44
timestamp 1698431365
transform 1 0 6272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_96
timestamp 1698431365
transform 1 0 12096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_100
timestamp 1698431365
transform 1 0 12544 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_173
timestamp 1698431365
transform 1 0 20720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_264
timestamp 1698431365
transform 1 0 30912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_290
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_317
timestamp 1698431365
transform 1 0 36848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_354
timestamp 1698431365
transform 1 0 40992 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_428
timestamp 1698431365
transform 1 0 49280 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_31
timestamp 1698431365
transform 1 0 4816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_87
timestamp 1698431365
transform 1 0 11088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_91
timestamp 1698431365
transform 1 0 11536 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_95
timestamp 1698431365
transform 1 0 11984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_157
timestamp 1698431365
transform 1 0 18928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_161
timestamp 1698431365
transform 1 0 19376 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_179
timestamp 1698431365
transform 1 0 21392 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_182
timestamp 1698431365
transform 1 0 21728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_186
timestamp 1698431365
transform 1 0 22176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_190
timestamp 1698431365
transform 1 0 22624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_194
timestamp 1698431365
transform 1 0 23072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_235
timestamp 1698431365
transform 1 0 27664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_255
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_285
timestamp 1698431365
transform 1 0 33264 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_10
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_14
timestamp 1698431365
transform 1 0 2912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_16
timestamp 1698431365
transform 1 0 3136 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698431365
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_82
timestamp 1698431365
transform 1 0 10528 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_112
timestamp 1698431365
transform 1 0 13888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_152
timestamp 1698431365
transform 1 0 18368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_154
timestamp 1698431365
transform 1 0 18592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_171
timestamp 1698431365
transform 1 0 20496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_175
timestamp 1698431365
transform 1 0 20944 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_198
timestamp 1698431365
transform 1 0 23520 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_222
timestamp 1698431365
transform 1 0 26208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_255
timestamp 1698431365
transform 1 0 29904 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_394
timestamp 1698431365
transform 1 0 45472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_428
timestamp 1698431365
transform 1 0 49280 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_31
timestamp 1698431365
transform 1 0 4816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_84
timestamp 1698431365
transform 1 0 10752 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_144
timestamp 1698431365
transform 1 0 17472 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_179
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_186
timestamp 1698431365
transform 1 0 22176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_227
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_229
timestamp 1698431365
transform 1 0 26992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_307
timestamp 1698431365
transform 1 0 35728 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_331
timestamp 1698431365
transform 1 0 38416 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_384
timestamp 1698431365
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_10
timestamp 1698431365
transform 1 0 2464 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_14
timestamp 1698431365
transform 1 0 2912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_33
timestamp 1698431365
transform 1 0 5040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_35
timestamp 1698431365
transform 1 0 5264 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_58
timestamp 1698431365
transform 1 0 7840 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_96
timestamp 1698431365
transform 1 0 12096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_103
timestamp 1698431365
transform 1 0 12880 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_133
timestamp 1698431365
transform 1 0 16240 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_137
timestamp 1698431365
transform 1 0 16688 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_158
timestamp 1698431365
transform 1 0 19040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_160
timestamp 1698431365
transform 1 0 19264 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_222
timestamp 1698431365
transform 1 0 26208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_224
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_233
timestamp 1698431365
transform 1 0 27440 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_239
timestamp 1698431365
transform 1 0 28112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_243
timestamp 1698431365
transform 1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_302
timestamp 1698431365
transform 1 0 35168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_428
timestamp 1698431365
transform 1 0 49280 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_31
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_54
timestamp 1698431365
transform 1 0 7392 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_58
timestamp 1698431365
transform 1 0 7840 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_67
timestamp 1698431365
transform 1 0 8848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_140
timestamp 1698431365
transform 1 0 17024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_144
timestamp 1698431365
transform 1 0 17472 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_146
timestamp 1698431365
transform 1 0 17696 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_155
timestamp 1698431365
transform 1 0 18704 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_277
timestamp 1698431365
transform 1 0 32368 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_307
timestamp 1698431365
transform 1 0 35728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_350
timestamp 1698431365
transform 1 0 40544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_354
timestamp 1698431365
transform 1 0 40992 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_53
timestamp 1698431365
transform 1 0 7280 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_55
timestamp 1698431365
transform 1 0 7504 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_132
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_134
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698431365
transform 1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_148
timestamp 1698431365
transform 1 0 17920 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_159
timestamp 1698431365
transform 1 0 19152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_163
timestamp 1698431365
transform 1 0 19600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_169
timestamp 1698431365
transform 1 0 20272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_219
timestamp 1698431365
transform 1 0 25872 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_315
timestamp 1698431365
transform 1 0 36624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_347
timestamp 1698431365
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_39
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_69
timestamp 1698431365
transform 1 0 9072 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_98
timestamp 1698431365
transform 1 0 12320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_115
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_134
timestamp 1698431365
transform 1 0 16352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_136
timestamp 1698431365
transform 1 0 16576 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_184
timestamp 1698431365
transform 1 0 21952 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_196
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_229
timestamp 1698431365
transform 1 0 26992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_251
timestamp 1698431365
transform 1 0 29456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_255
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_258
timestamp 1698431365
transform 1 0 30240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_262
timestamp 1698431365
transform 1 0 30688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_264
timestamp 1698431365
transform 1 0 30912 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_427
timestamp 1698431365
transform 1 0 49168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_135
timestamp 1698431365
transform 1 0 16464 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_144
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_192
timestamp 1698431365
transform 1 0 22848 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_198
timestamp 1698431365
transform 1 0 23520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_202
timestamp 1698431365
transform 1 0 23968 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_220
timestamp 1698431365
transform 1 0 25984 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_223
timestamp 1698431365
transform 1 0 26320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_260
timestamp 1698431365
transform 1 0 30464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_266
timestamp 1698431365
transform 1 0 31136 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_303
timestamp 1698431365
transform 1 0 35280 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_428
timestamp 1698431365
transform 1 0 49280 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_31
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_39
timestamp 1698431365
transform 1 0 5712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_96
timestamp 1698431365
transform 1 0 12096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_98
timestamp 1698431365
transform 1 0 12320 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_165
timestamp 1698431365
transform 1 0 19824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_199
timestamp 1698431365
transform 1 0 23632 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_230
timestamp 1698431365
transform 1 0 27104 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_253
timestamp 1698431365
transform 1 0 29680 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_298
timestamp 1698431365
transform 1 0 34720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_312
timestamp 1698431365
transform 1 0 36288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_339
timestamp 1698431365
transform 1 0 39312 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_369
timestamp 1698431365
transform 1 0 42672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_373
timestamp 1698431365
transform 1 0 43120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_6
timestamp 1698431365
transform 1 0 2016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_42
timestamp 1698431365
transform 1 0 6048 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_52
timestamp 1698431365
transform 1 0 7168 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_59
timestamp 1698431365
transform 1 0 7952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_77
timestamp 1698431365
transform 1 0 9968 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_81
timestamp 1698431365
transform 1 0 10416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_157
timestamp 1698431365
transform 1 0 18928 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_170
timestamp 1698431365
transform 1 0 20384 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_174
timestamp 1698431365
transform 1 0 20832 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_206
timestamp 1698431365
transform 1 0 24416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_222
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_227
timestamp 1698431365
transform 1 0 26768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_229
timestamp 1698431365
transform 1 0 26992 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_259
timestamp 1698431365
transform 1 0 30352 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_316
timestamp 1698431365
transform 1 0 36736 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_370
timestamp 1698431365
transform 1 0 42784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_372
timestamp 1698431365
transform 1 0 43008 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_428
timestamp 1698431365
transform 1 0 49280 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_31
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_50
timestamp 1698431365
transform 1 0 6944 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_59
timestamp 1698431365
transform 1 0 7952 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_74
timestamp 1698431365
transform 1 0 9632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_78
timestamp 1698431365
transform 1 0 10080 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_86
timestamp 1698431365
transform 1 0 10976 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_90
timestamp 1698431365
transform 1 0 11424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_98
timestamp 1698431365
transform 1 0 12320 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_102
timestamp 1698431365
transform 1 0 12768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_204
timestamp 1698431365
transform 1 0 24192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_208
timestamp 1698431365
transform 1 0 24640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_212
timestamp 1698431365
transform 1 0 25088 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_277
timestamp 1698431365
transform 1 0 32368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_281
timestamp 1698431365
transform 1 0 32816 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_367
timestamp 1698431365
transform 1 0 42448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_378
timestamp 1698431365
transform 1 0 43680 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_50
timestamp 1698431365
transform 1 0 6944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_77
timestamp 1698431365
transform 1 0 9968 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_93
timestamp 1698431365
transform 1 0 11760 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_101
timestamp 1698431365
transform 1 0 12656 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_105
timestamp 1698431365
transform 1 0 13104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_121
timestamp 1698431365
transform 1 0 14896 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_123
timestamp 1698431365
transform 1 0 15120 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_151
timestamp 1698431365
transform 1 0 18256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_186
timestamp 1698431365
transform 1 0 22176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_188
timestamp 1698431365
transform 1 0 22400 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_262
timestamp 1698431365
transform 1 0 30688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_268
timestamp 1698431365
transform 1 0 31360 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_272
timestamp 1698431365
transform 1 0 31808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_286
timestamp 1698431365
transform 1 0 33376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_288
timestamp 1698431365
transform 1 0 33600 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_297
timestamp 1698431365
transform 1 0 34608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_299
timestamp 1698431365
transform 1 0 34832 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_361
timestamp 1698431365
transform 1 0 41776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_363
timestamp 1698431365
transform 1 0 42000 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_401
timestamp 1698431365
transform 1 0 46256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_428
timestamp 1698431365
transform 1 0 49280 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_31
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_142
timestamp 1698431365
transform 1 0 17248 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_166
timestamp 1698431365
transform 1 0 19936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_168
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_184
timestamp 1698431365
transform 1 0 21952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_186
timestamp 1698431365
transform 1 0 22176 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_197
timestamp 1698431365
transform 1 0 23408 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698431365
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_249
timestamp 1698431365
transform 1 0 29232 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_258
timestamp 1698431365
transform 1 0 30240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_260
timestamp 1698431365
transform 1 0 30464 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_295
timestamp 1698431365
transform 1 0 34384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_297
timestamp 1698431365
transform 1 0 34608 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_359
timestamp 1698431365
transform 1 0 41552 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_361
timestamp 1698431365
transform 1 0 41776 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_10
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_15
timestamp 1698431365
transform 1 0 3024 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_31
timestamp 1698431365
transform 1 0 4816 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_77
timestamp 1698431365
transform 1 0 9968 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_118
timestamp 1698431365
transform 1 0 14560 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_126
timestamp 1698431365
transform 1 0 15456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_132
timestamp 1698431365
transform 1 0 16128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_171
timestamp 1698431365
transform 1 0 20496 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_237
timestamp 1698431365
transform 1 0 27888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_263
timestamp 1698431365
transform 1 0 30800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_275
timestamp 1698431365
transform 1 0 32144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_295
timestamp 1698431365
transform 1 0 34384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_299
timestamp 1698431365
transform 1 0 34832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_364
timestamp 1698431365
transform 1 0 42112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_417
timestamp 1698431365
transform 1 0 48048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_419
timestamp 1698431365
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_428
timestamp 1698431365
transform 1 0 49280 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_31
timestamp 1698431365
transform 1 0 4816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_87
timestamp 1698431365
transform 1 0 11088 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_91
timestamp 1698431365
transform 1 0 11536 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_99
timestamp 1698431365
transform 1 0 12432 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_103
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_170
timestamp 1698431365
transform 1 0 20384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_210
timestamp 1698431365
transform 1 0 24864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_241
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_257
timestamp 1698431365
transform 1 0 30128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_261
timestamp 1698431365
transform 1 0 30576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_265
timestamp 1698431365
transform 1 0 31024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_277
timestamp 1698431365
transform 1 0 32368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_281
timestamp 1698431365
transform 1 0 32816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_285
timestamp 1698431365
transform 1 0 33264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_295
timestamp 1698431365
transform 1 0 34384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_299
timestamp 1698431365
transform 1 0 34832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_307
timestamp 1698431365
transform 1 0 35728 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_327
timestamp 1698431365
transform 1 0 37968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_347
timestamp 1698431365
transform 1 0 40208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_371
timestamp 1698431365
transform 1 0 42896 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_396
timestamp 1698431365
transform 1 0 45696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_10
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_14
timestamp 1698431365
transform 1 0 2912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_16
timestamp 1698431365
transform 1 0 3136 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_88
timestamp 1698431365
transform 1 0 11200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_90
timestamp 1698431365
transform 1 0 11424 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698431365
transform 1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_154
timestamp 1698431365
transform 1 0 18592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_173
timestamp 1698431365
transform 1 0 20720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_252
timestamp 1698431365
transform 1 0 29568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_256
timestamp 1698431365
transform 1 0 30016 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_271
timestamp 1698431365
transform 1 0 31696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_275
timestamp 1698431365
transform 1 0 32144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_306
timestamp 1698431365
transform 1 0 35616 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_321
timestamp 1698431365
transform 1 0 37296 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_332
timestamp 1698431365
transform 1 0 38528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_336
timestamp 1698431365
transform 1 0 38976 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_340
timestamp 1698431365
transform 1 0 39424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_344
timestamp 1698431365
transform 1 0 39872 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_348
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_358
timestamp 1698431365
transform 1 0 41440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_426
timestamp 1698431365
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_428
timestamp 1698431365
transform 1 0 49280 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_45
timestamp 1698431365
transform 1 0 6384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_49
timestamp 1698431365
transform 1 0 6832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_63
timestamp 1698431365
transform 1 0 8400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_67
timestamp 1698431365
transform 1 0 8848 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_284
timestamp 1698431365
transform 1 0 33152 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_286
timestamp 1698431365
transform 1 0 33376 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_292
timestamp 1698431365
transform 1 0 34048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_306
timestamp 1698431365
transform 1 0 35616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_308
timestamp 1698431365
transform 1 0 35840 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_425
timestamp 1698431365
transform 1 0 48944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_31
timestamp 1698431365
transform 1 0 4816 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_50
timestamp 1698431365
transform 1 0 6944 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_54
timestamp 1698431365
transform 1 0 7392 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_61
timestamp 1698431365
transform 1 0 8176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_65
timestamp 1698431365
transform 1 0 8624 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_82
timestamp 1698431365
transform 1 0 10528 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_90
timestamp 1698431365
transform 1 0 11424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_116
timestamp 1698431365
transform 1 0 14336 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_196
timestamp 1698431365
transform 1 0 23296 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_200
timestamp 1698431365
transform 1 0 23744 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_203
timestamp 1698431365
transform 1 0 24080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698431365
transform 1 0 24528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_317
timestamp 1698431365
transform 1 0 36848 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_354
timestamp 1698431365
transform 1 0 40992 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_407
timestamp 1698431365
transform 1 0 46928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_411
timestamp 1698431365
transform 1 0 47376 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_426
timestamp 1698431365
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_428
timestamp 1698431365
transform 1 0 49280 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_18
timestamp 1698431365
transform 1 0 3360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_20
timestamp 1698431365
transform 1 0 3584 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_67
timestamp 1698431365
transform 1 0 8848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_71
timestamp 1698431365
transform 1 0 9296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_73
timestamp 1698431365
transform 1 0 9520 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_88
timestamp 1698431365
transform 1 0 11200 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_92
timestamp 1698431365
transform 1 0 11648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_94
timestamp 1698431365
transform 1 0 11872 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_127
timestamp 1698431365
transform 1 0 15568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_159
timestamp 1698431365
transform 1 0 19152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_161
timestamp 1698431365
transform 1 0 19376 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_181
timestamp 1698431365
transform 1 0 21616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_217
timestamp 1698431365
transform 1 0 25648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_221
timestamp 1698431365
transform 1 0 26096 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_229
timestamp 1698431365
transform 1 0 26992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_240
timestamp 1698431365
transform 1 0 28224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_276
timestamp 1698431365
transform 1 0 32256 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_278
timestamp 1698431365
transform 1 0 32480 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_389
timestamp 1698431365
transform 1 0 44912 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_428
timestamp 1698431365
transform 1 0 49280 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_37
timestamp 1698431365
transform 1 0 5488 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_126
timestamp 1698431365
transform 1 0 15456 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_155
timestamp 1698431365
transform 1 0 18704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_159
timestamp 1698431365
transform 1 0 19152 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_162
timestamp 1698431365
transform 1 0 19488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_166
timestamp 1698431365
transform 1 0 19936 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_174
timestamp 1698431365
transform 1 0 20832 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_253
timestamp 1698431365
transform 1 0 29680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_255
timestamp 1698431365
transform 1 0 29904 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_272
timestamp 1698431365
transform 1 0 31808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1698431365
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_426
timestamp 1698431365
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_428
timestamp 1698431365
transform 1 0 49280 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_6
timestamp 1698431365
transform 1 0 2016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_8
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_99
timestamp 1698431365
transform 1 0 12432 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_163
timestamp 1698431365
transform 1 0 19600 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_167
timestamp 1698431365
transform 1 0 20048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_206
timestamp 1698431365
transform 1 0 24416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_208
timestamp 1698431365
transform 1 0 24640 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_238
timestamp 1698431365
transform 1 0 28000 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_256
timestamp 1698431365
transform 1 0 30016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_260
timestamp 1698431365
transform 1 0 30464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_322
timestamp 1698431365
transform 1 0 37408 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_391
timestamp 1698431365
transform 1 0 45136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_395
timestamp 1698431365
transform 1 0 45584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_399
timestamp 1698431365
transform 1 0 46032 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_80
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_84
timestamp 1698431365
transform 1 0 10752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_106
timestamp 1698431365
transform 1 0 13216 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_108
timestamp 1698431365
transform 1 0 13440 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_168
timestamp 1698431365
transform 1 0 20160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_172
timestamp 1698431365
transform 1 0 20608 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_216
timestamp 1698431365
transform 1 0 25536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_260
timestamp 1698431365
transform 1 0 30464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_264
timestamp 1698431365
transform 1 0 30912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_268
timestamp 1698431365
transform 1 0 31360 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_272
timestamp 1698431365
transform 1 0 31808 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_314
timestamp 1698431365
transform 1 0 36512 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_316
timestamp 1698431365
transform 1 0 36736 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_410
timestamp 1698431365
transform 1 0 47264 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_415
timestamp 1698431365
transform 1 0 47824 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_426
timestamp 1698431365
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_428
timestamp 1698431365
transform 1 0 49280 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_10
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_14
timestamp 1698431365
transform 1 0 2912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_102
timestamp 1698431365
transform 1 0 12768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_111
timestamp 1698431365
transform 1 0 13776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_131
timestamp 1698431365
transform 1 0 16016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_143
timestamp 1698431365
transform 1 0 17360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_192
timestamp 1698431365
transform 1 0 22848 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_230
timestamp 1698431365
transform 1 0 27104 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_240
timestamp 1698431365
transform 1 0 28224 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_305
timestamp 1698431365
transform 1 0 35504 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_10
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_14
timestamp 1698431365
transform 1 0 2912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_40
timestamp 1698431365
transform 1 0 5824 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_48
timestamp 1698431365
transform 1 0 6720 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_80
timestamp 1698431365
transform 1 0 10304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_88
timestamp 1698431365
transform 1 0 11200 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_92
timestamp 1698431365
transform 1 0 11648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_94
timestamp 1698431365
transform 1 0 11872 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_103
timestamp 1698431365
transform 1 0 12880 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_204
timestamp 1698431365
transform 1 0 24192 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_278
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_317
timestamp 1698431365
transform 1 0 36848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_364
timestamp 1698431365
transform 1 0 42112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_426
timestamp 1698431365
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_428
timestamp 1698431365
transform 1 0 49280 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_31
timestamp 1698431365
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_63
timestamp 1698431365
transform 1 0 8400 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_67
timestamp 1698431365
transform 1 0 8848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_109
timestamp 1698431365
transform 1 0 13552 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_207
timestamp 1698431365
transform 1 0 24528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_209
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_218
timestamp 1698431365
transform 1 0 25760 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_251
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_255
timestamp 1698431365
transform 1 0 29904 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_257
timestamp 1698431365
transform 1 0 30128 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_260
timestamp 1698431365
transform 1 0 30464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_280
timestamp 1698431365
transform 1 0 32704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_346
timestamp 1698431365
transform 1 0 40096 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_426
timestamp 1698431365
transform 1 0 49056 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_428
timestamp 1698431365
transform 1 0 49280 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_6
timestamp 1698431365
transform 1 0 2016 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_21
timestamp 1698431365
transform 1 0 3696 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_33
timestamp 1698431365
transform 1 0 5040 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_67
timestamp 1698431365
transform 1 0 8848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_162
timestamp 1698431365
transform 1 0 19488 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_164
timestamp 1698431365
transform 1 0 19712 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_175
timestamp 1698431365
transform 1 0 20944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_214
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_221
timestamp 1698431365
transform 1 0 26096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_225
timestamp 1698431365
transform 1 0 26544 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_228
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_232
timestamp 1698431365
transform 1 0 27328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_236
timestamp 1698431365
transform 1 0 27776 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_240
timestamp 1698431365
transform 1 0 28224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_244
timestamp 1698431365
transform 1 0 28672 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_250
timestamp 1698431365
transform 1 0 29344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_258
timestamp 1698431365
transform 1 0 30240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_262
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_266
timestamp 1698431365
transform 1 0 31136 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_275
timestamp 1698431365
transform 1 0 32144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_277
timestamp 1698431365
transform 1 0 32368 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_409
timestamp 1698431365
transform 1 0 47152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_428
timestamp 1698431365
transform 1 0 49280 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_31
timestamp 1698431365
transform 1 0 4816 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_68
timestamp 1698431365
transform 1 0 8960 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_88
timestamp 1698431365
transform 1 0 11200 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_204
timestamp 1698431365
transform 1 0 24192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_235
timestamp 1698431365
transform 1 0 27664 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_240
timestamp 1698431365
transform 1 0 28224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_274
timestamp 1698431365
transform 1 0 32032 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_352
timestamp 1698431365
transform 1 0 40768 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_399
timestamp 1698431365
transform 1 0 46032 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_89
timestamp 1698431365
transform 1 0 11312 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_147
timestamp 1698431365
transform 1 0 17808 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_157
timestamp 1698431365
transform 1 0 18928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_172
timestamp 1698431365
transform 1 0 20608 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_208
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_222
timestamp 1698431365
transform 1 0 26208 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_238
timestamp 1698431365
transform 1 0 28000 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_256
timestamp 1698431365
transform 1 0 30016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_260
timestamp 1698431365
transform 1 0 30464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_264
timestamp 1698431365
transform 1 0 30912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_385
timestamp 1698431365
transform 1 0 44464 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_428
timestamp 1698431365
transform 1 0 49280 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_47
timestamp 1698431365
transform 1 0 6608 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_52
timestamp 1698431365
transform 1 0 7168 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_61
timestamp 1698431365
transform 1 0 8176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_65
timestamp 1698431365
transform 1 0 8624 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_103
timestamp 1698431365
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_113
timestamp 1698431365
transform 1 0 14000 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_145
timestamp 1698431365
transform 1 0 17584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_147
timestamp 1698431365
transform 1 0 17808 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_187
timestamp 1698431365
transform 1 0 22288 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_191
timestamp 1698431365
transform 1 0 22736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_193
timestamp 1698431365
transform 1 0 22960 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_243
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_264
timestamp 1698431365
transform 1 0 30912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_268
timestamp 1698431365
transform 1 0 31360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_276
timestamp 1698431365
transform 1 0 32256 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_282
timestamp 1698431365
transform 1 0 32928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_383
timestamp 1698431365
transform 1 0 44240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_398
timestamp 1698431365
transform 1 0 45920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_20
timestamp 1698431365
transform 1 0 3584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_22
timestamp 1698431365
transform 1 0 3808 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_33
timestamp 1698431365
transform 1 0 5040 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_49
timestamp 1698431365
transform 1 0 6832 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_60
timestamp 1698431365
transform 1 0 8064 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_68
timestamp 1698431365
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_98
timestamp 1698431365
transform 1 0 12320 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_120
timestamp 1698431365
transform 1 0 14784 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_128
timestamp 1698431365
transform 1 0 15680 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_137
timestamp 1698431365
transform 1 0 16688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_146
timestamp 1698431365
transform 1 0 17696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_148
timestamp 1698431365
transform 1 0 17920 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_151
timestamp 1698431365
transform 1 0 18256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_167
timestamp 1698431365
transform 1 0 20048 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_171
timestamp 1698431365
transform 1 0 20496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_246
timestamp 1698431365
transform 1 0 28896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_266
timestamp 1698431365
transform 1 0 31136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_288
timestamp 1698431365
transform 1 0 33600 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_290
timestamp 1698431365
transform 1 0 33824 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_293
timestamp 1698431365
transform 1 0 34160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_329
timestamp 1698431365
transform 1 0 38192 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_333
timestamp 1698431365
transform 1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_358
timestamp 1698431365
transform 1 0 41440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_360
timestamp 1698431365
transform 1 0 41664 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_374
timestamp 1698431365
transform 1 0 43232 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_376
timestamp 1698431365
transform 1 0 43456 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_389
timestamp 1698431365
transform 1 0 44912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_428
timestamp 1698431365
transform 1 0 49280 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_103
timestamp 1698431365
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_136
timestamp 1698431365
transform 1 0 16576 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_140
timestamp 1698431365
transform 1 0 17024 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_159
timestamp 1698431365
transform 1 0 19152 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_167
timestamp 1698431365
transform 1 0 20048 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_174
timestamp 1698431365
transform 1 0 20832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_252
timestamp 1698431365
transform 1 0 29568 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_261
timestamp 1698431365
transform 1 0 30576 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_269
timestamp 1698431365
transform 1 0 31472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_319
timestamp 1698431365
transform 1 0 37072 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_349
timestamp 1698431365
transform 1 0 40432 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_351
timestamp 1698431365
transform 1 0 40656 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_428
timestamp 1698431365
transform 1 0 49280 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_14
timestamp 1698431365
transform 1 0 2912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_122
timestamp 1698431365
transform 1 0 15008 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_135
timestamp 1698431365
transform 1 0 16464 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_173
timestamp 1698431365
transform 1 0 20720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_205
timestamp 1698431365
transform 1 0 24304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_220
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_224
timestamp 1698431365
transform 1 0 26432 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_260
timestamp 1698431365
transform 1 0 30464 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_268
timestamp 1698431365
transform 1 0 31360 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_358
timestamp 1698431365
transform 1 0 41440 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_428
timestamp 1698431365
transform 1 0 49280 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_41
timestamp 1698431365
transform 1 0 5936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_72
timestamp 1698431365
transform 1 0 9408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_74
timestamp 1698431365
transform 1 0 9632 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_96
timestamp 1698431365
transform 1 0 12096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_98
timestamp 1698431365
transform 1 0 12320 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_109
timestamp 1698431365
transform 1 0 13552 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_132
timestamp 1698431365
transform 1 0 16128 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_140
timestamp 1698431365
transform 1 0 17024 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_152
timestamp 1698431365
transform 1 0 18368 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_156
timestamp 1698431365
transform 1 0 18816 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_170
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_206
timestamp 1698431365
transform 1 0 24416 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_236
timestamp 1698431365
transform 1 0 27776 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_276
timestamp 1698431365
transform 1 0 32256 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_319
timestamp 1698431365
transform 1 0 37072 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_337
timestamp 1698431365
transform 1 0 39088 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_362
timestamp 1698431365
transform 1 0 41888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_366
timestamp 1698431365
transform 1 0 42336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_368
timestamp 1698431365
transform 1 0 42560 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_10
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_21
timestamp 1698431365
transform 1 0 3696 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_25
timestamp 1698431365
transform 1 0 4144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_27
timestamp 1698431365
transform 1 0 4368 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_34
timestamp 1698431365
transform 1 0 5152 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_38
timestamp 1698431365
transform 1 0 5600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_40
timestamp 1698431365
transform 1 0 5824 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_47
timestamp 1698431365
transform 1 0 6608 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_55
timestamp 1698431365
transform 1 0 7504 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_67
timestamp 1698431365
transform 1 0 8848 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_69
timestamp 1698431365
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698431365
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_150
timestamp 1698431365
transform 1 0 18144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_152
timestamp 1698431365
transform 1 0 18368 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_204
timestamp 1698431365
transform 1 0 24192 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_230
timestamp 1698431365
transform 1 0 27104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_238
timestamp 1698431365
transform 1 0 28000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_242
timestamp 1698431365
transform 1 0 28448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_244
timestamp 1698431365
transform 1 0 28672 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_253
timestamp 1698431365
transform 1 0 29680 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_263
timestamp 1698431365
transform 1 0 30800 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_356
timestamp 1698431365
transform 1 0 41216 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_360
timestamp 1698431365
transform 1 0 41664 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_410
timestamp 1698431365
transform 1 0 47264 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_418
timestamp 1698431365
transform 1 0 48160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_428
timestamp 1698431365
transform 1 0 49280 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_16
timestamp 1698431365
transform 1 0 3136 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_32
timestamp 1698431365
transform 1 0 4928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_43
timestamp 1698431365
transform 1 0 6160 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_75
timestamp 1698431365
transform 1 0 9744 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_79
timestamp 1698431365
transform 1 0 10192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_87
timestamp 1698431365
transform 1 0 11088 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_103
timestamp 1698431365
transform 1 0 12880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_116
timestamp 1698431365
transform 1 0 14336 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_118
timestamp 1698431365
transform 1 0 14560 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_137
timestamp 1698431365
transform 1 0 16688 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_179
timestamp 1698431365
transform 1 0 21392 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_228
timestamp 1698431365
transform 1 0 26880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698431365
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_236
timestamp 1698431365
transform 1 0 27776 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_239
timestamp 1698431365
transform 1 0 28112 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_258
timestamp 1698431365
transform 1 0 30240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_260
timestamp 1698431365
transform 1 0 30464 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698431365
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_321
timestamp 1698431365
transform 1 0 37296 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_380
timestamp 1698431365
transform 1 0 43904 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_31
timestamp 1698431365
transform 1 0 4816 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_46
timestamp 1698431365
transform 1 0 6496 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_58
timestamp 1698431365
transform 1 0 7840 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_60
timestamp 1698431365
transform 1 0 8064 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_80
timestamp 1698431365
transform 1 0 10304 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_96
timestamp 1698431365
transform 1 0 12096 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_139
timestamp 1698431365
transform 1 0 16912 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_158
timestamp 1698431365
transform 1 0 19040 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_166
timestamp 1698431365
transform 1 0 19936 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_168
timestamp 1698431365
transform 1 0 20160 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_216
timestamp 1698431365
transform 1 0 25536 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_220
timestamp 1698431365
transform 1 0 25984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_237
timestamp 1698431365
transform 1 0 27888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_278
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_286
timestamp 1698431365
transform 1 0 33376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_290
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_292
timestamp 1698431365
transform 1 0 34048 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_361
timestamp 1698431365
transform 1 0 41776 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_365
timestamp 1698431365
transform 1 0 42224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_369
timestamp 1698431365
transform 1 0 42672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_373
timestamp 1698431365
transform 1 0 43120 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_394
timestamp 1698431365
transform 1 0 45472 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_415
timestamp 1698431365
transform 1 0 47824 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_428
timestamp 1698431365
transform 1 0 49280 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_45
timestamp 1698431365
transform 1 0 6384 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_117
timestamp 1698431365
transform 1 0 14448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_119
timestamp 1698431365
transform 1 0 14672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_140
timestamp 1698431365
transform 1 0 17024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_148
timestamp 1698431365
transform 1 0 17920 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_152
timestamp 1698431365
transform 1 0 18368 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_186
timestamp 1698431365
transform 1 0 22176 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_297
timestamp 1698431365
transform 1 0 34608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_310
timestamp 1698431365
transform 1 0 36064 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_338
timestamp 1698431365
transform 1 0 39200 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_380
timestamp 1698431365
transform 1 0 43904 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_398
timestamp 1698431365
transform 1 0 45920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_420
timestamp 1698431365
transform 1 0 48384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_428
timestamp 1698431365
transform 1 0 49280 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_16
timestamp 1698431365
transform 1 0 3136 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_49
timestamp 1698431365
transform 1 0 6832 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_53
timestamp 1698431365
transform 1 0 7280 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_62
timestamp 1698431365
transform 1 0 8288 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_69
timestamp 1698431365
transform 1 0 9072 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_87
timestamp 1698431365
transform 1 0 11088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_89
timestamp 1698431365
transform 1 0 11312 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_160
timestamp 1698431365
transform 1 0 19264 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_187
timestamp 1698431365
transform 1 0 22288 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_204
timestamp 1698431365
transform 1 0 24192 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_223
timestamp 1698431365
transform 1 0 26320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_229
timestamp 1698431365
transform 1 0 26992 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_239
timestamp 1698431365
transform 1 0 28112 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_278
timestamp 1698431365
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_300
timestamp 1698431365
transform 1 0 34944 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_330
timestamp 1698431365
transform 1 0 38304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_332
timestamp 1698431365
transform 1 0 38528 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_356
timestamp 1698431365
transform 1 0 41216 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_428
timestamp 1698431365
transform 1 0 49280 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_31
timestamp 1698431365
transform 1 0 4816 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_67
timestamp 1698431365
transform 1 0 8848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_71
timestamp 1698431365
transform 1 0 9296 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_159
timestamp 1698431365
transform 1 0 19152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_206
timestamp 1698431365
transform 1 0 24416 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_237
timestamp 1698431365
transform 1 0 27888 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_321
timestamp 1698431365
transform 1 0 37296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_396
timestamp 1698431365
transform 1 0 45696 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_4
timestamp 1698431365
transform 1 0 1792 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_55
timestamp 1698431365
transform 1 0 7504 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_63
timestamp 1698431365
transform 1 0 8400 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_67
timestamp 1698431365
transform 1 0 8848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_69
timestamp 1698431365
transform 1 0 9072 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_74
timestamp 1698431365
transform 1 0 9632 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_104
timestamp 1698431365
transform 1 0 12992 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_106
timestamp 1698431365
transform 1 0 13216 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_113
timestamp 1698431365
transform 1 0 14000 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_121
timestamp 1698431365
transform 1 0 14896 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_125
timestamp 1698431365
transform 1 0 15344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_127
timestamp 1698431365
transform 1 0 15568 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_150
timestamp 1698431365
transform 1 0 18144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_162
timestamp 1698431365
transform 1 0 19488 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_164
timestamp 1698431365
transform 1 0 19712 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_169
timestamp 1698431365
transform 1 0 20272 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_185
timestamp 1698431365
transform 1 0 22064 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_192
timestamp 1698431365
transform 1 0 22848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_196
timestamp 1698431365
transform 1 0 23296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_200
timestamp 1698431365
transform 1 0 23744 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_292
timestamp 1698431365
transform 1 0 34048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_356
timestamp 1698431365
transform 1 0 41216 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_403
timestamp 1698431365
transform 1 0 46480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_415
timestamp 1698431365
transform 1 0 47824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698431365
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_31
timestamp 1698431365
transform 1 0 4816 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_100
timestamp 1698431365
transform 1 0 12544 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_115
timestamp 1698431365
transform 1 0 14224 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_125
timestamp 1698431365
transform 1 0 15344 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_133
timestamp 1698431365
transform 1 0 16240 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_142
timestamp 1698431365
transform 1 0 17248 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_154
timestamp 1698431365
transform 1 0 18592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_156
timestamp 1698431365
transform 1 0 18816 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_161
timestamp 1698431365
transform 1 0 19376 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_169
timestamp 1698431365
transform 1 0 20272 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_173
timestamp 1698431365
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_179
timestamp 1698431365
transform 1 0 21392 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_200
timestamp 1698431365
transform 1 0 23744 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_243
timestamp 1698431365
transform 1 0 28560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_251
timestamp 1698431365
transform 1 0 29456 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_253
timestamp 1698431365
transform 1 0 29680 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_263
timestamp 1698431365
transform 1 0 30800 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_286
timestamp 1698431365
transform 1 0 33376 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_310
timestamp 1698431365
transform 1 0 36064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_314
timestamp 1698431365
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_325
timestamp 1698431365
transform 1 0 37744 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_327
timestamp 1698431365
transform 1 0 37968 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_384
timestamp 1698431365
transform 1 0 44352 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_398
timestamp 1698431365
transform 1 0 45920 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_10
timestamp 1698431365
transform 1 0 2464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_12
timestamp 1698431365
transform 1 0 2688 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_92
timestamp 1698431365
transform 1 0 11648 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_108
timestamp 1698431365
transform 1 0 13440 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_110
timestamp 1698431365
transform 1 0 13664 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_148
timestamp 1698431365
transform 1 0 17920 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_208
timestamp 1698431365
transform 1 0 24640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_216
timestamp 1698431365
transform 1 0 25536 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_218
timestamp 1698431365
transform 1 0 25760 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_225
timestamp 1698431365
transform 1 0 26544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_227
timestamp 1698431365
transform 1 0 26768 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_259
timestamp 1698431365
transform 1 0 30352 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_265
timestamp 1698431365
transform 1 0 31024 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_278
timestamp 1698431365
transform 1 0 32480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_395
timestamp 1698431365
transform 1 0 45584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_415
timestamp 1698431365
transform 1 0 47824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_419
timestamp 1698431365
transform 1 0 48272 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_428
timestamp 1698431365
transform 1 0 49280 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_31
timestamp 1698431365
transform 1 0 4816 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_48
timestamp 1698431365
transform 1 0 6720 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_99
timestamp 1698431365
transform 1 0 12432 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_103
timestamp 1698431365
transform 1 0 12880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_123
timestamp 1698431365
transform 1 0 15120 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_131
timestamp 1698431365
transform 1 0 16016 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_162
timestamp 1698431365
transform 1 0 19488 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_166
timestamp 1698431365
transform 1 0 19936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_172
timestamp 1698431365
transform 1 0 20608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_196
timestamp 1698431365
transform 1 0 23296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_198
timestamp 1698431365
transform 1 0 23520 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_242
timestamp 1698431365
transform 1 0 28448 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_244
timestamp 1698431365
transform 1 0 28672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_280
timestamp 1698431365
transform 1 0 32704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_313
timestamp 1698431365
transform 1 0 36400 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_360
timestamp 1698431365
transform 1 0 41664 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_362
timestamp 1698431365
transform 1 0 41888 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_424
timestamp 1698431365
transform 1 0 48832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_428
timestamp 1698431365
transform 1 0 49280 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_6
timestamp 1698431365
transform 1 0 2016 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_36
timestamp 1698431365
transform 1 0 5376 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_40
timestamp 1698431365
transform 1 0 5824 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_78
timestamp 1698431365
transform 1 0 10080 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_110
timestamp 1698431365
transform 1 0 13664 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_126
timestamp 1698431365
transform 1 0 15456 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_134
timestamp 1698431365
transform 1 0 16352 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_138
timestamp 1698431365
transform 1 0 16800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_150
timestamp 1698431365
transform 1 0 18144 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_218
timestamp 1698431365
transform 1 0 25760 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_248
timestamp 1698431365
transform 1 0 29120 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_252
timestamp 1698431365
transform 1 0 29568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_293
timestamp 1698431365
transform 1 0 34160 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_315
timestamp 1698431365
transform 1 0 36624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_317
timestamp 1698431365
transform 1 0 36848 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698431365
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_354
timestamp 1698431365
transform 1 0 40992 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_428
timestamp 1698431365
transform 1 0 49280 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_18
timestamp 1698431365
transform 1 0 3360 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_44
timestamp 1698431365
transform 1 0 6272 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_46
timestamp 1698431365
transform 1 0 6496 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_84
timestamp 1698431365
transform 1 0 10752 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_100
timestamp 1698431365
transform 1 0 12544 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_107 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_209
timestamp 1698431365
transform 1 0 24752 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_217
timestamp 1698431365
transform 1 0 25648 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_221
timestamp 1698431365
transform 1 0 26096 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_244
timestamp 1698431365
transform 1 0 28672 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_255
timestamp 1698431365
transform 1 0 29904 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_352
timestamp 1698431365
transform 1 0 40768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_354
timestamp 1698431365
transform 1 0 40992 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_391
timestamp 1698431365
transform 1 0 45136 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_10
timestamp 1698431365
transform 1 0 2464 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_14
timestamp 1698431365
transform 1 0 2912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_16
timestamp 1698431365
transform 1 0 3136 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_65
timestamp 1698431365
transform 1 0 8624 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_69
timestamp 1698431365
transform 1 0 9072 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_136
timestamp 1698431365
transform 1 0 16576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_150
timestamp 1698431365
transform 1 0 18144 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_154
timestamp 1698431365
transform 1 0 18592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_184
timestamp 1698431365
transform 1 0 21952 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_200
timestamp 1698431365
transform 1 0 23744 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_208
timestamp 1698431365
transform 1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_241
timestamp 1698431365
transform 1 0 28336 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_243
timestamp 1698431365
transform 1 0 28560 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_279
timestamp 1698431365
transform 1 0 32592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_286
timestamp 1698431365
transform 1 0 33376 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_290
timestamp 1698431365
transform 1 0 33824 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_323
timestamp 1698431365
transform 1 0 37520 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_333
timestamp 1698431365
transform 1 0 38640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_337
timestamp 1698431365
transform 1 0 39088 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_341
timestamp 1698431365
transform 1 0 39536 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_345
timestamp 1698431365
transform 1 0 39984 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_347
timestamp 1698431365
transform 1 0 40208 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_381
timestamp 1698431365
transform 1 0 44016 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_417
timestamp 1698431365
transform 1 0 48048 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_419
timestamp 1698431365
transform 1 0 48272 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_428
timestamp 1698431365
transform 1 0 49280 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_36
timestamp 1698431365
transform 1 0 5376 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_44
timestamp 1698431365
transform 1 0 6272 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_51
timestamp 1698431365
transform 1 0 7056 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_67
timestamp 1698431365
transform 1 0 8848 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_70
timestamp 1698431365
transform 1 0 9184 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_104
timestamp 1698431365
transform 1 0 12992 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_138
timestamp 1698431365
transform 1 0 16800 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_154
timestamp 1698431365
transform 1 0 18592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_156
timestamp 1698431365
transform 1 0 18816 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_167
timestamp 1698431365
transform 1 0 20048 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_169
timestamp 1698431365
transform 1 0 20272 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_172
timestamp 1698431365
transform 1 0 20608 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_206
timestamp 1698431365
transform 1 0 24416 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_214
timestamp 1698431365
transform 1 0 25312 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_218
timestamp 1698431365
transform 1 0 25760 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_220
timestamp 1698431365
transform 1 0 25984 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_227
timestamp 1698431365
transform 1 0 26768 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_235
timestamp 1698431365
transform 1 0 27664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_237
timestamp 1698431365
transform 1 0 27888 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_240
timestamp 1698431365
transform 1 0 28224 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_248
timestamp 1698431365
transform 1 0 29120 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_255
timestamp 1698431365
transform 1 0 29904 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_259
timestamp 1698431365
transform 1 0 30352 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_261
timestamp 1698431365
transform 1 0 30576 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_303
timestamp 1698431365
transform 1 0 35280 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_305
timestamp 1698431365
transform 1 0 35504 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_314
timestamp 1698431365
transform 1 0 36512 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_318
timestamp 1698431365
transform 1 0 36960 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_320
timestamp 1698431365
transform 1 0 37184 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_323
timestamp 1698431365
transform 1 0 37520 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_327
timestamp 1698431365
transform 1 0 37968 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_331
timestamp 1698431365
transform 1 0 38416 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_335
timestamp 1698431365
transform 1 0 38864 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_339
timestamp 1698431365
transform 1 0 39312 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_342
timestamp 1698431365
transform 1 0 39648 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_344
timestamp 1698431365
transform 1 0 39872 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_347
timestamp 1698431365
transform 1 0 40208 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_351
timestamp 1698431365
transform 1 0 40656 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_373
timestamp 1698431365
transform 1 0 43120 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_382
timestamp 1698431365
transform 1 0 44128 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_405
timestamp 1698431365
transform 1 0 46704 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_407
timestamp 1698431365
transform 1 0 46928 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_410
timestamp 1698431365
transform 1 0 47264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_412
timestamp 1698431365
transform 1 0 47488 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 49392 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2
timestamp 1698431365
transform -1 0 49392 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform -1 0 48496 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input4
timestamp 1698431365
transform -1 0 49392 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input5
timestamp 1698431365
transform -1 0 49392 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input6
timestamp 1698431365
transform -1 0 48384 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input7
timestamp 1698431365
transform -1 0 49392 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input8
timestamp 1698431365
transform -1 0 44464 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input9
timestamp 1698431365
transform -1 0 48384 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1698431365
transform -1 0 49392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform -1 0 48384 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input12
timestamp 1698431365
transform -1 0 31808 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input13
timestamp 1698431365
transform -1 0 45136 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input14
timestamp 1698431365
transform 1 0 19152 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698431365
transform -1 0 31808 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform 1 0 38304 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform 1 0 37408 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform 1 0 41328 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform 1 0 17360 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_57 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 49616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 49616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 49616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 49616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 49616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 49616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 49616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 49616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 49616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 49616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 49616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 49616 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 49616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 49616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 49616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 49616 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 49616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 49616 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 49616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 49616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 49616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 49616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 49616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 49616 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 49616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 49616 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 49616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 49616 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 49616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 49616 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 49616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 49616 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 49616 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 49616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 49616 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 49616 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 49616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 49616 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 49616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 49616 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 49616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 49616 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 49616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 49616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 49616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 49616 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 49616 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 49616 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 49616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 49616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 49616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 49616 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 49616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_110
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 49616 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_111
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 49616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_112
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 49616 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_113
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 49616 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_118
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_119
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_120
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_121
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_122
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_123
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_124
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_125
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_126
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_127
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_128
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_129
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_130
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_131
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_132
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_133
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_134
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_135
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_136
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_137
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_138
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_139
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_140
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_141
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_142
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_143
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_144
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_145
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_146
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_147
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_148
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_149
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_150
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_151
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_152
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_153
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_154
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_155
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_156
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_157
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_158
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_159
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_160
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_161
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_162
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_163
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_164
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_165
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_166
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_167
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_168
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_169
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_170
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_171
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_172
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_173
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_174
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_175
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_176
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_177
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_178
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_179
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_180
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_181
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_182
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_183
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_184
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_185
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_186
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_187
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_188
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_189
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_190
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_191
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_192
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_193
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_194
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_195
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_196
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_197
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_198
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_199
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_200
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_201
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_202
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_203
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_204
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_205
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_206
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_207
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_208
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_209
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_210
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_211
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_212
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_213
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_214
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_215
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_216
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_217
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_218
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_219
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_220
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_221
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_222
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_223
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_224
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_225
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_226
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_227
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_228
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_229
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_230
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_231
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_232
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_233
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_234
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_235
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_236
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_237
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_238
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_239
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_240
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_241
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_242
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_243
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_244
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_245
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_246
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_247
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_248
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_249
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_250
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_251
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_252
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_253
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_254
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_255
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_256
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_257
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_258
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_259
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_260
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_261
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_262
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_263
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_264
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_265
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_266
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_267
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_268
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_269
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_270
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_271
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_272
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_273
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_274
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_275
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_276
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_277
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_278
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_279
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_280
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_281
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_282
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_283
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_284
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_285
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_286
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_287
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_288
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_289
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_290
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_291
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_292
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_293
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_294
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_295
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_296
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_297
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_298
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_299
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_300
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_301
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_302
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_303
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_304
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_305
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_306
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_307
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_308
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_309
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_310
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_311
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_312
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_313
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_314
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_315
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_316
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_317
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_318
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_319
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_320
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_321
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_322
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_323
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_324
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_325
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_326
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_327
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_328
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_329
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_330
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_331
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_332
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_333
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_334
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_335
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_336
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_337
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_338
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_339
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_340
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_341
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_342
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_343
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_344
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_345
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_346
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_347
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_348
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_349
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_350
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_351
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_352
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_353
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_354
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_355
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_356
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_357
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_358
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_359
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_360
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_361
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_362
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_363
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_364
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_365
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_366
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_367
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_368
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_369
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_370
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_371
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_372
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_373
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_374
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_375
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_376
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_377
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_378
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_379
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_380
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_381
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_382
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_383
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_384
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_385
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_386
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_387
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_388
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_389
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_390
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_391
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_392
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_393
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_394
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_395
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_396
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_397
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_398
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_399
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_400
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_401
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_402
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_403
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_404
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_405
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_406
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_407
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_408
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_409
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_410
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_411
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_412
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_413
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_414
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_415
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_416
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_417
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_418
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_419
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_420
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_421
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_422
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_423
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_424
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_425
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_426
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_427
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_428
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_429
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_430
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_431
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_432
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_433
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_434
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_435
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_436
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_437
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_438
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_439
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_440
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_441
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_442
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_443
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_444
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_445
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_446
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_447
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_448
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_449
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_450
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_451
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_452
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_453
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_454
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_455
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_456
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_457
timestamp 1698431365
transform 1 0 8960 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_458
timestamp 1698431365
transform 1 0 12768 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_459
timestamp 1698431365
transform 1 0 16576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_460
timestamp 1698431365
transform 1 0 20384 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_461
timestamp 1698431365
transform 1 0 24192 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_462
timestamp 1698431365
transform 1 0 28000 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_463
timestamp 1698431365
transform 1 0 31808 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_464
timestamp 1698431365
transform 1 0 35616 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_465
timestamp 1698431365
transform 1 0 39424 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_466
timestamp 1698431365
transform 1 0 43232 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_467
timestamp 1698431365
transform 1 0 47040 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_24 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_25
timestamp 1698431365
transform -1 0 3472 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_26
timestamp 1698431365
transform -1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_27
timestamp 1698431365
transform -1 0 7056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_28
timestamp 1698431365
transform 1 0 7168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_29
timestamp 1698431365
transform 1 0 7616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_30
timestamp 1698431365
transform 1 0 8064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_31
timestamp 1698431365
transform 1 0 8512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_32
timestamp 1698431365
transform -1 0 25088 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_33
timestamp 1698431365
transform -1 0 28672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_34
timestamp 1698431365
transform -1 0 28448 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_35
timestamp 1698431365
transform -1 0 31920 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_36
timestamp 1698431365
transform -1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_37
timestamp 1698431365
transform -1 0 48384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_38
timestamp 1698431365
transform -1 0 48384 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_39
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_40
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_41
timestamp 1698431365
transform 1 0 47040 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_42
timestamp 1698431365
transform -1 0 45136 0 1 4704
box -86 -86 534 870
<< labels >>
flabel metal3 s 50200 36064 51000 36176 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 50200 40320 51000 40432 0 FreeSans 448 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal3 s 50200 44576 51000 44688 0 FreeSans 448 0 0 0 custom_settings[2]
port 2 nsew signal input
flabel metal3 s 50200 48832 51000 48944 0 FreeSans 448 0 0 0 custom_settings[3]
port 3 nsew signal input
flabel metal3 s 50200 2016 51000 2128 0 FreeSans 448 0 0 0 io_in_1[0]
port 4 nsew signal input
flabel metal3 s 50200 6272 51000 6384 0 FreeSans 448 0 0 0 io_in_1[1]
port 5 nsew signal input
flabel metal3 s 50200 10528 51000 10640 0 FreeSans 448 0 0 0 io_in_1[2]
port 6 nsew signal input
flabel metal3 s 50200 14784 51000 14896 0 FreeSans 448 0 0 0 io_in_1[3]
port 7 nsew signal input
flabel metal3 s 50200 19040 51000 19152 0 FreeSans 448 0 0 0 io_in_1[4]
port 8 nsew signal input
flabel metal3 s 50200 23296 51000 23408 0 FreeSans 448 0 0 0 io_in_1[5]
port 9 nsew signal input
flabel metal3 s 50200 27552 51000 27664 0 FreeSans 448 0 0 0 io_in_1[6]
port 10 nsew signal input
flabel metal3 s 50200 31808 51000 31920 0 FreeSans 448 0 0 0 io_in_1[7]
port 11 nsew signal input
flabel metal2 s 31808 50200 31920 51000 0 FreeSans 448 90 0 0 io_in_2[0]
port 12 nsew signal input
flabel metal2 s 44576 50200 44688 51000 0 FreeSans 448 90 0 0 io_in_2[1]
port 13 nsew signal input
flabel metal2 s 1120 0 1232 800 0 FreeSans 448 90 0 0 io_out[0]
port 14 nsew signal tristate
flabel metal2 s 19040 0 19152 800 0 FreeSans 448 90 0 0 io_out[10]
port 15 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 io_out[11]
port 16 nsew signal tristate
flabel metal2 s 22624 0 22736 800 0 FreeSans 448 90 0 0 io_out[12]
port 17 nsew signal tristate
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 io_out[13]
port 18 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 io_out[14]
port 19 nsew signal tristate
flabel metal2 s 28000 0 28112 800 0 FreeSans 448 90 0 0 io_out[15]
port 20 nsew signal tristate
flabel metal2 s 29792 0 29904 800 0 FreeSans 448 90 0 0 io_out[16]
port 21 nsew signal tristate
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 io_out[17]
port 22 nsew signal tristate
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 io_out[18]
port 23 nsew signal tristate
flabel metal2 s 35168 0 35280 800 0 FreeSans 448 90 0 0 io_out[19]
port 24 nsew signal tristate
flabel metal2 s 2912 0 3024 800 0 FreeSans 448 90 0 0 io_out[1]
port 25 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 io_out[20]
port 26 nsew signal tristate
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 io_out[21]
port 27 nsew signal tristate
flabel metal2 s 40544 0 40656 800 0 FreeSans 448 90 0 0 io_out[22]
port 28 nsew signal tristate
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 io_out[23]
port 29 nsew signal tristate
flabel metal2 s 44128 0 44240 800 0 FreeSans 448 90 0 0 io_out[24]
port 30 nsew signal tristate
flabel metal2 s 45920 0 46032 800 0 FreeSans 448 90 0 0 io_out[25]
port 31 nsew signal tristate
flabel metal2 s 47712 0 47824 800 0 FreeSans 448 90 0 0 io_out[26]
port 32 nsew signal tristate
flabel metal2 s 49504 0 49616 800 0 FreeSans 448 90 0 0 io_out[27]
port 33 nsew signal tristate
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 io_out[2]
port 34 nsew signal tristate
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 io_out[3]
port 35 nsew signal tristate
flabel metal2 s 8288 0 8400 800 0 FreeSans 448 90 0 0 io_out[4]
port 36 nsew signal tristate
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 io_out[5]
port 37 nsew signal tristate
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 io_out[6]
port 38 nsew signal tristate
flabel metal2 s 13664 0 13776 800 0 FreeSans 448 90 0 0 io_out[7]
port 39 nsew signal tristate
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 io_out[8]
port 40 nsew signal tristate
flabel metal2 s 17248 0 17360 800 0 FreeSans 448 90 0 0 io_out[9]
port 41 nsew signal tristate
flabel metal2 s 19040 50200 19152 51000 0 FreeSans 448 90 0 0 rst_n
port 42 nsew signal input
flabel metal4 s 4448 3076 4768 47884 0 FreeSans 1280 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 35168 3076 35488 47884 0 FreeSans 1280 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 19808 3076 20128 47884 0 FreeSans 1280 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal2 s 6272 50200 6384 51000 0 FreeSans 448 90 0 0 wb_clk_i
port 45 nsew signal input
rlabel metal1 25480 47824 25480 47824 0 vdd
rlabel metal1 25480 47040 25480 47040 0 vss
rlabel metal2 8232 45864 8232 45864 0 _0000_
rlabel metal2 5544 47376 5544 47376 0 _0001_
rlabel metal2 3080 45472 3080 45472 0 _0002_
rlabel metal2 2520 43932 2520 43932 0 _0003_
rlabel metal2 9576 45360 9576 45360 0 _0004_
rlabel metal2 7896 42224 7896 42224 0 _0005_
rlabel metal2 10696 41216 10696 41216 0 _0006_
rlabel metal2 2520 43064 2520 43064 0 _0007_
rlabel metal2 2632 40656 2632 40656 0 _0008_
rlabel metal2 2968 39424 2968 39424 0 _0009_
rlabel metal2 2576 38248 2576 38248 0 _0010_
rlabel metal2 8904 38976 8904 38976 0 _0011_
rlabel metal2 10136 39200 10136 39200 0 _0012_
rlabel metal2 8456 36624 8456 36624 0 _0013_
rlabel metal2 11816 37576 11816 37576 0 _0014_
rlabel metal2 10584 34720 10584 34720 0 _0015_
rlabel metal3 10024 33208 10024 33208 0 _0016_
rlabel metal2 6664 32480 6664 32480 0 _0017_
rlabel metal2 10136 30968 10136 30968 0 _0018_
rlabel metal2 8232 28280 8232 28280 0 _0019_
rlabel metal2 4312 23296 4312 23296 0 _0020_
rlabel metal2 2744 22008 2744 22008 0 _0021_
rlabel metal3 4368 24584 4368 24584 0 _0022_
rlabel metal2 6832 26152 6832 26152 0 _0023_
rlabel metal2 2520 26656 2520 26656 0 _0024_
rlabel metal2 2520 27496 2520 27496 0 _0025_
rlabel metal2 2520 30352 2520 30352 0 _0026_
rlabel metal2 2520 31892 2520 31892 0 _0027_
rlabel metal2 2576 35896 2576 35896 0 _0028_
rlabel metal2 3192 32984 3192 32984 0 _0029_
rlabel metal2 4144 35560 4144 35560 0 _0030_
rlabel metal2 6440 34552 6440 34552 0 _0031_
rlabel metal2 33096 31976 33096 31976 0 _0032_
rlabel metal3 34328 30184 34328 30184 0 _0033_
rlabel metal2 33320 32984 33320 32984 0 _0034_
rlabel metal2 40936 32984 40936 32984 0 _0035_
rlabel metal3 37800 30072 37800 30072 0 _0036_
rlabel metal2 19544 21896 19544 21896 0 _0037_
rlabel metal2 19432 21952 19432 21952 0 _0038_
rlabel metal2 22624 19880 22624 19880 0 _0039_
rlabel metal2 22792 21560 22792 21560 0 _0040_
rlabel metal3 29736 4200 29736 4200 0 _0041_
rlabel metal2 28616 6216 28616 6216 0 _0042_
rlabel metal2 25368 3696 25368 3696 0 _0043_
rlabel metal2 25032 5320 25032 5320 0 _0044_
rlabel metal2 24136 8512 24136 8512 0 _0045_
rlabel metal2 20776 7000 20776 7000 0 _0046_
rlabel metal3 24360 4200 24360 4200 0 _0047_
rlabel metal2 17864 6328 17864 6328 0 _0048_
rlabel metal2 23016 4816 23016 4816 0 _0049_
rlabel metal2 37464 5264 37464 5264 0 _0050_
rlabel metal2 39480 7224 39480 7224 0 _0051_
rlabel metal2 47544 4312 47544 4312 0 _0052_
rlabel metal2 33936 7336 33936 7336 0 _0053_
rlabel metal2 44744 4760 44744 4760 0 _0054_
rlabel metal2 32200 3472 32200 3472 0 _0055_
rlabel metal2 44464 13832 44464 13832 0 _0056_
rlabel metal2 47096 8568 47096 8568 0 _0057_
rlabel metal2 47096 7280 47096 7280 0 _0058_
rlabel metal2 48888 7896 48888 7896 0 _0059_
rlabel metal2 25704 10192 25704 10192 0 _0060_
rlabel metal2 24472 11760 24472 11760 0 _0061_
rlabel metal2 21672 13384 21672 13384 0 _0062_
rlabel metal2 18536 13272 18536 13272 0 _0063_
rlabel metal2 14112 15176 14112 15176 0 _0064_
rlabel metal2 15904 11928 15904 11928 0 _0065_
rlabel metal2 13832 10920 13832 10920 0 _0066_
rlabel metal3 16856 8344 16856 8344 0 _0067_
rlabel metal2 24696 37688 24696 37688 0 _0068_
rlabel metal2 26824 36792 26824 36792 0 _0069_
rlabel metal2 27832 39928 27832 39928 0 _0070_
rlabel metal2 24584 39928 24584 39928 0 _0071_
rlabel metal2 23464 41496 23464 41496 0 _0072_
rlabel metal3 23408 43624 23408 43624 0 _0073_
rlabel metal2 20440 45528 20440 45528 0 _0074_
rlabel metal2 19992 43176 19992 43176 0 _0075_
rlabel metal2 26488 23380 26488 23380 0 _0076_
rlabel metal2 26488 22008 26488 22008 0 _0077_
rlabel metal2 29344 24024 29344 24024 0 _0078_
rlabel metal3 30632 23800 30632 23800 0 _0079_
rlabel metal2 37128 37576 37128 37576 0 _0080_
rlabel metal3 32088 37464 32088 37464 0 _0081_
rlabel metal3 33544 38584 33544 38584 0 _0082_
rlabel metal2 36456 40096 36456 40096 0 _0083_
rlabel metal2 30016 43736 30016 43736 0 _0084_
rlabel metal2 29960 39312 29960 39312 0 _0085_
rlabel metal2 24696 42392 24696 42392 0 _0086_
rlabel metal2 25592 41720 25592 41720 0 _0087_
rlabel metal2 35112 4648 35112 4648 0 _0088_
rlabel metal2 36624 9128 36624 9128 0 _0089_
rlabel metal2 32536 9408 32536 9408 0 _0090_
rlabel metal3 33600 5096 33600 5096 0 _0091_
rlabel metal2 32088 7000 32088 7000 0 _0092_
rlabel metal2 21784 10192 21784 10192 0 _0093_
rlabel metal2 18424 11312 18424 11312 0 _0094_
rlabel metal2 18200 9296 18200 9296 0 _0095_
rlabel metal2 9464 10136 9464 10136 0 _0096_
rlabel metal2 9576 7560 9576 7560 0 _0097_
rlabel metal2 13608 6720 13608 6720 0 _0098_
rlabel metal2 16072 7616 16072 7616 0 _0099_
rlabel metal2 15288 7896 15288 7896 0 _0100_
rlabel metal2 5992 9352 5992 9352 0 _0101_
rlabel metal2 5320 7784 5320 7784 0 _0102_
rlabel metal2 6216 6440 6216 6440 0 _0103_
rlabel metal3 7168 4200 7168 4200 0 _0104_
rlabel metal2 9912 3976 9912 3976 0 _0105_
rlabel metal2 11816 4312 11816 4312 0 _0106_
rlabel metal2 16072 4536 16072 4536 0 _0107_
rlabel metal2 17304 4200 17304 4200 0 _0108_
rlabel metal2 24472 13496 24472 13496 0 _0109_
rlabel metal2 27888 14616 27888 14616 0 _0110_
rlabel metal2 41048 37688 41048 37688 0 _0111_
rlabel metal2 39816 38360 39816 38360 0 _0112_
rlabel metal2 40376 39256 40376 39256 0 _0113_
rlabel metal2 39984 40600 39984 40600 0 _0114_
rlabel metal3 37800 44408 37800 44408 0 _0115_
rlabel metal2 38080 45192 38080 45192 0 _0116_
rlabel metal2 38472 46200 38472 46200 0 _0117_
rlabel metal3 39480 41888 39480 41888 0 _0118_
rlabel metal2 27048 27776 27048 27776 0 _0119_
rlabel metal3 29960 28616 29960 28616 0 _0120_
rlabel metal3 24584 27720 24584 27720 0 _0121_
rlabel metal2 26824 25928 26824 25928 0 _0122_
rlabel metal2 23464 23744 23464 23744 0 _0123_
rlabel metal2 23128 25928 23128 25928 0 _0124_
rlabel metal2 19992 24304 19992 24304 0 _0125_
rlabel metal3 22456 26936 22456 26936 0 _0126_
rlabel metal2 32928 3640 32928 3640 0 _0127_
rlabel metal2 39144 5656 39144 5656 0 _0128_
rlabel metal2 36792 3864 36792 3864 0 _0129_
rlabel metal3 12096 11256 12096 11256 0 _0130_
rlabel metal2 24696 16632 24696 16632 0 _0131_
rlabel metal2 30744 17976 30744 17976 0 _0132_
rlabel metal3 28056 16968 28056 16968 0 _0133_
rlabel metal3 25032 17640 25032 17640 0 _0134_
rlabel metal2 30016 14616 30016 14616 0 _0135_
rlabel metal3 33600 18424 33600 18424 0 _0136_
rlabel metal2 42056 21168 42056 21168 0 _0137_
rlabel metal2 45080 13328 45080 13328 0 _0138_
rlabel metal3 46648 12712 46648 12712 0 _0139_
rlabel metal3 47992 9912 47992 9912 0 _0140_
rlabel metal2 45640 11536 45640 11536 0 _0141_
rlabel metal2 47880 17136 47880 17136 0 _0142_
rlabel metal2 47096 20944 47096 20944 0 _0143_
rlabel metal2 39536 35000 39536 35000 0 _0144_
rlabel metal3 41944 33432 41944 33432 0 _0145_
rlabel metal2 41664 35000 41664 35000 0 _0146_
rlabel metal2 42168 33208 42168 33208 0 _0147_
rlabel metal2 48888 34440 48888 34440 0 _0148_
rlabel metal3 46480 33432 46480 33432 0 _0149_
rlabel metal3 48160 40264 48160 40264 0 _0150_
rlabel metal2 48552 39704 48552 39704 0 _0151_
rlabel metal3 44240 38696 44240 38696 0 _0152_
rlabel metal3 47544 39368 47544 39368 0 _0153_
rlabel metal2 47096 41720 47096 41720 0 _0154_
rlabel metal2 47096 42896 47096 42896 0 _0155_
rlabel metal2 48104 45136 48104 45136 0 _0156_
rlabel metal2 45080 47040 45080 47040 0 _0157_
rlabel metal2 41720 46984 41720 46984 0 _0158_
rlabel metal2 42616 43120 42616 43120 0 _0159_
rlabel metal2 45528 16968 45528 16968 0 _0160_
rlabel metal2 14616 15288 14616 15288 0 _0161_
rlabel metal2 11704 16520 11704 16520 0 _0162_
rlabel metal2 10808 14168 10808 14168 0 _0163_
rlabel metal2 8120 16240 8120 16240 0 _0164_
rlabel metal2 8680 18032 8680 18032 0 _0165_
rlabel metal2 7560 20216 7560 20216 0 _0166_
rlabel metal2 6216 21000 6216 21000 0 _0167_
rlabel metal2 5992 19432 5992 19432 0 _0168_
rlabel metal2 3080 20440 3080 20440 0 _0169_
rlabel metal3 3192 18312 3192 18312 0 _0170_
rlabel metal2 2352 16744 2352 16744 0 _0171_
rlabel metal2 3416 15736 3416 15736 0 _0172_
rlabel metal2 2520 14112 2520 14112 0 _0173_
rlabel metal2 5992 12880 5992 12880 0 _0174_
rlabel metal2 2520 11760 2520 11760 0 _0175_
rlabel metal2 7392 10472 7392 10472 0 _0176_
rlabel metal2 9800 13104 9800 13104 0 _0177_
rlabel metal2 35672 12096 35672 12096 0 _0178_
rlabel metal2 32200 27888 32200 27888 0 _0179_
rlabel metal2 35168 26152 35168 26152 0 _0180_
rlabel metal2 33880 24360 33880 24360 0 _0181_
rlabel metal2 39256 25032 39256 25032 0 _0182_
rlabel metal2 38024 25872 38024 25872 0 _0183_
rlabel metal2 47096 19768 47096 19768 0 _0184_
rlabel metal2 22568 32200 22568 32200 0 _0185_
rlabel metal2 21672 34776 21672 34776 0 _0186_
rlabel metal2 18648 34944 18648 34944 0 _0187_
rlabel metal2 14840 43008 14840 43008 0 _0188_
rlabel metal2 17416 43960 17416 43960 0 _0189_
rlabel metal2 14056 41272 14056 41272 0 _0190_
rlabel metal2 13272 39144 13272 39144 0 _0191_
rlabel metal2 13720 36680 13720 36680 0 _0192_
rlabel metal3 13664 35000 13664 35000 0 _0193_
rlabel metal2 13160 32872 13160 32872 0 _0194_
rlabel metal2 14168 30464 14168 30464 0 _0195_
rlabel metal2 18424 28672 18424 28672 0 _0196_
rlabel metal2 28056 18928 28056 18928 0 _0197_
rlabel metal3 32200 35000 32200 35000 0 _0198_
rlabel metal2 32536 36120 32536 36120 0 _0199_
rlabel metal2 37464 42000 37464 42000 0 _0200_
rlabel metal2 35224 46984 35224 46984 0 _0201_
rlabel metal2 32424 47096 32424 47096 0 _0202_
rlabel metal2 29624 46984 29624 46984 0 _0203_
rlabel metal3 24920 44408 24920 44408 0 _0204_
rlabel metal2 26040 46984 26040 46984 0 _0205_
rlabel metal3 30408 36568 30408 36568 0 _0206_
rlabel metal2 25816 33376 25816 33376 0 _0207_
rlabel metal2 25592 31416 25592 31416 0 _0208_
rlabel metal2 28168 28952 28168 28952 0 _0209_
rlabel metal2 32872 20944 32872 20944 0 _0210_
rlabel metal2 22568 29848 22568 29848 0 _0211_
rlabel metal2 21392 29512 21392 29512 0 _0212_
rlabel metal2 15512 28896 15512 28896 0 _0213_
rlabel metal2 10472 29120 10472 29120 0 _0214_
rlabel metal2 12488 30464 12488 30464 0 _0215_
rlabel metal2 10136 25760 10136 25760 0 _0216_
rlabel metal2 13384 24024 13384 24024 0 _0217_
rlabel metal2 9968 24024 9968 24024 0 _0218_
rlabel metal2 10808 21280 10808 21280 0 _0219_
rlabel metal2 14168 17192 14168 17192 0 _0220_
rlabel metal2 11816 18760 11816 18760 0 _0221_
rlabel metal2 14952 20608 14952 20608 0 _0222_
rlabel metal3 25256 20888 25256 20888 0 _0223_
rlabel metal2 40040 15568 40040 15568 0 _0224_
rlabel metal2 39480 13160 39480 13160 0 _0225_
rlabel metal2 42840 12320 42840 12320 0 _0226_
rlabel metal2 45136 9128 45136 9128 0 _0227_
rlabel metal2 40040 6664 40040 6664 0 _0228_
rlabel metal2 38248 10248 38248 10248 0 _0229_
rlabel metal2 44744 11200 44744 11200 0 _0230_
rlabel metal2 37352 12880 37352 12880 0 _0231_
rlabel metal3 36232 14616 36232 14616 0 _0232_
rlabel metal3 39144 15848 39144 15848 0 _0233_
rlabel metal2 34328 19768 34328 19768 0 _0234_
rlabel metal2 39480 21168 39480 21168 0 _0235_
rlabel metal2 6888 24024 6888 24024 0 _0236_
rlabel metal2 19992 16464 19992 16464 0 _0237_
rlabel metal2 20328 17192 20328 17192 0 _0238_
rlabel metal3 22792 17752 22792 17752 0 _0239_
rlabel metal2 21448 19600 21448 19600 0 _0240_
rlabel metal2 44408 28392 44408 28392 0 _0241_
rlabel metal2 40040 28168 40040 28168 0 _0242_
rlabel metal2 43232 22232 43232 22232 0 _0243_
rlabel metal3 45304 24584 45304 24584 0 _0244_
rlabel metal2 45640 24080 45640 24080 0 _0245_
rlabel metal2 47096 23464 47096 23464 0 _0246_
rlabel metal3 47320 26936 47320 26936 0 _0247_
rlabel metal2 46984 25648 46984 25648 0 _0248_
rlabel metal3 30184 11480 30184 11480 0 _0249_
rlabel metal3 30352 10808 30352 10808 0 _0250_
rlabel metal2 33432 13720 33432 13720 0 _0251_
rlabel metal3 32368 13608 32368 13608 0 _0252_
rlabel metal2 44968 18088 44968 18088 0 _0253_
rlabel metal2 44408 20328 44408 20328 0 _0254_
rlabel metal2 42168 17472 42168 17472 0 _0255_
rlabel metal2 40488 17752 40488 17752 0 _0256_
rlabel metal2 39704 41776 39704 41776 0 _0257_
rlabel metal3 39900 44408 39900 44408 0 _0258_
rlabel metal2 40376 42224 40376 42224 0 _0259_
rlabel metal2 43288 20496 43288 20496 0 _0260_
rlabel metal2 25480 25872 25480 25872 0 _0261_
rlabel metal2 29176 26208 29176 26208 0 _0262_
rlabel metal2 24808 25592 24808 25592 0 _0263_
rlabel metal2 26600 28224 26600 28224 0 _0264_
rlabel metal2 26768 28056 26768 28056 0 _0265_
rlabel metal2 25816 16016 25816 16016 0 _0266_
rlabel metal2 29512 27832 29512 27832 0 _0267_
rlabel metal2 41720 22960 41720 22960 0 _0268_
rlabel metal2 25368 28280 25368 28280 0 _0269_
rlabel metal2 24864 17080 24864 17080 0 _0270_
rlabel metal3 27216 25368 27216 25368 0 _0271_
rlabel metal3 21392 25480 21392 25480 0 _0272_
rlabel metal3 21392 25256 21392 25256 0 _0273_
rlabel metal3 22064 24920 22064 24920 0 _0274_
rlabel metal3 23408 25368 23408 25368 0 _0275_
rlabel metal3 20048 25480 20048 25480 0 _0276_
rlabel metal2 22120 25872 22120 25872 0 _0277_
rlabel metal2 22008 11088 22008 11088 0 _0278_
rlabel metal3 41664 5992 41664 5992 0 _0279_
rlabel metal2 36456 5488 36456 5488 0 _0280_
rlabel metal2 12992 11368 12992 11368 0 _0281_
rlabel metal2 33880 18704 33880 18704 0 _0282_
rlabel metal2 29736 18592 29736 18592 0 _0283_
rlabel metal2 32312 17752 32312 17752 0 _0284_
rlabel metal2 29400 18760 29400 18760 0 _0285_
rlabel metal2 25816 18704 25816 18704 0 _0286_
rlabel metal2 31472 18648 31472 18648 0 _0287_
rlabel metal2 28560 17528 28560 17528 0 _0288_
rlabel metal2 27720 18088 27720 18088 0 _0289_
rlabel metal2 30968 17024 30968 17024 0 _0290_
rlabel metal3 33544 17752 33544 17752 0 _0291_
rlabel metal2 40936 19208 40936 19208 0 _0292_
rlabel metal2 45864 21336 45864 21336 0 _0293_
rlabel metal3 49336 10696 49336 10696 0 _0294_
rlabel metal2 47320 15596 47320 15596 0 _0295_
rlabel metal2 49000 20160 49000 20160 0 _0296_
rlabel metal2 48776 17024 48776 17024 0 _0297_
rlabel metal2 46760 19264 46760 19264 0 _0298_
rlabel metal2 44072 19544 44072 19544 0 _0299_
rlabel metal3 44744 16520 44744 16520 0 _0300_
rlabel metal2 45416 13104 45416 13104 0 _0301_
rlabel metal4 45864 15848 45864 15848 0 _0302_
rlabel metal2 48328 12992 48328 12992 0 _0303_
rlabel metal2 48160 11480 48160 11480 0 _0304_
rlabel metal2 47544 12208 47544 12208 0 _0305_
rlabel metal2 48776 11144 48776 11144 0 _0306_
rlabel metal2 49112 11648 49112 11648 0 _0307_
rlabel metal2 46704 12264 46704 12264 0 _0308_
rlabel metal2 48160 16296 48160 16296 0 _0309_
rlabel metal2 48776 15792 48776 15792 0 _0310_
rlabel metal2 48216 19320 48216 19320 0 _0311_
rlabel metal2 48552 29904 48552 29904 0 _0312_
rlabel metal2 48776 29960 48776 29960 0 _0313_
rlabel metal2 47880 29680 47880 29680 0 _0314_
rlabel metal2 44184 35672 44184 35672 0 _0315_
rlabel metal3 46928 30408 46928 30408 0 _0316_
rlabel metal2 44856 29512 44856 29512 0 _0317_
rlabel metal2 45304 30464 45304 30464 0 _0318_
rlabel metal2 45080 30408 45080 30408 0 _0319_
rlabel metal2 43624 31024 43624 31024 0 _0320_
rlabel metal2 42168 30184 42168 30184 0 _0321_
rlabel metal2 42728 30184 42728 30184 0 _0322_
rlabel metal2 41216 30968 41216 30968 0 _0323_
rlabel metal2 44352 31752 44352 31752 0 _0324_
rlabel metal2 42392 30520 42392 30520 0 _0325_
rlabel metal2 42784 29624 42784 29624 0 _0326_
rlabel metal2 45752 31808 45752 31808 0 _0327_
rlabel metal2 46984 29120 46984 29120 0 _0328_
rlabel metal3 45864 31864 45864 31864 0 _0329_
rlabel metal2 47432 29232 47432 29232 0 _0330_
rlabel metal2 47152 28728 47152 28728 0 _0331_
rlabel metal3 45472 36456 45472 36456 0 _0332_
rlabel metal2 48048 35448 48048 35448 0 _0333_
rlabel metal3 48048 32536 48048 32536 0 _0334_
rlabel metal3 46704 30968 46704 30968 0 _0335_
rlabel metal3 43400 44296 43400 44296 0 _0336_
rlabel metal3 44688 44184 44688 44184 0 _0337_
rlabel metal2 44800 42952 44800 42952 0 _0338_
rlabel metal3 45640 38808 45640 38808 0 _0339_
rlabel metal3 44912 38584 44912 38584 0 _0340_
rlabel metal2 45304 39424 45304 39424 0 _0341_
rlabel metal3 48888 39592 48888 39592 0 _0342_
rlabel metal2 43176 39816 43176 39816 0 _0343_
rlabel metal3 44464 39592 44464 39592 0 _0344_
rlabel metal2 47992 39816 47992 39816 0 _0345_
rlabel metal2 43400 40152 43400 40152 0 _0346_
rlabel metal2 43960 46536 43960 46536 0 _0347_
rlabel metal2 42728 45416 42728 45416 0 _0348_
rlabel metal3 44184 45640 44184 45640 0 _0349_
rlabel metal2 43624 42000 43624 42000 0 _0350_
rlabel metal2 42392 40768 42392 40768 0 _0351_
rlabel metal2 42840 43400 42840 43400 0 _0352_
rlabel metal2 44968 41216 44968 41216 0 _0353_
rlabel metal2 42616 44296 42616 44296 0 _0354_
rlabel metal2 43120 41944 43120 41944 0 _0355_
rlabel metal3 47040 44296 47040 44296 0 _0356_
rlabel metal2 44240 43288 44240 43288 0 _0357_
rlabel metal2 45416 43120 45416 43120 0 _0358_
rlabel metal2 44072 41496 44072 41496 0 _0359_
rlabel metal2 45528 41664 45528 41664 0 _0360_
rlabel metal2 45640 43232 45640 43232 0 _0361_
rlabel metal2 45304 38752 45304 38752 0 _0362_
rlabel metal3 45360 41720 45360 41720 0 _0363_
rlabel metal2 42616 40376 42616 40376 0 _0364_
rlabel metal3 43232 38136 43232 38136 0 _0365_
rlabel metal2 43512 30688 43512 30688 0 _0366_
rlabel metal2 46536 31360 46536 31360 0 _0367_
rlabel metal2 42560 41720 42560 41720 0 _0368_
rlabel metal2 42728 42336 42728 42336 0 _0369_
rlabel metal2 44968 42504 44968 42504 0 _0370_
rlabel metal2 43120 40264 43120 40264 0 _0371_
rlabel metal2 45864 30072 45864 30072 0 _0372_
rlabel metal3 45752 28840 45752 28840 0 _0373_
rlabel metal3 45976 30016 45976 30016 0 _0374_
rlabel metal2 46032 30184 46032 30184 0 _0375_
rlabel metal2 43960 30128 43960 30128 0 _0376_
rlabel metal2 44408 29288 44408 29288 0 _0377_
rlabel metal2 44072 12880 44072 12880 0 _0378_
rlabel metal3 42728 21560 42728 21560 0 _0379_
rlabel metal2 42616 16072 42616 16072 0 _0380_
rlabel metal2 42168 24640 42168 24640 0 _0381_
rlabel metal2 45528 28672 45528 28672 0 _0382_
rlabel metal2 46984 22400 46984 22400 0 _0383_
rlabel metal3 47320 21784 47320 21784 0 _0384_
rlabel metal3 45640 34104 45640 34104 0 _0385_
rlabel metal3 41216 47656 41216 47656 0 _0386_
rlabel metal2 26488 34440 26488 34440 0 _0387_
rlabel metal2 25816 32144 25816 32144 0 _0388_
rlabel metal3 31808 29400 31808 29400 0 _0389_
rlabel metal3 34048 26264 34048 26264 0 _0390_
rlabel metal3 26264 30240 26264 30240 0 _0391_
rlabel metal2 37576 36120 37576 36120 0 _0392_
rlabel metal3 41720 36288 41720 36288 0 _0393_
rlabel metal3 42560 34328 42560 34328 0 _0394_
rlabel metal2 24584 36064 24584 36064 0 _0395_
rlabel metal2 41048 29680 41048 29680 0 _0396_
rlabel metal2 39256 33544 39256 33544 0 _0397_
rlabel metal2 40264 32200 40264 32200 0 _0398_
rlabel metal2 40712 32312 40712 32312 0 _0399_
rlabel metal2 40936 35840 40936 35840 0 _0400_
rlabel metal3 43848 33208 43848 33208 0 _0401_
rlabel metal3 44128 32536 44128 32536 0 _0402_
rlabel metal3 43400 34104 43400 34104 0 _0403_
rlabel metal2 49000 42112 49000 42112 0 _0404_
rlabel metal2 48104 32368 48104 32368 0 _0405_
rlabel metal2 47208 34776 47208 34776 0 _0406_
rlabel metal3 45864 33880 45864 33880 0 _0407_
rlabel metal3 48104 34328 48104 34328 0 _0408_
rlabel metal2 47656 41944 47656 41944 0 _0409_
rlabel metal2 45528 34048 45528 34048 0 _0410_
rlabel metal2 45920 36456 45920 36456 0 _0411_
rlabel metal2 46872 37296 46872 37296 0 _0412_
rlabel metal3 47712 38920 47712 38920 0 _0413_
rlabel metal3 47768 40152 47768 40152 0 _0414_
rlabel metal3 46088 35000 46088 35000 0 _0415_
rlabel metal2 49056 39032 49056 39032 0 _0416_
rlabel metal2 45752 37744 45752 37744 0 _0417_
rlabel metal2 46032 38248 46032 38248 0 _0418_
rlabel metal3 47320 39480 47320 39480 0 _0419_
rlabel metal2 47600 38920 47600 38920 0 _0420_
rlabel metal2 47768 40152 47768 40152 0 _0421_
rlabel metal2 46088 44576 46088 44576 0 _0422_
rlabel metal2 47320 44016 47320 44016 0 _0423_
rlabel metal2 45416 45976 45416 45976 0 _0424_
rlabel metal3 43792 47208 43792 47208 0 _0425_
rlabel metal2 48440 44912 48440 44912 0 _0426_
rlabel metal2 48160 44072 48160 44072 0 _0427_
rlabel metal2 45640 46536 45640 46536 0 _0428_
rlabel metal2 44296 46144 44296 46144 0 _0429_
rlabel metal2 44184 46704 44184 46704 0 _0430_
rlabel metal2 41272 46760 41272 46760 0 _0431_
rlabel metal3 42168 42728 42168 42728 0 _0432_
rlabel metal2 45976 18816 45976 18816 0 _0433_
rlabel metal2 47488 20104 47488 20104 0 _0434_
rlabel metal2 46984 18144 46984 18144 0 _0435_
rlabel metal2 45528 18312 45528 18312 0 _0436_
rlabel metal2 45528 14784 45528 14784 0 _0437_
rlabel metal3 12096 12936 12096 12936 0 _0438_
rlabel metal3 10976 13832 10976 13832 0 _0439_
rlabel metal2 11144 16744 11144 16744 0 _0440_
rlabel metal2 13720 16016 13720 16016 0 _0441_
rlabel metal2 7672 13552 7672 13552 0 _0442_
rlabel metal2 6328 18032 6328 18032 0 _0443_
rlabel metal2 12208 17528 12208 17528 0 _0444_
rlabel metal2 13272 16072 13272 16072 0 _0445_
rlabel metal2 6552 15232 6552 15232 0 _0446_
rlabel metal3 22008 15792 22008 15792 0 _0447_
rlabel metal2 11816 15960 11816 15960 0 _0448_
rlabel metal2 11592 16744 11592 16744 0 _0449_
rlabel metal3 9464 13720 9464 13720 0 _0450_
rlabel metal2 10584 14000 10584 14000 0 _0451_
rlabel metal2 7336 15624 7336 15624 0 _0452_
rlabel metal2 7784 18480 7784 18480 0 _0453_
rlabel metal3 9240 16856 9240 16856 0 _0454_
rlabel metal2 8120 17136 8120 17136 0 _0455_
rlabel metal2 8344 19264 8344 19264 0 _0456_
rlabel metal2 8568 18592 8568 18592 0 _0457_
rlabel metal2 6720 18648 6720 18648 0 _0458_
rlabel metal2 9240 18424 9240 18424 0 _0459_
rlabel metal2 8568 20384 8568 20384 0 _0460_
rlabel metal2 9016 19600 9016 19600 0 _0461_
rlabel metal3 6776 19208 6776 19208 0 _0462_
rlabel metal2 6552 21056 6552 21056 0 _0463_
rlabel metal2 2968 14784 2968 14784 0 _0464_
rlabel metal2 5320 18984 5320 18984 0 _0465_
rlabel metal2 6328 19096 6328 19096 0 _0466_
rlabel metal2 3976 18256 3976 18256 0 _0467_
rlabel metal3 3864 18200 3864 18200 0 _0468_
rlabel metal2 5992 17080 5992 17080 0 _0469_
rlabel metal2 2800 20104 2800 20104 0 _0470_
rlabel metal3 3024 18424 3024 18424 0 _0471_
rlabel metal2 3304 18480 3304 18480 0 _0472_
rlabel metal2 2632 15232 2632 15232 0 _0473_
rlabel metal2 2072 16240 2072 16240 0 _0474_
rlabel metal2 3192 13888 3192 13888 0 _0475_
rlabel metal2 6888 14616 6888 14616 0 _0476_
rlabel metal3 5040 15288 5040 15288 0 _0477_
rlabel metal2 3864 15232 3864 15232 0 _0478_
rlabel metal2 4536 13888 4536 13888 0 _0479_
rlabel metal2 6776 11704 6776 11704 0 _0480_
rlabel metal2 4144 13832 4144 13832 0 _0481_
rlabel metal2 5880 13328 5880 13328 0 _0482_
rlabel metal2 6216 12992 6216 12992 0 _0483_
rlabel metal3 4928 10808 4928 10808 0 _0484_
rlabel metal2 3752 12208 3752 12208 0 _0485_
rlabel metal2 7448 11704 7448 11704 0 _0486_
rlabel metal2 6888 10640 6888 10640 0 _0487_
rlabel metal3 9464 20216 9464 20216 0 _0488_
rlabel metal2 6216 14224 6216 14224 0 _0489_
rlabel metal2 6104 12992 6104 12992 0 _0490_
rlabel metal3 7420 16072 7420 16072 0 _0491_
rlabel metal2 10304 15960 10304 15960 0 _0492_
rlabel metal2 9016 15624 9016 15624 0 _0493_
rlabel metal2 8680 15120 8680 15120 0 _0494_
rlabel metal2 8624 13720 8624 13720 0 _0495_
rlabel metal2 9688 12544 9688 12544 0 _0496_
rlabel metal3 36736 24024 36736 24024 0 _0497_
rlabel metal2 33936 27944 33936 27944 0 _0498_
rlabel metal2 35784 29064 35784 29064 0 _0499_
rlabel metal2 34104 28280 34104 28280 0 _0500_
rlabel metal2 35672 28112 35672 28112 0 _0501_
rlabel metal2 37352 27832 37352 27832 0 _0502_
rlabel metal2 38696 28896 38696 28896 0 _0503_
rlabel metal2 39144 28168 39144 28168 0 _0504_
rlabel metal2 38248 24528 38248 24528 0 _0505_
rlabel metal2 38808 28112 38808 28112 0 _0506_
rlabel metal2 38528 24136 38528 24136 0 _0507_
rlabel metal2 22568 12880 22568 12880 0 _0508_
rlabel metal2 35168 12824 35168 12824 0 _0509_
rlabel metal3 33488 27832 33488 27832 0 _0510_
rlabel metal3 39816 25424 39816 25424 0 _0511_
rlabel metal2 36680 25144 36680 25144 0 _0512_
rlabel metal2 26152 21280 26152 21280 0 _0513_
rlabel metal3 34552 25592 34552 25592 0 _0514_
rlabel metal2 37576 24640 37576 24640 0 _0515_
rlabel metal2 35448 23744 35448 23744 0 _0516_
rlabel metal2 39592 25760 39592 25760 0 _0517_
rlabel metal2 37352 23352 37352 23352 0 _0518_
rlabel metal2 22680 36848 22680 36848 0 _0519_
rlabel metal2 26264 19320 26264 19320 0 _0520_
rlabel metal2 22568 31696 22568 31696 0 _0521_
rlabel metal3 17864 33320 17864 33320 0 _0522_
rlabel metal3 19320 31528 19320 31528 0 _0523_
rlabel metal2 20216 32648 20216 32648 0 _0524_
rlabel metal2 17528 32256 17528 32256 0 _0525_
rlabel metal2 19712 32760 19712 32760 0 _0526_
rlabel metal2 19320 33712 19320 33712 0 _0527_
rlabel metal3 17136 32760 17136 32760 0 _0528_
rlabel metal3 19208 32536 19208 32536 0 _0529_
rlabel metal2 18760 31864 18760 31864 0 _0530_
rlabel metal2 19208 31304 19208 31304 0 _0531_
rlabel metal2 17416 33152 17416 33152 0 _0532_
rlabel metal2 18648 32536 18648 32536 0 _0533_
rlabel metal3 19824 32760 19824 32760 0 _0534_
rlabel metal2 20104 36736 20104 36736 0 _0535_
rlabel metal3 20216 39480 20216 39480 0 _0536_
rlabel metal2 18200 40264 18200 40264 0 _0537_
rlabel metal2 21672 39984 21672 39984 0 _0538_
rlabel metal2 21280 40600 21280 40600 0 _0539_
rlabel metal3 23464 35896 23464 35896 0 _0540_
rlabel metal3 22232 38136 22232 38136 0 _0541_
rlabel metal2 20552 40992 20552 40992 0 _0542_
rlabel via2 17080 41048 17080 41048 0 _0543_
rlabel metal2 19544 41440 19544 41440 0 _0544_
rlabel metal2 20048 39592 20048 39592 0 _0545_
rlabel metal3 21168 40376 21168 40376 0 _0546_
rlabel metal2 19768 40600 19768 40600 0 _0547_
rlabel metal3 20272 40264 20272 40264 0 _0548_
rlabel metal2 20776 39088 20776 39088 0 _0549_
rlabel metal3 20440 38584 20440 38584 0 _0550_
rlabel metal2 18200 39928 18200 39928 0 _0551_
rlabel via2 17752 38024 17752 38024 0 _0552_
rlabel metal3 16464 38024 16464 38024 0 _0553_
rlabel metal2 17976 37912 17976 37912 0 _0554_
rlabel metal2 18200 38080 18200 38080 0 _0555_
rlabel metal2 18312 37576 18312 37576 0 _0556_
rlabel metal2 18928 37912 18928 37912 0 _0557_
rlabel metal2 22400 38696 22400 38696 0 _0558_
rlabel metal2 19544 37128 19544 37128 0 _0559_
rlabel metal3 21336 37912 21336 37912 0 _0560_
rlabel metal2 19376 39592 19376 39592 0 _0561_
rlabel metal2 21784 38528 21784 38528 0 _0562_
rlabel metal2 22120 38864 22120 38864 0 _0563_
rlabel metal2 20216 39704 20216 39704 0 _0564_
rlabel metal3 19320 37464 19320 37464 0 _0565_
rlabel metal2 19320 37464 19320 37464 0 _0566_
rlabel metal2 19096 36960 19096 36960 0 _0567_
rlabel metal2 19768 36904 19768 36904 0 _0568_
rlabel metal2 19264 32760 19264 32760 0 _0569_
rlabel metal2 19432 32872 19432 32872 0 _0570_
rlabel metal2 20776 35336 20776 35336 0 _0571_
rlabel metal2 19712 26488 19712 26488 0 _0572_
rlabel metal2 21224 32256 21224 32256 0 _0573_
rlabel metal2 17416 41048 17416 41048 0 _0574_
rlabel metal2 20888 33096 20888 33096 0 _0575_
rlabel metal3 22624 35224 22624 35224 0 _0576_
rlabel metal3 22120 35672 22120 35672 0 _0577_
rlabel metal2 23576 35728 23576 35728 0 _0578_
rlabel metal2 18312 35728 18312 35728 0 _0579_
rlabel metal2 18872 35056 18872 35056 0 _0580_
rlabel metal3 17472 41160 17472 41160 0 _0581_
rlabel metal2 16856 42392 16856 42392 0 _0582_
rlabel metal3 15848 42616 15848 42616 0 _0583_
rlabel metal2 17640 40768 17640 40768 0 _0584_
rlabel metal2 17752 41496 17752 41496 0 _0585_
rlabel metal2 17976 42840 17976 42840 0 _0586_
rlabel metal2 14392 35392 14392 35392 0 _0587_
rlabel metal2 15344 39368 15344 39368 0 _0588_
rlabel via2 16184 39480 16184 39480 0 _0589_
rlabel metal3 14560 39592 14560 39592 0 _0590_
rlabel metal2 13608 39816 13608 39816 0 _0591_
rlabel metal3 14840 38696 14840 38696 0 _0592_
rlabel metal3 13160 38248 13160 38248 0 _0593_
rlabel metal2 16184 34832 16184 34832 0 _0594_
rlabel metal2 16184 37576 16184 37576 0 _0595_
rlabel metal2 14952 36904 14952 36904 0 _0596_
rlabel metal2 15568 36456 15568 36456 0 _0597_
rlabel metal2 14168 36120 14168 36120 0 _0598_
rlabel metal2 12712 36400 12712 36400 0 _0599_
rlabel metal2 17080 33544 17080 33544 0 _0600_
rlabel metal2 16296 33376 16296 33376 0 _0601_
rlabel metal2 17640 32928 17640 32928 0 _0602_
rlabel metal3 14784 33208 14784 33208 0 _0603_
rlabel metal3 16968 32536 16968 32536 0 _0604_
rlabel metal3 18200 30744 18200 30744 0 _0605_
rlabel metal2 16072 31640 16072 31640 0 _0606_
rlabel metal2 18424 21112 18424 21112 0 _0607_
rlabel metal3 29064 20552 29064 20552 0 _0608_
rlabel metal2 29512 20832 29512 20832 0 _0609_
rlabel metal2 35504 35000 35504 35000 0 _0610_
rlabel metal2 31528 35056 31528 35056 0 _0611_
rlabel via2 29848 34328 29848 34328 0 _0612_
rlabel metal3 29344 30744 29344 30744 0 _0613_
rlabel metal2 30184 32592 30184 32592 0 _0614_
rlabel metal2 27832 31640 27832 31640 0 _0615_
rlabel metal2 29960 32984 29960 32984 0 _0616_
rlabel metal2 29624 34272 29624 34272 0 _0617_
rlabel metal2 29400 34384 29400 34384 0 _0618_
rlabel metal2 29512 33768 29512 33768 0 _0619_
rlabel metal3 29344 32648 29344 32648 0 _0620_
rlabel metal3 28896 32312 28896 32312 0 _0621_
rlabel metal2 27888 34776 27888 34776 0 _0622_
rlabel metal2 29008 34776 29008 34776 0 _0623_
rlabel metal3 29792 34888 29792 34888 0 _0624_
rlabel metal2 30856 40712 30856 40712 0 _0625_
rlabel via2 35448 43624 35448 43624 0 _0626_
rlabel metal2 35112 44576 35112 44576 0 _0627_
rlabel metal2 35336 42784 35336 42784 0 _0628_
rlabel metal2 33096 42224 33096 42224 0 _0629_
rlabel metal2 36232 40600 36232 40600 0 _0630_
rlabel metal2 33320 41160 33320 41160 0 _0631_
rlabel metal2 31192 41440 31192 41440 0 _0632_
rlabel metal2 33768 44688 33768 44688 0 _0633_
rlabel metal2 32088 43400 32088 43400 0 _0634_
rlabel metal3 32144 42168 32144 42168 0 _0635_
rlabel metal2 33656 43652 33656 43652 0 _0636_
rlabel metal2 33208 43848 33208 43848 0 _0637_
rlabel metal2 32704 41944 32704 41944 0 _0638_
rlabel metal3 32984 41832 32984 41832 0 _0639_
rlabel metal2 33992 41496 33992 41496 0 _0640_
rlabel metal2 28392 43008 28392 43008 0 _0641_
rlabel metal2 28504 43120 28504 43120 0 _0642_
rlabel metal3 28112 44072 28112 44072 0 _0643_
rlabel metal2 28280 42952 28280 42952 0 _0644_
rlabel metal2 28560 41272 28560 41272 0 _0645_
rlabel metal2 29512 42224 29512 42224 0 _0646_
rlabel metal2 29848 40712 29848 40712 0 _0647_
rlabel metal2 38808 39872 38808 39872 0 _0648_
rlabel metal2 36232 38752 36232 38752 0 _0649_
rlabel metal2 31864 40656 31864 40656 0 _0650_
rlabel metal3 32648 42952 32648 42952 0 _0651_
rlabel metal3 35280 41384 35280 41384 0 _0652_
rlabel metal2 33712 40600 33712 40600 0 _0653_
rlabel metal2 33544 40432 33544 40432 0 _0654_
rlabel metal2 32760 43176 32760 43176 0 _0655_
rlabel metal2 28672 41048 28672 41048 0 _0656_
rlabel metal2 31528 42392 31528 42392 0 _0657_
rlabel metal2 31528 41496 31528 41496 0 _0658_
rlabel metal2 29904 35448 29904 35448 0 _0659_
rlabel metal2 30464 33544 30464 33544 0 _0660_
rlabel metal3 30576 37352 30576 37352 0 _0661_
rlabel metal2 30688 41384 30688 41384 0 _0662_
rlabel metal2 31864 33712 31864 33712 0 _0663_
rlabel metal2 30856 44744 30856 44744 0 _0664_
rlabel metal2 32088 33376 32088 33376 0 _0665_
rlabel metal2 37016 45080 37016 45080 0 _0666_
rlabel metal2 32760 37240 32760 37240 0 _0667_
rlabel metal2 32312 36400 32312 36400 0 _0668_
rlabel metal2 37240 43176 37240 43176 0 _0669_
rlabel metal3 36736 42952 36736 42952 0 _0670_
rlabel metal2 35224 45080 35224 45080 0 _0671_
rlabel metal2 36120 45136 36120 45136 0 _0672_
rlabel metal2 36400 45304 36400 45304 0 _0673_
rlabel metal3 33320 44968 33320 44968 0 _0674_
rlabel metal2 31528 45528 31528 45528 0 _0675_
rlabel metal2 30296 46144 30296 46144 0 _0676_
rlabel metal2 27608 43988 27608 43988 0 _0677_
rlabel metal2 30296 45192 30296 45192 0 _0678_
rlabel metal3 31472 45192 31472 45192 0 _0679_
rlabel metal2 30072 45584 30072 45584 0 _0680_
rlabel metal2 29736 46704 29736 46704 0 _0681_
rlabel metal2 27384 44744 27384 44744 0 _0682_
rlabel metal2 27048 44800 27048 44800 0 _0683_
rlabel metal2 26488 45472 26488 45472 0 _0684_
rlabel metal3 27384 45752 27384 45752 0 _0685_
rlabel metal3 26992 45864 26992 45864 0 _0686_
rlabel metal2 27048 46704 27048 46704 0 _0687_
rlabel metal2 27944 35896 27944 35896 0 _0688_
rlabel metal2 28616 36736 28616 36736 0 _0689_
rlabel metal2 27496 35168 27496 35168 0 _0690_
rlabel metal2 27384 33992 27384 33992 0 _0691_
rlabel metal2 27272 33712 27272 33712 0 _0692_
rlabel metal2 25592 32648 25592 32648 0 _0693_
rlabel metal2 27272 32760 27272 32760 0 _0694_
rlabel metal2 28336 33544 28336 33544 0 _0695_
rlabel metal2 25928 31696 25928 31696 0 _0696_
rlabel metal2 33320 22176 33320 22176 0 _0697_
rlabel metal2 31976 21728 31976 21728 0 _0698_
rlabel metal3 20160 28616 20160 28616 0 _0699_
rlabel metal2 22568 28560 22568 28560 0 _0700_
rlabel metal3 15624 18648 15624 18648 0 _0701_
rlabel metal2 17416 20720 17416 20720 0 _0702_
rlabel metal2 18760 20468 18760 20468 0 _0703_
rlabel via2 16296 19096 16296 19096 0 _0704_
rlabel metal3 17304 18424 17304 18424 0 _0705_
rlabel metal2 18200 19096 18200 19096 0 _0706_
rlabel metal2 16744 15568 16744 15568 0 _0707_
rlabel metal2 18704 18536 18704 18536 0 _0708_
rlabel metal3 17976 18200 17976 18200 0 _0709_
rlabel metal2 16744 17360 16744 17360 0 _0710_
rlabel metal2 15288 17920 15288 17920 0 _0711_
rlabel metal2 18536 18256 18536 18256 0 _0712_
rlabel metal2 18648 18256 18648 18256 0 _0713_
rlabel metal3 18480 23912 18480 23912 0 _0714_
rlabel metal2 15960 27552 15960 27552 0 _0715_
rlabel metal2 16632 28168 16632 28168 0 _0716_
rlabel metal2 16296 28336 16296 28336 0 _0717_
rlabel metal2 17192 27776 17192 27776 0 _0718_
rlabel metal2 21448 29848 21448 29848 0 _0719_
rlabel metal2 18312 27160 18312 27160 0 _0720_
rlabel metal3 17080 26264 17080 26264 0 _0721_
rlabel metal2 14280 26320 14280 26320 0 _0722_
rlabel metal3 15344 25704 15344 25704 0 _0723_
rlabel metal2 17696 26488 17696 26488 0 _0724_
rlabel metal2 15400 26264 15400 26264 0 _0725_
rlabel metal2 15008 25704 15008 25704 0 _0726_
rlabel metal2 16464 26936 16464 26936 0 _0727_
rlabel metal2 17584 27272 17584 27272 0 _0728_
rlabel metal2 18648 25536 18648 25536 0 _0729_
rlabel metal2 15624 25088 15624 25088 0 _0730_
rlabel metal3 15008 24584 15008 24584 0 _0731_
rlabel metal2 13160 23968 13160 23968 0 _0732_
rlabel metal2 16184 25144 16184 25144 0 _0733_
rlabel metal2 16296 24864 16296 24864 0 _0734_
rlabel metal2 16072 23968 16072 23968 0 _0735_
rlabel metal2 16968 24808 16968 24808 0 _0736_
rlabel metal2 19320 27272 19320 27272 0 _0737_
rlabel metal2 18760 26040 18760 26040 0 _0738_
rlabel metal2 18200 25032 18200 25032 0 _0739_
rlabel metal2 18256 26264 18256 26264 0 _0740_
rlabel metal2 18536 26992 18536 26992 0 _0741_
rlabel metal2 16856 27160 16856 27160 0 _0742_
rlabel metal2 17416 26600 17416 26600 0 _0743_
rlabel metal3 17248 25480 17248 25480 0 _0744_
rlabel metal2 16520 23744 16520 23744 0 _0745_
rlabel metal2 16744 24416 16744 24416 0 _0746_
rlabel metal2 20776 24416 20776 24416 0 _0747_
rlabel metal2 17864 17304 17864 17304 0 _0748_
rlabel metal2 18984 20468 18984 20468 0 _0749_
rlabel metal2 21112 23408 21112 23408 0 _0750_
rlabel metal3 25704 20552 25704 20552 0 _0751_
rlabel metal2 21448 27496 21448 27496 0 _0752_
rlabel via2 21112 28504 21112 28504 0 _0753_
rlabel metal2 14224 21560 14224 21560 0 _0754_
rlabel metal2 21896 28672 21896 28672 0 _0755_
rlabel metal2 21784 29288 21784 29288 0 _0756_
rlabel metal2 21280 28840 21280 28840 0 _0757_
rlabel metal2 15064 28896 15064 28896 0 _0758_
rlabel metal2 15736 29288 15736 29288 0 _0759_
rlabel metal3 13272 27720 13272 27720 0 _0760_
rlabel metal3 11760 27720 11760 27720 0 _0761_
rlabel metal2 11144 28728 11144 28728 0 _0762_
rlabel metal2 14056 26600 14056 26600 0 _0763_
rlabel metal2 13496 27608 13496 27608 0 _0764_
rlabel metal2 12712 29904 12712 29904 0 _0765_
rlabel metal2 11032 24304 11032 24304 0 _0766_
rlabel metal3 13328 25480 13328 25480 0 _0767_
rlabel metal2 12600 24584 12600 24584 0 _0768_
rlabel metal3 11536 25480 11536 25480 0 _0769_
rlabel metal3 10136 25480 10136 25480 0 _0770_
rlabel metal2 12544 24136 12544 24136 0 _0771_
rlabel metal3 13496 24136 13496 24136 0 _0772_
rlabel metal2 13496 24192 13496 24192 0 _0773_
rlabel metal2 11816 23912 11816 23912 0 _0774_
rlabel metal2 10808 23856 10808 23856 0 _0775_
rlabel metal2 10472 24024 10472 24024 0 _0776_
rlabel metal3 11536 21448 11536 21448 0 _0777_
rlabel metal3 10584 21672 10584 21672 0 _0778_
rlabel metal2 16240 20328 16240 20328 0 _0779_
rlabel metal2 14280 18704 14280 18704 0 _0780_
rlabel metal3 15232 19992 15232 19992 0 _0781_
rlabel metal2 12768 17640 12768 17640 0 _0782_
rlabel metal3 14448 19208 14448 19208 0 _0783_
rlabel metal2 15400 19768 15400 19768 0 _0784_
rlabel metal2 12152 19040 12152 19040 0 _0785_
rlabel metal2 25816 21280 25816 21280 0 _0786_
rlabel metal2 26040 20860 26040 20860 0 _0787_
rlabel metal3 40544 15400 40544 15400 0 _0788_
rlabel metal2 42056 15204 42056 15204 0 _0789_
rlabel metal2 40040 12544 40040 12544 0 _0790_
rlabel metal3 40824 13720 40824 13720 0 _0791_
rlabel metal2 42504 12432 42504 12432 0 _0792_
rlabel metal2 42448 11928 42448 11928 0 _0793_
rlabel metal3 43568 9800 43568 9800 0 _0794_
rlabel metal2 42504 8456 42504 8456 0 _0795_
rlabel metal2 45416 10640 45416 10640 0 _0796_
rlabel metal2 39256 8904 39256 8904 0 _0797_
rlabel metal2 40152 6832 40152 6832 0 _0798_
rlabel metal2 41720 11984 41720 11984 0 _0799_
rlabel metal2 39704 10528 39704 10528 0 _0800_
rlabel metal3 42504 12152 42504 12152 0 _0801_
rlabel metal3 43960 11592 43960 11592 0 _0802_
rlabel metal2 40376 21000 40376 21000 0 _0803_
rlabel metal2 40152 21056 40152 21056 0 _0804_
rlabel metal3 35896 17528 35896 17528 0 _0805_
rlabel metal2 39368 15456 39368 15456 0 _0806_
rlabel metal2 37688 14000 37688 14000 0 _0807_
rlabel metal2 38584 15904 38584 15904 0 _0808_
rlabel metal3 38808 14504 38808 14504 0 _0809_
rlabel metal2 39536 15288 39536 15288 0 _0810_
rlabel metal2 36344 21280 36344 21280 0 _0811_
rlabel metal3 39424 17640 39424 17640 0 _0812_
rlabel metal2 8232 24360 8232 24360 0 _0813_
rlabel metal2 24080 19208 24080 19208 0 _0814_
rlabel metal2 21336 19264 21336 19264 0 _0815_
rlabel metal2 21784 17360 21784 17360 0 _0816_
rlabel metal2 21336 16800 21336 16800 0 _0817_
rlabel metal2 21784 16576 21784 16576 0 _0818_
rlabel metal2 20888 17696 20888 17696 0 _0819_
rlabel metal2 22792 17640 22792 17640 0 _0820_
rlabel metal2 22008 19208 22008 19208 0 _0821_
rlabel metal2 44296 25872 44296 25872 0 _0822_
rlabel metal2 42952 25368 42952 25368 0 _0823_
rlabel metal2 44184 23800 44184 23800 0 _0824_
rlabel metal2 43400 24920 43400 24920 0 _0825_
rlabel metal2 44072 27832 44072 27832 0 _0826_
rlabel metal2 42840 28224 42840 28224 0 _0827_
rlabel metal2 43344 22456 43344 22456 0 _0828_
rlabel metal3 43960 24808 43960 24808 0 _0829_
rlabel metal2 47544 25816 47544 25816 0 _0830_
rlabel metal2 47880 25032 47880 25032 0 _0831_
rlabel metal2 46760 24920 46760 24920 0 _0832_
rlabel metal2 48664 24024 48664 24024 0 _0833_
rlabel metal2 47768 26684 47768 26684 0 _0834_
rlabel metal3 47824 26152 47824 26152 0 _0835_
rlabel metal2 31864 10976 31864 10976 0 _0836_
rlabel metal2 31416 10920 31416 10920 0 _0837_
rlabel metal2 33544 13104 33544 13104 0 _0838_
rlabel metal2 32928 12936 32928 12936 0 _0839_
rlabel metal2 32704 16632 32704 16632 0 _0840_
rlabel metal2 34216 14392 34216 14392 0 _0841_
rlabel metal2 41384 19880 41384 19880 0 _0842_
rlabel metal2 44856 19152 44856 19152 0 _0843_
rlabel metal3 43232 20664 43232 20664 0 _0844_
rlabel metal2 42616 18928 42616 18928 0 _0845_
rlabel metal2 41272 20832 41272 20832 0 _0846_
rlabel metal2 21896 5544 21896 5544 0 _0847_
rlabel metal2 21448 6328 21448 6328 0 _0848_
rlabel metal2 22456 5880 22456 5880 0 _0849_
rlabel metal2 16296 6440 16296 6440 0 _0850_
rlabel metal2 19096 5544 19096 5544 0 _0851_
rlabel metal2 20440 4872 20440 4872 0 _0852_
rlabel metal3 30520 12936 30520 12936 0 _0853_
rlabel metal2 31192 11368 31192 11368 0 _0854_
rlabel metal2 31864 12880 31864 12880 0 _0855_
rlabel metal2 31304 10920 31304 10920 0 _0856_
rlabel metal2 31528 13328 31528 13328 0 _0857_
rlabel metal2 28616 14504 28616 14504 0 _0858_
rlabel metal2 28448 11368 28448 11368 0 _0859_
rlabel metal3 26992 11144 26992 11144 0 _0860_
rlabel metal3 31920 15176 31920 15176 0 _0861_
rlabel metal2 31416 13160 31416 13160 0 _0862_
rlabel metal2 29456 10584 29456 10584 0 _0863_
rlabel metal2 26152 15904 26152 15904 0 _0864_
rlabel metal2 29288 15568 29288 15568 0 _0865_
rlabel metal2 28280 18368 28280 18368 0 _0866_
rlabel metal2 29624 10528 29624 10528 0 _0867_
rlabel metal2 24696 10304 24696 10304 0 _0868_
rlabel metal3 30296 7448 30296 7448 0 _0869_
rlabel metal2 28168 9744 28168 9744 0 _0870_
rlabel metal3 28672 8232 28672 8232 0 _0871_
rlabel metal2 30240 9128 30240 9128 0 _0872_
rlabel metal3 30408 9016 30408 9016 0 _0873_
rlabel metal4 6104 44744 6104 44744 0 _0874_
rlabel metal2 7224 33712 7224 33712 0 _0875_
rlabel metal2 8344 32088 8344 32088 0 _0876_
rlabel metal2 5992 39312 5992 39312 0 _0877_
rlabel metal2 7560 36456 7560 36456 0 _0878_
rlabel metal2 7896 34272 7896 34272 0 _0879_
rlabel metal2 7952 30968 7952 30968 0 _0880_
rlabel metal3 7280 31080 7280 31080 0 _0881_
rlabel metal2 5880 25256 5880 25256 0 _0882_
rlabel metal2 6048 28840 6048 28840 0 _0883_
rlabel metal2 6440 31024 6440 31024 0 _0884_
rlabel metal2 6496 33208 6496 33208 0 _0885_
rlabel metal3 7224 30856 7224 30856 0 _0886_
rlabel metal2 6440 30464 6440 30464 0 _0887_
rlabel metal3 7672 29400 7672 29400 0 _0888_
rlabel metal2 8232 25200 8232 25200 0 _0889_
rlabel metal3 7560 46760 7560 46760 0 _0890_
rlabel metal2 6776 46648 6776 46648 0 _0891_
rlabel metal2 5656 29400 5656 29400 0 _0892_
rlabel metal2 4032 43288 4032 43288 0 _0893_
rlabel metal3 5264 43624 5264 43624 0 _0894_
rlabel metal3 6104 45752 6104 45752 0 _0895_
rlabel metal3 5432 43400 5432 43400 0 _0896_
rlabel metal2 6608 42728 6608 42728 0 _0897_
rlabel metal2 7112 43568 7112 43568 0 _0898_
rlabel metal2 9912 44072 9912 44072 0 _0899_
rlabel metal2 8904 43008 8904 43008 0 _0900_
rlabel metal2 8232 42280 8232 42280 0 _0901_
rlabel metal2 10584 40656 10584 40656 0 _0902_
rlabel metal2 10920 41888 10920 41888 0 _0903_
rlabel metal3 9016 42952 9016 42952 0 _0904_
rlabel metal3 9464 43288 9464 43288 0 _0905_
rlabel metal2 2744 37968 2744 37968 0 _0906_
rlabel metal3 6160 43288 6160 43288 0 _0907_
rlabel metal2 5096 40432 5096 40432 0 _0908_
rlabel metal2 2968 40320 2968 40320 0 _0909_
rlabel metal2 6272 39592 6272 39592 0 _0910_
rlabel metal2 6664 40656 6664 40656 0 _0911_
rlabel metal2 7448 40264 7448 40264 0 _0912_
rlabel metal2 5880 39144 5880 39144 0 _0913_
rlabel metal2 5656 39760 5656 39760 0 _0914_
rlabel metal2 2968 38472 2968 38472 0 _0915_
rlabel metal2 8568 39032 8568 39032 0 _0916_
rlabel metal2 8904 39816 8904 39816 0 _0917_
rlabel metal2 9800 39480 9800 39480 0 _0918_
rlabel metal3 8288 38808 8288 38808 0 _0919_
rlabel metal2 6552 36288 6552 36288 0 _0920_
rlabel via2 8120 36568 8120 36568 0 _0921_
rlabel metal2 10920 37296 10920 37296 0 _0922_
rlabel metal2 8344 29456 8344 29456 0 _0923_
rlabel metal2 9240 35672 9240 35672 0 _0924_
rlabel metal3 8680 35112 8680 35112 0 _0925_
rlabel metal2 11032 33040 11032 33040 0 _0926_
rlabel metal2 7336 33264 7336 33264 0 _0927_
rlabel metal2 7448 30800 7448 30800 0 _0928_
rlabel metal2 7112 31752 7112 31752 0 _0929_
rlabel metal2 10808 31696 10808 31696 0 _0930_
rlabel metal2 7112 27552 7112 27552 0 _0931_
rlabel metal2 4872 25760 4872 25760 0 _0932_
rlabel metal2 8680 28504 8680 28504 0 _0933_
rlabel metal3 5320 25592 5320 25592 0 _0934_
rlabel metal2 4592 23128 4592 23128 0 _0935_
rlabel via2 4872 23800 4872 23800 0 _0936_
rlabel metal3 4704 23128 4704 23128 0 _0937_
rlabel metal2 2856 22344 2856 22344 0 _0938_
rlabel metal2 6104 24080 6104 24080 0 _0939_
rlabel metal3 7392 25368 7392 25368 0 _0940_
rlabel metal3 7784 25480 7784 25480 0 _0941_
rlabel metal2 5320 25872 5320 25872 0 _0942_
rlabel metal2 5208 26656 5208 26656 0 _0943_
rlabel metal2 3304 27160 3304 27160 0 _0944_
rlabel metal2 3304 29008 3304 29008 0 _0945_
rlabel metal2 5320 29848 5320 29848 0 _0946_
rlabel metal2 3976 28672 3976 28672 0 _0947_
rlabel metal2 2632 27888 2632 27888 0 _0948_
rlabel metal2 3080 30576 3080 30576 0 _0949_
rlabel metal2 3304 30184 3304 30184 0 _0950_
rlabel metal3 3360 30968 3360 30968 0 _0951_
rlabel metal2 2184 30856 2184 30856 0 _0952_
rlabel metal2 2968 33992 2968 33992 0 _0953_
rlabel metal2 3080 36232 3080 36232 0 _0954_
rlabel metal2 2632 37464 2632 37464 0 _0955_
rlabel metal2 2520 35280 2520 35280 0 _0956_
rlabel metal2 2632 35280 2632 35280 0 _0957_
rlabel metal2 2744 34496 2744 34496 0 _0958_
rlabel metal3 2520 32424 2520 32424 0 _0959_
rlabel metal2 3304 33208 3304 33208 0 _0960_
rlabel metal2 4424 33992 4424 33992 0 _0961_
rlabel metal2 4032 34216 4032 34216 0 _0962_
rlabel metal2 4536 34216 4536 34216 0 _0963_
rlabel metal3 43008 38920 43008 38920 0 _0964_
rlabel metal2 37072 20776 37072 20776 0 _0965_
rlabel metal2 35504 21000 35504 21000 0 _0966_
rlabel metal3 35392 23016 35392 23016 0 _0967_
rlabel metal2 38920 16520 38920 16520 0 _0968_
rlabel metal3 41160 18424 41160 18424 0 _0969_
rlabel metal2 37128 17976 37128 17976 0 _0970_
rlabel metal3 34888 16968 34888 16968 0 _0971_
rlabel metal2 36568 25116 36568 25116 0 _0972_
rlabel metal2 36120 31472 36120 31472 0 _0973_
rlabel metal3 34832 23352 34832 23352 0 _0974_
rlabel metal2 39256 22736 39256 22736 0 _0975_
rlabel metal2 40152 35952 40152 35952 0 _0976_
rlabel metal2 36568 30072 36568 30072 0 _0977_
rlabel metal2 35784 31416 35784 31416 0 _0978_
rlabel metal3 34832 31864 34832 31864 0 _0979_
rlabel metal3 41272 38696 41272 38696 0 _0980_
rlabel metal2 35000 29680 35000 29680 0 _0981_
rlabel metal2 39032 43568 39032 43568 0 _0982_
rlabel metal3 33824 32424 33824 32424 0 _0983_
rlabel metal2 25928 40712 25928 40712 0 _0984_
rlabel metal2 38472 32144 38472 32144 0 _0985_
rlabel metal2 23576 41776 23576 41776 0 _0986_
rlabel metal2 36344 30856 36344 30856 0 _0987_
rlabel metal2 29512 13160 29512 13160 0 _0988_
rlabel metal2 20216 22904 20216 22904 0 _0989_
rlabel metal2 38248 14392 38248 14392 0 _0990_
rlabel metal2 34552 16912 34552 16912 0 _0991_
rlabel metal3 22008 20664 22008 20664 0 _0992_
rlabel metal2 20440 21056 20440 21056 0 _0993_
rlabel metal2 27104 13720 27104 13720 0 _0994_
rlabel metal2 21224 15848 21224 15848 0 _0995_
rlabel metal2 21448 22512 21448 22512 0 _0996_
rlabel metal2 21784 20944 21784 20944 0 _0997_
rlabel metal2 21448 21336 21448 21336 0 _0998_
rlabel metal2 21000 21560 21000 21560 0 _0999_
rlabel metal2 18984 22344 18984 22344 0 _1000_
rlabel metal2 22904 19432 22904 19432 0 _1001_
rlabel metal2 26824 8316 26824 8316 0 _1002_
rlabel metal2 28280 20384 28280 20384 0 _1003_
rlabel metal2 23352 20664 23352 20664 0 _1004_
rlabel metal2 22904 21784 22904 21784 0 _1005_
rlabel metal3 23408 20104 23408 20104 0 _1006_
rlabel metal2 21448 11200 21448 11200 0 _1007_
rlabel metal2 29344 5096 29344 5096 0 _1008_
rlabel metal2 30744 4648 30744 4648 0 _1009_
rlabel metal2 30184 16296 30184 16296 0 _1010_
rlabel metal2 37128 9856 37128 9856 0 _1011_
rlabel metal2 30856 7056 30856 7056 0 _1012_
rlabel metal2 30856 8232 30856 8232 0 _1013_
rlabel metal2 30296 7840 30296 7840 0 _1014_
rlabel metal2 29568 6664 29568 6664 0 _1015_
rlabel metal2 30576 6888 30576 6888 0 _1016_
rlabel metal2 28056 7000 28056 7000 0 _1017_
rlabel metal3 28896 7448 28896 7448 0 _1018_
rlabel metal2 27496 5488 27496 5488 0 _1019_
rlabel metal2 26488 4704 26488 4704 0 _1020_
rlabel metal2 23016 7784 23016 7784 0 _1021_
rlabel via2 25704 4424 25704 4424 0 _1022_
rlabel metal3 25368 4088 25368 4088 0 _1023_
rlabel metal2 25816 7000 25816 7000 0 _1024_
rlabel metal3 26096 7336 26096 7336 0 _1025_
rlabel metal2 25928 7336 25928 7336 0 _1026_
rlabel metal2 25368 7616 25368 7616 0 _1027_
rlabel metal2 23856 9016 23856 9016 0 _1028_
rlabel metal3 24192 8232 24192 8232 0 _1029_
rlabel metal3 25032 9240 25032 9240 0 _1030_
rlabel metal2 25592 7896 25592 7896 0 _1031_
rlabel metal3 23464 8008 23464 8008 0 _1032_
rlabel metal2 23800 6328 23800 6328 0 _1033_
rlabel metal2 23240 11816 23240 11816 0 _1034_
rlabel metal3 22232 8904 22232 8904 0 _1035_
rlabel metal2 25928 4424 25928 4424 0 _1036_
rlabel metal2 15624 6608 15624 6608 0 _1037_
rlabel metal3 21056 8232 21056 8232 0 _1038_
rlabel metal2 17976 7056 17976 7056 0 _1039_
rlabel metal2 24472 6552 24472 6552 0 _1040_
rlabel metal2 35784 7392 35784 7392 0 _1041_
rlabel metal3 34160 8120 34160 8120 0 _1042_
rlabel metal3 36568 6664 36568 6664 0 _1043_
rlabel metal3 36960 6552 36960 6552 0 _1044_
rlabel metal2 36120 7448 36120 7448 0 _1045_
rlabel metal3 40712 7448 40712 7448 0 _1046_
rlabel metal2 34776 7896 34776 7896 0 _1047_
rlabel metal2 31640 8736 31640 8736 0 _1048_
rlabel metal3 40376 7336 40376 7336 0 _1049_
rlabel metal2 34832 7448 34832 7448 0 _1050_
rlabel metal2 27496 9800 27496 9800 0 _1051_
rlabel metal2 32368 10808 32368 10808 0 _1052_
rlabel metal2 39256 7728 39256 7728 0 _1053_
rlabel metal3 24696 21784 24696 21784 0 _1054_
rlabel metal2 22008 5880 22008 5880 0 _1055_
rlabel metal2 12208 2968 12208 2968 0 _1056_
rlabel metal2 38360 6496 38360 6496 0 _1057_
rlabel metal2 43960 4816 43960 4816 0 _1058_
rlabel metal2 47432 5264 47432 5264 0 _1059_
rlabel metal2 36904 6720 36904 6720 0 _1060_
rlabel metal2 43288 6832 43288 6832 0 _1061_
rlabel metal2 48104 9072 48104 9072 0 _1062_
rlabel metal2 45528 8512 45528 8512 0 _1063_
rlabel metal3 35224 4424 35224 4424 0 _1064_
rlabel metal2 49000 7504 49000 7504 0 _1065_
rlabel metal2 46872 6832 46872 6832 0 _1066_
rlabel metal2 47768 9296 47768 9296 0 _1067_
rlabel metal2 46704 9240 46704 9240 0 _1068_
rlabel metal2 45416 7000 45416 7000 0 _1069_
rlabel metal2 25536 12376 25536 12376 0 _1070_
rlabel metal2 25816 10136 25816 10136 0 _1071_
rlabel metal2 24472 12488 24472 12488 0 _1072_
rlabel metal3 25144 12040 25144 12040 0 _1073_
rlabel metal2 21672 12824 21672 12824 0 _1074_
rlabel metal3 22456 12824 22456 12824 0 _1075_
rlabel metal3 18872 14280 18872 14280 0 _1076_
rlabel metal2 17304 13608 17304 13608 0 _1077_
rlabel metal2 22120 11592 22120 11592 0 _1078_
rlabel metal2 18872 13552 18872 13552 0 _1079_
rlabel metal2 15400 11368 15400 11368 0 _1080_
rlabel metal2 15848 12432 15848 12432 0 _1081_
rlabel metal2 18032 26040 18032 26040 0 _1082_
rlabel metal2 16632 12880 16632 12880 0 _1083_
rlabel metal3 17080 12152 17080 12152 0 _1084_
rlabel metal2 15064 11480 15064 11480 0 _1085_
rlabel metal2 25312 21560 25312 21560 0 _1086_
rlabel metal2 16408 9352 16408 9352 0 _1087_
rlabel metal2 33432 17136 33432 17136 0 _1088_
rlabel metal2 24136 40600 24136 40600 0 _1089_
rlabel metal2 26152 39704 26152 39704 0 _1090_
rlabel metal2 24136 38808 24136 38808 0 _1091_
rlabel metal2 26600 39480 26600 39480 0 _1092_
rlabel metal3 25088 37128 25088 37128 0 _1093_
rlabel metal2 26600 37688 26600 37688 0 _1094_
rlabel metal2 26712 39648 26712 39648 0 _1095_
rlabel metal2 24472 40320 24472 40320 0 _1096_
rlabel metal2 22568 43400 22568 43400 0 _1097_
rlabel metal2 22904 39704 22904 39704 0 _1098_
rlabel metal2 23016 40824 23016 40824 0 _1099_
rlabel metal2 23912 25592 23912 25592 0 _1100_
rlabel metal2 23128 42840 23128 42840 0 _1101_
rlabel metal3 22120 26488 22120 26488 0 _1102_
rlabel metal3 21336 44184 21336 44184 0 _1103_
rlabel metal2 22232 25648 22232 25648 0 _1104_
rlabel metal3 21168 42616 21168 42616 0 _1105_
rlabel metal3 37856 20776 37856 20776 0 _1106_
rlabel metal2 34216 20944 34216 20944 0 _1107_
rlabel metal2 38360 21784 38360 21784 0 _1108_
rlabel metal2 31528 23408 31528 23408 0 _1109_
rlabel metal2 26376 22736 26376 22736 0 _1110_
rlabel metal3 31752 24696 31752 24696 0 _1111_
rlabel metal2 27608 23912 27608 23912 0 _1112_
rlabel metal2 27048 21504 27048 21504 0 _1113_
rlabel metal2 30856 24528 30856 24528 0 _1114_
rlabel metal2 29848 24192 29848 24192 0 _1115_
rlabel metal2 31136 23128 31136 23128 0 _1116_
rlabel metal2 28728 38724 28728 38724 0 _1117_
rlabel metal2 40712 37744 40712 37744 0 _1118_
rlabel metal2 31304 37072 31304 37072 0 _1119_
rlabel metal2 35504 39592 35504 39592 0 _1120_
rlabel metal3 36288 38136 36288 38136 0 _1121_
rlabel metal2 32536 37576 32536 37576 0 _1122_
rlabel metal2 33096 39928 33096 39928 0 _1123_
rlabel metal3 36848 39480 36848 39480 0 _1124_
rlabel metal2 29960 43120 29960 43120 0 _1125_
rlabel metal2 30464 42504 30464 42504 0 _1126_
rlabel metal2 30184 43120 30184 43120 0 _1127_
rlabel metal3 29008 39368 29008 39368 0 _1128_
rlabel metal2 24584 42672 24584 42672 0 _1129_
rlabel metal2 26376 42000 26376 42000 0 _1130_
rlabel metal2 35000 6328 35000 6328 0 _1131_
rlabel metal3 31976 8792 31976 8792 0 _1132_
rlabel metal2 32312 7840 32312 7840 0 _1133_
rlabel metal3 37968 11368 37968 11368 0 _1134_
rlabel metal2 36120 10528 36120 10528 0 _1135_
rlabel metal2 32200 9576 32200 9576 0 _1136_
rlabel metal3 32480 7448 32480 7448 0 _1137_
rlabel metal2 34104 5488 34104 5488 0 _1138_
rlabel metal2 32648 7560 32648 7560 0 _1139_
rlabel metal2 21672 9744 21672 9744 0 _1140_
rlabel metal2 22792 9744 22792 9744 0 _1141_
rlabel metal2 18872 9632 18872 9632 0 _1142_
rlabel metal2 19768 11480 19768 11480 0 _1143_
rlabel metal2 18312 9408 18312 9408 0 _1144_
rlabel metal2 18760 8792 18760 8792 0 _1145_
rlabel metal2 11872 10024 11872 10024 0 _1146_
rlabel metal2 11032 9856 11032 9856 0 _1147_
rlabel metal2 11536 9240 11536 9240 0 _1148_
rlabel metal2 13160 8680 13160 8680 0 _1149_
rlabel metal3 11368 7672 11368 7672 0 _1150_
rlabel metal3 10304 8120 10304 8120 0 _1151_
rlabel metal3 13552 6664 13552 6664 0 _1152_
rlabel metal2 13944 8680 13944 8680 0 _1153_
rlabel metal2 15008 8120 15008 8120 0 _1154_
rlabel metal2 15624 8456 15624 8456 0 _1155_
rlabel metal2 8680 9352 8680 9352 0 _1156_
rlabel metal2 7560 9800 7560 9800 0 _1157_
rlabel metal2 7840 7560 7840 7560 0 _1158_
rlabel metal2 7448 8232 7448 8232 0 _1159_
rlabel metal2 7504 6440 7504 6440 0 _1160_
rlabel metal2 10248 11480 10248 11480 0 _1161_
rlabel metal2 7448 6944 7448 6944 0 _1162_
rlabel metal2 8568 4704 8568 4704 0 _1163_
rlabel metal2 8344 4032 8344 4032 0 _1164_
rlabel metal3 9744 3752 9744 3752 0 _1165_
rlabel metal2 11704 4032 11704 4032 0 _1166_
rlabel metal2 9576 4312 9576 4312 0 _1167_
rlabel metal2 12264 3696 12264 3696 0 _1168_
rlabel metal2 13272 4424 13272 4424 0 _1169_
rlabel metal2 14784 5096 14784 5096 0 _1170_
rlabel metal2 17080 5824 17080 5824 0 _1171_
rlabel metal2 39704 21448 39704 21448 0 _1172_
rlabel metal2 38416 21000 38416 21000 0 _1173_
rlabel metal2 26488 15736 26488 15736 0 _1174_
rlabel metal2 27160 15736 27160 15736 0 _1175_
rlabel metal2 24752 23016 24752 23016 0 _1176_
rlabel metal2 31640 11284 31640 11284 0 _1177_
rlabel metal2 28392 15344 28392 15344 0 _1178_
rlabel metal2 39144 24640 39144 24640 0 _1179_
rlabel metal2 39032 39312 39032 39312 0 _1180_
rlabel metal2 38024 40264 38024 40264 0 _1181_
rlabel metal2 39256 40040 39256 40040 0 _1182_
rlabel metal3 40432 37128 40432 37128 0 _1183_
rlabel metal2 38808 37128 38808 37128 0 _1184_
rlabel metal3 39704 38696 39704 38696 0 _1185_
rlabel metal2 41272 39424 41272 39424 0 _1186_
rlabel metal2 39368 41776 39368 41776 0 _1187_
rlabel metal3 40488 42168 40488 42168 0 _1188_
rlabel metal2 36792 43904 36792 43904 0 _1189_
rlabel metal2 7784 23856 7784 23856 0 blink.LED
rlabel metal2 6048 44968 6048 44968 0 blink.counter\[0\]
rlabel metal2 5768 40880 5768 40880 0 blink.counter\[10\]
rlabel metal2 7672 40432 7672 40432 0 blink.counter\[11\]
rlabel metal2 7784 39256 7784 39256 0 blink.counter\[12\]
rlabel metal3 9184 35672 9184 35672 0 blink.counter\[13\]
rlabel metal3 11088 36456 11088 36456 0 blink.counter\[14\]
rlabel metal2 10528 34104 10528 34104 0 blink.counter\[15\]
rlabel metal2 10808 32592 10808 32592 0 blink.counter\[16\]
rlabel metal2 9912 31584 9912 31584 0 blink.counter\[17\]
rlabel metal2 10472 32088 10472 32088 0 blink.counter\[18\]
rlabel metal2 7784 28224 7784 28224 0 blink.counter\[19\]
rlabel metal2 7112 46592 7112 46592 0 blink.counter\[1\]
rlabel metal2 5096 25312 5096 25312 0 blink.counter\[20\]
rlabel metal2 4648 22512 4648 22512 0 blink.counter\[21\]
rlabel metal2 5208 24304 5208 24304 0 blink.counter\[22\]
rlabel metal2 8680 25816 8680 25816 0 blink.counter\[23\]
rlabel metal2 4648 26208 4648 26208 0 blink.counter\[24\]
rlabel metal3 5096 29400 5096 29400 0 blink.counter\[25\]
rlabel metal2 4872 28728 4872 28728 0 blink.counter\[26\]
rlabel metal2 2352 31192 2352 31192 0 blink.counter\[27\]
rlabel metal2 2296 36960 2296 36960 0 blink.counter\[28\]
rlabel metal2 6048 33544 6048 33544 0 blink.counter\[29\]
rlabel metal3 5992 44968 5992 44968 0 blink.counter\[2\]
rlabel metal2 6216 34552 6216 34552 0 blink.counter\[30\]
rlabel metal2 7336 34608 7336 34608 0 blink.counter\[31\]
rlabel metal2 5768 44016 5768 44016 0 blink.counter\[3\]
rlabel metal3 11648 43512 11648 43512 0 blink.counter\[4\]
rlabel via2 11480 42728 11480 42728 0 blink.counter\[5\]
rlabel metal2 12824 41776 12824 41776 0 blink.counter\[6\]
rlabel metal2 5320 43288 5320 43288 0 blink.counter\[7\]
rlabel metal2 4648 40824 4648 40824 0 blink.counter\[8\]
rlabel metal2 6104 40152 6104 40152 0 blink.counter\[9\]
rlabel metal2 18760 19544 18760 19544 0 clknet_0_wb_clk_i
rlabel metal2 22680 7112 22680 7112 0 clknet_2_0__leaf_wb_clk_i
rlabel metal2 23296 41944 23296 41944 0 clknet_2_1__leaf_wb_clk_i
rlabel metal2 22232 15512 22232 15512 0 clknet_2_2__leaf_wb_clk_i
rlabel metal2 38808 23352 38808 23352 0 clknet_2_3__leaf_wb_clk_i
rlabel metal2 12712 21952 12712 21952 0 clknet_leaf_0_wb_clk_i
rlabel metal2 23912 45472 23912 45472 0 clknet_leaf_10_wb_clk_i
rlabel metal2 20888 34160 20888 34160 0 clknet_leaf_11_wb_clk_i
rlabel metal2 24584 31360 24584 31360 0 clknet_leaf_12_wb_clk_i
rlabel metal2 31976 36736 31976 36736 0 clknet_leaf_13_wb_clk_i
rlabel metal2 26264 38808 26264 38808 0 clknet_leaf_14_wb_clk_i
rlabel metal2 28952 45472 28952 45472 0 clknet_leaf_15_wb_clk_i
rlabel metal2 39256 42336 39256 42336 0 clknet_leaf_16_wb_clk_i
rlabel metal2 45304 45528 45304 45528 0 clknet_leaf_17_wb_clk_i
rlabel metal2 46424 40768 46424 40768 0 clknet_leaf_18_wb_clk_i
rlabel metal2 45304 35224 45304 35224 0 clknet_leaf_19_wb_clk_i
rlabel metal2 20832 23912 20832 23912 0 clknet_leaf_1_wb_clk_i
rlabel metal2 45416 26152 45416 26152 0 clknet_leaf_20_wb_clk_i
rlabel metal2 39256 26572 39256 26572 0 clknet_leaf_21_wb_clk_i
rlabel metal2 36232 31304 36232 31304 0 clknet_leaf_22_wb_clk_i
rlabel metal2 33208 24920 33208 24920 0 clknet_leaf_23_wb_clk_i
rlabel metal2 39592 18368 39592 18368 0 clknet_leaf_24_wb_clk_i
rlabel metal2 43512 24304 43512 24304 0 clknet_leaf_25_wb_clk_i
rlabel metal2 46312 18032 46312 18032 0 clknet_leaf_26_wb_clk_i
rlabel metal2 44856 3920 44856 3920 0 clknet_leaf_27_wb_clk_i
rlabel metal2 38248 7112 38248 7112 0 clknet_leaf_28_wb_clk_i
rlabel metal2 37576 10752 37576 10752 0 clknet_leaf_29_wb_clk_i
rlabel metal2 17528 30520 17528 30520 0 clknet_leaf_2_wb_clk_i
rlabel metal2 27832 5096 27832 5096 0 clknet_leaf_30_wb_clk_i
rlabel metal3 31640 11760 31640 11760 0 clknet_leaf_31_wb_clk_i
rlabel metal2 29288 14112 29288 14112 0 clknet_leaf_32_wb_clk_i
rlabel metal2 25368 22400 25368 22400 0 clknet_leaf_33_wb_clk_i
rlabel metal2 23632 11368 23632 11368 0 clknet_leaf_34_wb_clk_i
rlabel metal2 23464 7448 23464 7448 0 clknet_leaf_35_wb_clk_i
rlabel metal2 17752 7000 17752 7000 0 clknet_leaf_36_wb_clk_i
rlabel metal2 8792 9744 8792 9744 0 clknet_leaf_37_wb_clk_i
rlabel metal2 10024 5432 10024 5432 0 clknet_leaf_38_wb_clk_i
rlabel metal2 1848 11424 1848 11424 0 clknet_leaf_39_wb_clk_i
rlabel metal3 4032 26264 4032 26264 0 clknet_leaf_3_wb_clk_i
rlabel metal2 8008 16912 8008 16912 0 clknet_leaf_40_wb_clk_i
rlabel metal2 1848 16520 1848 16520 0 clknet_leaf_41_wb_clk_i
rlabel metal2 6272 23128 6272 23128 0 clknet_leaf_42_wb_clk_i
rlabel metal2 1848 30968 1848 30968 0 clknet_leaf_4_wb_clk_i
rlabel metal2 9912 35224 9912 35224 0 clknet_leaf_5_wb_clk_i
rlabel metal2 1848 44688 1848 44688 0 clknet_leaf_6_wb_clk_i
rlabel metal2 9016 44744 9016 44744 0 clknet_leaf_7_wb_clk_i
rlabel metal2 13608 42336 13608 42336 0 clknet_leaf_8_wb_clk_i
rlabel metal2 21672 45920 21672 45920 0 clknet_leaf_9_wb_clk_i
rlabel metal2 49280 41944 49280 41944 0 custom_settings[0]
rlabel metal2 49112 47376 49112 47376 0 custom_settings[1]
rlabel metal2 48216 47712 48216 47712 0 custom_settings[3]
rlabel metal3 50106 2072 50106 2072 0 io_in_1[0]
rlabel metal3 28000 2744 28000 2744 0 io_in_1[1]
rlabel metal3 26040 9968 26040 9968 0 io_in_1[2]
rlabel metal2 17080 22512 17080 22512 0 io_in_1[3]
rlabel metal3 20160 22960 20160 22960 0 io_in_1[4]
rlabel metal2 48104 24024 48104 24024 0 io_in_1[5]
rlabel metal4 46312 34720 46312 34720 0 io_in_1[6]
rlabel metal2 42000 39928 42000 39928 0 io_in_1[7]
rlabel metal2 31640 47824 31640 47824 0 io_in_2[0]
rlabel metal2 44856 47824 44856 47824 0 io_in_2[1]
rlabel metal2 19096 2030 19096 2030 0 io_out[10]
rlabel metal2 20888 854 20888 854 0 io_out[11]
rlabel metal2 31640 2198 31640 2198 0 io_out[17]
rlabel metal2 33432 2198 33432 2198 0 io_out[18]
rlabel metal2 35224 2254 35224 2254 0 io_out[19]
rlabel metal2 37016 2422 37016 2422 0 io_out[20]
rlabel metal2 38808 2814 38808 2814 0 io_out[21]
rlabel metal2 15512 2030 15512 2030 0 io_out[8]
rlabel metal2 17304 854 17304 854 0 io_out[9]
rlabel metal3 21560 21616 21560 21616 0 net1
rlabel metal2 47656 26544 47656 26544 0 net10
rlabel metal3 43736 26376 43736 26376 0 net11
rlabel metal2 23912 17472 23912 17472 0 net12
rlabel metal2 26264 21868 26264 21868 0 net13
rlabel metal2 15456 24920 15456 24920 0 net14
rlabel metal2 19712 3528 19712 3528 0 net15
rlabel metal2 21056 5096 21056 5096 0 net16
rlabel metal2 31416 4872 31416 4872 0 net17
rlabel metal2 35112 3584 35112 3584 0 net18
rlabel metal2 38976 3640 38976 3640 0 net19
rlabel metal3 43400 15960 43400 15960 0 net2
rlabel metal2 31640 7560 31640 7560 0 net20
rlabel metal3 31500 9128 31500 9128 0 net21
rlabel metal2 21784 5040 21784 5040 0 net22
rlabel metal3 17136 4312 17136 4312 0 net23
rlabel metal2 1176 2030 1176 2030 0 net24
rlabel metal2 2968 2030 2968 2030 0 net25
rlabel metal2 4760 2030 4760 2030 0 net26
rlabel metal2 6552 1190 6552 1190 0 net27
rlabel metal2 8344 1246 8344 1246 0 net28
rlabel metal2 10136 2030 10136 2030 0 net29
rlabel metal3 22344 6552 22344 6552 0 net3
rlabel metal2 8288 3304 8288 3304 0 net30
rlabel metal3 11256 3528 11256 3528 0 net31
rlabel metal2 22680 1470 22680 1470 0 net32
rlabel metal2 24472 2030 24472 2030 0 net33
rlabel metal2 26264 1582 26264 1582 0 net34
rlabel metal2 28056 2590 28056 2590 0 net35
rlabel metal2 29848 2086 29848 2086 0 net36
rlabel metal2 42392 2030 42392 2030 0 net37
rlabel metal2 44184 2058 44184 2058 0 net38
rlabel metal3 45472 4872 45472 4872 0 net39
rlabel metal2 21112 12432 21112 12432 0 net4
rlabel metal2 47712 3976 47712 3976 0 net40
rlabel metal3 48440 10248 48440 10248 0 net41
rlabel metal3 42728 4536 42728 4536 0 net42
rlabel metal2 24640 18312 24640 18312 0 net5
rlabel metal2 41272 9688 41272 9688 0 net6
rlabel metal2 26264 17136 26264 17136 0 net7
rlabel metal2 43848 20048 43848 20048 0 net8
rlabel metal2 43400 17864 43400 17864 0 net9
rlabel metal2 19096 48874 19096 48874 0 rst_n
rlabel metal3 39032 15400 39032 15400 0 tt_um_rejunity_ay8913.active
rlabel metal2 27496 16240 27496 16240 0 tt_um_rejunity_ay8913.amplitude_A\[0\]
rlabel metal2 33544 14448 33544 14448 0 tt_um_rejunity_ay8913.amplitude_B\[0\]
rlabel metal2 33096 11928 33096 11928 0 tt_um_rejunity_ay8913.amplitude_C\[0\]
rlabel metal2 41944 15792 41944 15792 0 tt_um_rejunity_ay8913.clk_counter\[0\]
rlabel metal2 41608 13160 41608 13160 0 tt_um_rejunity_ay8913.clk_counter\[1\]
rlabel metal2 42280 13608 42280 13608 0 tt_um_rejunity_ay8913.clk_counter\[2\]
rlabel metal3 42672 10696 42672 10696 0 tt_um_rejunity_ay8913.clk_counter\[3\]
rlabel metal2 41720 10136 41720 10136 0 tt_um_rejunity_ay8913.clk_counter\[4\]
rlabel metal3 42448 10360 42448 10360 0 tt_um_rejunity_ay8913.clk_counter\[5\]
rlabel metal2 41944 11368 41944 11368 0 tt_um_rejunity_ay8913.clk_counter\[6\]
rlabel metal4 28280 17696 28280 17696 0 tt_um_rejunity_ay8913.envelope_A
rlabel metal2 32088 13272 32088 13272 0 tt_um_rejunity_ay8913.envelope_B
rlabel metal2 27944 12544 27944 12544 0 tt_um_rejunity_ay8913.envelope_C
rlabel metal2 42280 19824 42280 19824 0 tt_um_rejunity_ay8913.envelope_alternate
rlabel metal2 45752 17976 45752 17976 0 tt_um_rejunity_ay8913.envelope_attack
rlabel metal3 43288 20104 43288 20104 0 tt_um_rejunity_ay8913.envelope_continue
rlabel metal2 46312 15596 46312 15596 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\]
rlabel metal2 47768 14224 47768 14224 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\]
rlabel metal2 47768 12600 47768 12600 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\]
rlabel metal2 47376 12936 47376 12936 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\]
rlabel metal2 43736 20104 43736 20104 0 tt_um_rejunity_ay8913.envelope_generator.hold
rlabel metal2 45976 16912 45976 16912 0 tt_um_rejunity_ay8913.envelope_generator.invert_output
rlabel metal2 42952 30296 42952 30296 0 tt_um_rejunity_ay8913.envelope_generator.period\[0\]
rlabel metal3 40656 40488 40656 40488 0 tt_um_rejunity_ay8913.envelope_generator.period\[10\]
rlabel metal2 41720 42000 41720 42000 0 tt_um_rejunity_ay8913.envelope_generator.period\[11\]
rlabel metal2 40488 44240 40488 44240 0 tt_um_rejunity_ay8913.envelope_generator.period\[12\]
rlabel metal2 40096 44968 40096 44968 0 tt_um_rejunity_ay8913.envelope_generator.period\[13\]
rlabel metal2 41216 45192 41216 45192 0 tt_um_rejunity_ay8913.envelope_generator.period\[14\]
rlabel metal2 40376 43288 40376 43288 0 tt_um_rejunity_ay8913.envelope_generator.period\[15\]
rlabel metal2 41608 31024 41608 31024 0 tt_um_rejunity_ay8913.envelope_generator.period\[1\]
rlabel metal3 42168 25368 42168 25368 0 tt_um_rejunity_ay8913.envelope_generator.period\[2\]
rlabel metal2 42280 24864 42280 24864 0 tt_um_rejunity_ay8913.envelope_generator.period\[3\]
rlabel metal2 45864 25312 45864 25312 0 tt_um_rejunity_ay8913.envelope_generator.period\[4\]
rlabel metal2 48888 23800 48888 23800 0 tt_um_rejunity_ay8913.envelope_generator.period\[5\]
rlabel metal3 48664 27160 48664 27160 0 tt_um_rejunity_ay8913.envelope_generator.period\[6\]
rlabel metal3 48664 25592 48664 25592 0 tt_um_rejunity_ay8913.envelope_generator.period\[7\]
rlabel metal2 43736 38080 43736 38080 0 tt_um_rejunity_ay8913.envelope_generator.period\[8\]
rlabel metal2 43456 38808 43456 38808 0 tt_um_rejunity_ay8913.envelope_generator.period\[9\]
rlabel metal2 49224 19040 49224 19040 0 tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
rlabel metal2 49224 21392 49224 21392 0 tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal
rlabel metal2 49224 17808 49224 17808 0 tt_um_rejunity_ay8913.envelope_generator.stop
rlabel metal2 39592 34048 39592 34048 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\]
rlabel metal3 46760 41272 46760 41272 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\]
rlabel metal2 47880 46312 47880 46312 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\]
rlabel metal2 46368 47432 46368 47432 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\]
rlabel metal2 43064 46648 43064 46648 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\]
rlabel metal2 43848 46032 43848 46032 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\]
rlabel metal2 44128 42840 44128 42840 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\]
rlabel metal2 40936 30576 40936 30576 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\]
rlabel metal2 43848 35056 43848 35056 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\]
rlabel metal2 44296 32368 44296 32368 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\]
rlabel metal2 45080 32984 45080 32984 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\]
rlabel metal3 48496 30968 48496 30968 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\]
rlabel metal2 49224 37016 49224 37016 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\]
rlabel metal3 48776 31864 48776 31864 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\]
rlabel metal2 44856 37184 44856 37184 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\]
rlabel metal2 49168 39704 49168 39704 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\]
rlabel metal2 36680 17640 36680 17640 0 tt_um_rejunity_ay8913.latched_register\[0\]
rlabel metal2 41048 16800 41048 16800 0 tt_um_rejunity_ay8913.latched_register\[1\]
rlabel metal2 35560 21504 35560 21504 0 tt_um_rejunity_ay8913.latched_register\[2\]
rlabel metal2 40040 21840 40040 21840 0 tt_um_rejunity_ay8913.latched_register\[3\]
rlabel metal3 28280 17528 28280 17528 0 tt_um_rejunity_ay8913.noise_disable_A
rlabel metal2 32200 14868 32200 14868 0 tt_um_rejunity_ay8913.noise_disable_B
rlabel metal2 34552 17976 34552 17976 0 tt_um_rejunity_ay8913.noise_disable_C
rlabel metal2 26488 12656 26488 12656 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[0\]
rlabel metal3 3248 15512 3248 15512 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[10\]
rlabel metal2 5880 15344 5880 15344 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[11\]
rlabel metal2 4648 14168 4648 14168 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[12\]
rlabel metal2 3304 13496 3304 13496 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[13\]
rlabel metal2 5096 12656 5096 12656 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[14\]
rlabel metal2 5992 11872 5992 11872 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[15\]
rlabel metal2 7672 12712 7672 12712 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[16\]
rlabel metal2 11816 17248 11816 17248 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[1\]
rlabel metal3 10360 17416 10360 17416 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[2\]
rlabel metal2 5992 15848 5992 15848 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[3\]
rlabel metal2 9688 17808 9688 17808 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[4\]
rlabel metal2 9688 20552 9688 20552 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[5\]
rlabel metal2 8624 21784 8624 21784 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[6\]
rlabel metal2 6776 19936 6776 19936 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[7\]
rlabel metal3 6048 20104 6048 20104 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[8\]
rlabel metal2 4536 18480 4536 18480 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[9\]
rlabel metal2 35224 31304 35224 31304 0 tt_um_rejunity_ay8913.noise_generator.period\[0\]
rlabel metal3 33656 29400 33656 29400 0 tt_um_rejunity_ay8913.noise_generator.period\[1\]
rlabel metal2 34776 33040 34776 33040 0 tt_um_rejunity_ay8913.noise_generator.period\[2\]
rlabel metal2 40488 29176 40488 29176 0 tt_um_rejunity_ay8913.noise_generator.period\[3\]
rlabel metal2 37744 29400 37744 29400 0 tt_um_rejunity_ay8913.noise_generator.period\[4\]
rlabel metal2 13720 12432 13720 12432 0 tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0
rlabel metal2 28056 13440 28056 13440 0 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal
rlabel metal2 36120 28672 36120 28672 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\]
rlabel metal2 33992 25816 33992 25816 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\]
rlabel metal2 36344 24976 36344 24976 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\]
rlabel metal2 36456 24304 36456 24304 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\]
rlabel metal2 36344 25816 36344 25816 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[4\]
rlabel metal2 7952 9800 7952 9800 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[2\]
rlabel metal3 8120 8232 8120 8232 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[3\]
rlabel metal2 8288 6776 8288 6776 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[4\]
rlabel metal2 7728 5096 7728 5096 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[5\]
rlabel metal2 10248 3808 10248 3808 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[6\]
rlabel metal2 12880 5208 12880 5208 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[7\]
rlabel metal2 13944 5432 13944 5432 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[8\]
rlabel metal2 15624 5040 15624 5040 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[9\]
rlabel metal2 23800 9688 23800 9688 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[2\]
rlabel metal2 20328 11256 20328 11256 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[3\]
rlabel metal2 19712 9912 19712 9912 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[4\]
rlabel metal3 12040 9912 12040 9912 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[5\]
rlabel metal2 11144 7504 11144 7504 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[6\]
rlabel metal2 13272 7728 13272 7728 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[7\]
rlabel metal2 13944 7280 13944 7280 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[8\]
rlabel metal2 17472 6776 17472 6776 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[9\]
rlabel metal2 27272 10808 27272 10808 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[2\]
rlabel metal2 25816 12376 25816 12376 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[3\]
rlabel metal2 23016 13272 23016 13272 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[4\]
rlabel metal2 19768 13384 19768 13384 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[5\]
rlabel metal2 16072 13664 16072 13664 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[6\]
rlabel metal2 17976 12992 17976 12992 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
rlabel metal2 15736 10136 15736 10136 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[8\]
rlabel metal2 18928 5208 18928 5208 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[9\]
rlabel metal2 20888 3920 20888 3920 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[10\]
rlabel metal2 30128 6776 30128 6776 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[2\]
rlabel metal2 30520 5432 30520 5432 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[3\]
rlabel metal2 27720 5544 27720 5544 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[4\]
rlabel metal2 27664 7448 27664 7448 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[5\]
rlabel metal2 26264 8372 26264 8372 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[6\]
rlabel metal2 22736 7672 22736 7672 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[7\]
rlabel metal3 23352 4312 23352 4312 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[8\]
rlabel metal2 21784 7504 21784 7504 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[9\]
rlabel metal2 45360 21448 45360 21448 0 tt_um_rejunity_ay8913.restart_envelope
rlabel metal2 37240 4256 37240 4256 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\]
rlabel metal3 35840 10696 35840 10696 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\]
rlabel metal2 34552 9856 34552 9856 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
rlabel metal2 31864 6328 31864 6328 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\]
rlabel metal2 34272 6776 34272 6776 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
rlabel metal2 46648 8344 46648 8344 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal2 44240 6552 44240 6552 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal3 36512 8232 36512 8232 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 41664 6776 41664 6776 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal2 43120 5208 43120 5208 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 43736 5824 43736 5824 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal2 45248 8120 45248 8120 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal2 46480 5992 46480 5992 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal2 46984 6272 46984 6272 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal3 48552 9016 48552 9016 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\]
rlabel metal2 26712 20524 26712 20524 0 tt_um_rejunity_ay8913.tone_A
rlabel metal2 23128 30072 23128 30072 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[0\]
rlabel metal2 15624 18480 15624 18480 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[10\]
rlabel metal3 18424 20776 18424 20776 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[11\]
rlabel metal2 24024 28952 24024 28952 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[1\]
rlabel metal2 18760 27832 18760 27832 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[2\]
rlabel metal2 15288 27160 15288 27160 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[3\]
rlabel metal2 15176 26656 15176 26656 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[4\]
rlabel metal3 16800 26376 16800 26376 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[5\]
rlabel metal3 15064 23016 15064 23016 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[6\]
rlabel metal2 15512 24360 15512 24360 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[7\]
rlabel metal2 13160 21168 13160 21168 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[8\]
rlabel metal2 16184 15680 16184 15680 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[9\]
rlabel metal2 24920 27384 24920 27384 0 tt_um_rejunity_ay8913.tone_A_generator.period\[0\]
rlabel metal2 21336 18144 21336 18144 0 tt_um_rejunity_ay8913.tone_A_generator.period\[10\]
rlabel metal2 22456 19320 22456 19320 0 tt_um_rejunity_ay8913.tone_A_generator.period\[11\]
rlabel metal2 19880 28840 19880 28840 0 tt_um_rejunity_ay8913.tone_A_generator.period\[1\]
rlabel metal2 21784 27832 21784 27832 0 tt_um_rejunity_ay8913.tone_A_generator.period\[2\]
rlabel metal2 25256 26040 25256 26040 0 tt_um_rejunity_ay8913.tone_A_generator.period\[3\]
rlabel metal2 22456 24920 22456 24920 0 tt_um_rejunity_ay8913.tone_A_generator.period\[4\]
rlabel metal2 21784 25872 21784 25872 0 tt_um_rejunity_ay8913.tone_A_generator.period\[5\]
rlabel metal2 17864 24584 17864 24584 0 tt_um_rejunity_ay8913.tone_A_generator.period\[6\]
rlabel metal2 22568 25424 22568 25424 0 tt_um_rejunity_ay8913.tone_A_generator.period\[7\]
rlabel metal2 17864 16128 17864 16128 0 tt_um_rejunity_ay8913.tone_A_generator.period\[8\]
rlabel metal2 18200 17080 18200 17080 0 tt_um_rejunity_ay8913.tone_A_generator.period\[9\]
rlabel metal3 31920 20888 31920 20888 0 tt_um_rejunity_ay8913.tone_B
rlabel metal2 34776 34552 34776 34552 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[0\]
rlabel metal2 27944 32928 27944 32928 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[10\]
rlabel metal2 30296 28504 30296 28504 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[11\]
rlabel metal2 36120 35784 36120 35784 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[1\]
rlabel metal2 35168 41832 35168 41832 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[2\]
rlabel metal3 36176 45080 36176 45080 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[3\]
rlabel metal2 34048 44296 34048 44296 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[4\]
rlabel metal3 32592 42504 32592 42504 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[5\]
rlabel metal2 27944 44352 27944 44352 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[6\]
rlabel metal3 28672 43400 28672 43400 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[7\]
rlabel metal3 29456 35672 29456 35672 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[8\]
rlabel metal2 28392 35112 28392 35112 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[9\]
rlabel metal2 39256 38024 39256 38024 0 tt_um_rejunity_ay8913.tone_B_generator.period\[0\]
rlabel metal2 31080 25312 31080 25312 0 tt_um_rejunity_ay8913.tone_B_generator.period\[10\]
rlabel metal2 32984 24472 32984 24472 0 tt_um_rejunity_ay8913.tone_B_generator.period\[11\]
rlabel metal2 36288 38920 36288 38920 0 tt_um_rejunity_ay8913.tone_B_generator.period\[1\]
rlabel metal2 36960 41048 36960 41048 0 tt_um_rejunity_ay8913.tone_B_generator.period\[2\]
rlabel metal2 35168 42728 35168 42728 0 tt_um_rejunity_ay8913.tone_B_generator.period\[3\]
rlabel metal3 31304 42728 31304 42728 0 tt_um_rejunity_ay8913.tone_B_generator.period\[4\]
rlabel metal3 31920 42504 31920 42504 0 tt_um_rejunity_ay8913.tone_B_generator.period\[5\]
rlabel metal3 28112 42840 28112 42840 0 tt_um_rejunity_ay8913.tone_B_generator.period\[6\]
rlabel metal2 27720 41664 27720 41664 0 tt_um_rejunity_ay8913.tone_B_generator.period\[7\]
rlabel metal3 29456 33320 29456 33320 0 tt_um_rejunity_ay8913.tone_B_generator.period\[8\]
rlabel metal2 28168 22960 28168 22960 0 tt_um_rejunity_ay8913.tone_B_generator.period\[9\]
rlabel metal2 29848 21280 29848 21280 0 tt_um_rejunity_ay8913.tone_C
rlabel metal2 24808 33656 24808 33656 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[0\]
rlabel metal3 17976 31192 17976 31192 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[10\]
rlabel metal2 20328 30072 20328 30072 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[11\]
rlabel metal2 23800 33600 23800 33600 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[1\]
rlabel metal2 22344 36512 22344 36512 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[2\]
rlabel metal2 16408 41888 16408 41888 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[3\]
rlabel metal2 19208 42112 19208 42112 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[4\]
rlabel metal2 16408 40432 16408 40432 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[5\]
rlabel metal2 15456 38696 15456 38696 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[6\]
rlabel metal2 17864 38668 17864 38668 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[7\]
rlabel metal3 16688 34104 16688 34104 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[8\]
rlabel metal2 15232 32424 15232 32424 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[9\]
rlabel metal2 23912 36792 23912 36792 0 tt_um_rejunity_ay8913.tone_C_generator.period\[0\]
rlabel metal2 24584 24164 24584 24164 0 tt_um_rejunity_ay8913.tone_C_generator.period\[10\]
rlabel metal3 22792 22456 22792 22456 0 tt_um_rejunity_ay8913.tone_C_generator.period\[11\]
rlabel metal2 24696 36736 24696 36736 0 tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
rlabel metal2 22680 39144 22680 39144 0 tt_um_rejunity_ay8913.tone_C_generator.period\[2\]
rlabel metal3 23800 40488 23800 40488 0 tt_um_rejunity_ay8913.tone_C_generator.period\[3\]
rlabel via2 21336 41048 21336 41048 0 tt_um_rejunity_ay8913.tone_C_generator.period\[4\]
rlabel metal2 21560 43176 21560 43176 0 tt_um_rejunity_ay8913.tone_C_generator.period\[5\]
rlabel metal2 18872 45864 18872 45864 0 tt_um_rejunity_ay8913.tone_C_generator.period\[6\]
rlabel metal2 21224 43120 21224 43120 0 tt_um_rejunity_ay8913.tone_C_generator.period\[7\]
rlabel metal2 21560 21056 21560 21056 0 tt_um_rejunity_ay8913.tone_C_generator.period\[8\]
rlabel metal2 19432 23016 19432 23016 0 tt_um_rejunity_ay8913.tone_C_generator.period\[9\]
rlabel metal2 26824 17416 26824 17416 0 tt_um_rejunity_ay8913.tone_disable_A
rlabel metal2 32928 17752 32928 17752 0 tt_um_rejunity_ay8913.tone_disable_B
rlabel metal2 31192 18872 31192 18872 0 tt_um_rejunity_ay8913.tone_disable_C
rlabel metal3 24584 24696 24584 24696 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 51000 51000
<< end >>
